// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Thu Jan 30 13:05:32 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_c_1, ENCODER0_B_c_0, 
        ENCODER1_A_c_1, ENCODER1_B_c_0, NEOPXL_c, DE_c, RX_c, INHC_c, 
        INLB_c, INHB_c, INLA_c, INHA_c;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(39[11:13])
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(41[13:25])
    
    wire hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(87[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(88[21:25])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(122[22:39])
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(123[21:45])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(124[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(125[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(126[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(127[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(128[22:24])
    
    wire n31327;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(130[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(131[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(132[22:35])
    
    wire n31195, n3957, n14, n31326;
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(162[22:33])
    
    wire n31325;
    wire [31:0]data;   // verilog/TinyFPGA_B.v(206[15:19])
    
    wire data_ready, n31194, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(229[11:24])
    
    wire read;
    wire [22:0]pwm_setpoint_22__N_11;
    
    wire RX_N_10;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [31:0]motor_state_23__N_82;
    wire [25:0]encoder0_position_scaled_23__N_34;
    wire [23:0]displacement_23__N_58;
    
    wire n5180, n31193, n31192, n31324, n31323, n31191;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    
    wire start, \neo_pixel_transmitter.done ;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n5442, n31190, n22424, n35562;
    wire [3:0]state_3__N_369;
    
    wire n34460, n27400, n31322, n28054, n22423, n22422, n31189, 
        n31321, n31320, n22421, n22420, n22419, n22418, n22417, 
        n22416, n22415, n22414, n22413, n22412, n22411, n20602, 
        n31188, \neo_pixel_transmitter.done_N_583 , n31319, n28050, 
        n31187, n31186, n425;
    wire [31:0]pwm_counter;   // verilog/pwm.v(11[9:20])
    
    wire n15, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
        n13, n14_adj_4855, n15_adj_4856, n16, n17, n18, n19, n20, 
        n21, n22, n23, n24, n25, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(91[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(95[12:19])
    
    wire n31318, n31185, n28040;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(97[12:26])
    
    wire tx_active, n31317, n31316, n14_adj_4857, n10_adj_4858, n31184, 
        n31315, n10_adj_4859, n12_adj_4860, n7_adj_4861, n31183, n20_adj_4862, 
        n18_adj_4863, n16_adj_4864, n31182, n31314, n31181, n31313, 
        n31180, n31179, n31312, n31178, n31177, n26980, n27990, 
        n31311, n27986, n31310, n31309, n31176, n31175, n31308, 
        n31174, n31307, n31173, n31172, n31171, n31306, n31170, 
        n31169, n31305, n31304, n31168, n31303, n27974, n31167, 
        n31302, n27942, n31166, n27938, n31165, n7_adj_4865, n31164, 
        n31163, n31301, n31300, n31162, n31161, n31160, n40105, 
        n31299, n31159, n31158, n31028, n31298, n31297, n31157, 
        n31296, n31027, n31156, n31155, n31154, n27926, n31026, 
        n31295, n31153, n31294, n40109, n31293, n31025, n40035, 
        n31292, n28004, n31291, n31024, n15_adj_4866, n14_adj_4867, 
        n40054, n37894, n4_adj_4868, n31152, n31023, n31151, n31022, 
        n31150, n31149, n31290, n31148, n12_adj_4869, n11_adj_4870, 
        n10_adj_4871, n40034, n31289, n31147, n31288, n31146, n31021, 
        n31287, n31286, n31145, n31144, n31020, n31285, n31284, 
        n31143, n31283, n31282, n31019, n31281, n27970, n31280, 
        n31279, n31278, n31018, n31277, n31276, n31275, n31017, 
        n39945, n31274, n39943, n31273, n31272, n31016, n39938, 
        n39932, n31015, n31271, n39926, n31270, n39924, n31014, 
        n39861, n31269, n31013, n31134, n31012, n31133, n31268, 
        n31267, n31011, n31010, n31132, n31266, n31131, n31009, 
        n31008, n31130, n31007, n31265, n31264, n6_adj_4872, n31129, 
        n31128, n31006, n31127, n31126, n31263, n31395, n31262, 
        n31394, n31125, n31393, n31124, n31261, n31260, n31392, 
        n31391, n31259, n31258, n31123, n31257, n31122, n31390, 
        n31256, n5440, n31255, n31254, n31389, n24_adj_4873, n21_adj_4874, 
        n20_adj_4875, n17_adj_4876, n31121, n31253, n31120, n39620, 
        n31252, n39610, n31119, n31388, n31251, n31118, n31250, 
        n31117, n31249, n31116, n30761, n30760, n31387, n31248, 
        n31115, n36330, n4_adj_4877, n30759, n31386, n31114, n31113, 
        n31112, n31111, n35561, n12_adj_4878, n37487, n35272, n31110, 
        n39875, n40291, n27830, n31385, n28094, n37529, n8_adj_4879, 
        n31384, n25_adj_4880, n24_adj_4881, n23_adj_4882, n22_adj_4883, 
        n21_adj_4884, n20_adj_4885, n19_adj_4886, n18_adj_4887, n17_adj_4888, 
        n16_adj_4889, n15_adj_4890, n14_adj_4891, n13_adj_4892, n12_adj_4893, 
        n11_adj_4894, n10_adj_4895, n9_adj_4896, n8_adj_4897, n7_adj_4898, 
        n6_adj_4899, n5_adj_4900, n22856, n22855, n22854, n22853, 
        n22852, n22851, n22850, n22849, n22848, n22847, n34, n22843, 
        n22840, n22839, n33, n32, n22838, n31, n22837, n22836, 
        n22835, n22834, n31247, n31109, n31383, n31382, n30758, 
        n31108, n31107, n31106, n30757, n31246, n31245, n31244, 
        n31243, n31242, n31105, n31381, n31241, n31240, n31380, 
        n30756, n30, n30755, n36440, n22833, n22832, n22831, n22830, 
        n22829, n22828, n22827, n22826, n22825, n22824, n22823, 
        n22822, n22821, n22820, n22819, n22818, n22817, n22814, 
        n39791, n22813, n22812, n22811, n22810, n22809, n22808, 
        n22807, n22806, n22805, n22804, n22803, n22802, n22801, 
        n22800, n22799, n22798, n22797, n32024, n32023, n32022, 
        n22796, n22795, n22794, n22793, n22792, n22791, n22790, 
        n22789, n22788, n32021, n32020, n22787, n22786, n22785, 
        n22784, n22783, n22782, n22781, n22780, n22779, n22778, 
        n22777, n15_adj_4901, n22776, n10_adj_4902, n22775, n22774, 
        n22773, n22772, n22771, n22770, n22769, n22768, n22767, 
        n22766, n22765, n22764, n22763, n22762, n22761, n22760, 
        n22759, n22758, n22757, n22756, n22755, n22754, n22753, 
        n22752, n22751, n36368, n22750, n22749, n31379, n31378, 
        n31239, n31238, n31237, n31236, n31377, n31376, n39793, 
        n31375, n31235, n31234, n31374, n31373, n31372, n31371, 
        n30754, n31370, n22748, n22747, n22746, n22745, n22744, 
        n22743, n22742, n22741, n22740, n22739, n22738, n22737, 
        n22736, n22735, n22734, n22733, n22732, n22731, n22730, 
        n22729, n22728, quadA_debounced, quadB_debounced, n3461, n22727, 
        n22726, n22725, n4_adj_4903, n3_adj_4904, n2, n22724, n27098, 
        n22721, n22720, n22719, n22718, quadA_debounced_adj_4905, 
        quadB_debounced_adj_4906, n22717, n22716, n22715, n22714, 
        n22713, n22712, n22711, n22710, n22709, n22708, n22707, 
        n22706, n22705, n22704, n22703, n22702, n22701, n22700, 
        n22699, n22698, n22697, n22696, n22695, n22694, n22693, 
        n22692, n22691, n22690, n22689, n22688, n22687, n22686, 
        n22685, n22684, n22683, n22682, n22681, n22680, n22679, 
        n22678, rw;
    wire [7:0]state_adj_5082;   // verilog/eeprom.v(22[11:16])
    
    wire n22677, n22676, n22675, n22674, n22673, n22672, n10_adj_4908, 
        n22671, n22670, n22370, n22669, n22668, n22667, n22666, 
        n22665, n22664, n22663, n22662, n22661, n22660, n22659, 
        n22658, n22657, n20604, n22369, n22656, n22655, n22654, 
        n22653, n22652, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    
    wire n22651, n22650, n31233, n22649, n22648, n22647, n22646, 
        n22645, n22644, n22643, n22642, n22641, n22640, n22639, 
        n22638, n22637, n22636, n22635, n22634, n30753, n22633, 
        n5445, n22632, n22_adj_4909, n22631, n22630, n22629, n20_adj_4910, 
        n22628, n22627, n22626, n22625, n22368, n22624, n22623, 
        n22622, n22621, n22620, n22619, n22618, n22617, n22616, 
        n22615, n22614, n22613, n22612, n18_adj_4911;
    wire [2:0]r_SM_Main_adj_5088;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_Bit_Index_adj_5090;   // verilog/uart_tx.v(33[16:27])
    
    wire n13_adj_4913;
    wire [2:0]r_SM_Main_2__N_3454;
    
    wire n22611, n22610, n28078, n22609, n22608, n4_adj_4914, n22367, 
        n22607, n22606, n22605, n22604, n22603, n22602, n22601, 
        n22600, n22599, n22598, n22597, n22596, n22595, n22594, 
        n22593, n22592, n22591, n22590, n22589, n22588, n22587, 
        n22586, n22585;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n22584, n22583, n22582, n22581, n22580, n22579, n22578;
    wire [1:0]reg_B_adj_5099;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n22577, n15_adj_4917, n22576, n22575, n22574;
    wire [7:0]state_adj_5111;   // verilog/i2c_controller.v(32[12:17])
    
    wire n37048;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(33[12:22])
    
    wire n22573, n22366, scl_enable_N_3958;
    wire [7:0]state_7__N_3865;
    
    wire n22291, n22572, n4_adj_4920, n39335, n22571, n4_adj_4921, 
        n22365, n4760, n5444, n22570, n22569, n22568;
    wire [7:0]state_7__N_3881;
    
    wire n22567, n39329, n22566, n22565, n22564, n22563, n22562, 
        n22561, n22560, n39327, n22559, n22558, n22557, n22556, 
        n22555, n22364, n22363, n22362, n22361, n22360, n22359, 
        n22358, n22357, n22554, n22553, n22552, n22551, n22550, 
        n22549, n22548, n15_adj_4922, n22547, n22546, n22545, n22544, 
        n22543, n22542, n20608, n22541, n22540, n22539, n22538, 
        n3_adj_4923, n5_adj_4924, n6_adj_4925, n7_adj_4926, n8_adj_4927, 
        n9_adj_4928, n10_adj_4929, n11_adj_4930, n12_adj_4931, n13_adj_4932, 
        n14_adj_4933, n15_adj_4934, n16_adj_4935, n17_adj_4936, n18_adj_4937, 
        n19_adj_4938, n20_adj_4939, n21_adj_4940, n22_adj_4941, n23_adj_4942, 
        n24_adj_4943, n25_adj_4944, n4_adj_4945, n22195, n509, n510, 
        n511, n513, n514, n515, n516, n517, n518, n519, n520, 
        n521, n522, n523, n524, n525, n526, n527, n528, n529, 
        n530, n531, n532, n22193, n22012, n39323, n39321, n619, 
        n674, n675, n676, n677, n678, n679, n700, n728, n729, 
        n730, n731, n732, n733, n752, n753, n754, n755, n756, 
        n757, n758, n778, n806, n807, n808, n809, n810, n811, 
        n812, n830, n831, n832, n833, n834, n835, n836, n837, 
        n856, n883, n884, n885, n886, n887, n888, n889, n890, 
        n891, n908, n909, n910, n911, n912, n913, n914, n915, 
        n916, n40392, n934, n37217, n961, n962, n963, n964, 
        n965, n966, n967, n968, n969, n970, n986, n987, n988, 
        n989, n990, n991, n992, n993, n994, n995, n1012, n1040, 
        n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, 
        n1049, n35575, n1064, n1065, n1066, n1067, n1068, n1069, 
        n1070, n1071, n1072, n1073, n1074, n1090, n1117, n1118, 
        n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, 
        n1127, n1128, n22157, n1142, n1143, n1144, n1145, n1146, 
        n1147, n1148, n1149, n1150, n1151, n1152, n1153, n40353, 
        n1168, n1195, n1196, n1197, n1198, n1199, n1200, n1201, 
        n1202, n1203, n1204, n1205, n1206, n1207, n21971, n1220, 
        n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, 
        n1229, n1230, n1231, n1232, n1246, n21969, n1273, n1274, 
        n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
        n1283, n1284, n1285, n1286, n1298, n1299, n1300, n1301, 
        n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, 
        n1310, n1311, n1324, n1351, n1352, n1353, n1354, n1355, 
        n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, 
        n1364, n1365, n1376, n1377, n1378, n1379, n1380, n1381, 
        n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, 
        n1390, n1402, n1429, n1430, n1431, n1432, n1433, n1434, 
        n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, 
        n1443, n1444, n1454, n1455, n1456, n1457, n1458, n1459, 
        n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, 
        n1468, n1469, n1480, n1507, n1508, n1509, n1510, n1511, 
        n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, 
        n1520, n1521, n1522, n1523, n1532, n1533, n1534, n1535, 
        n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, 
        n1544, n1545, n1546, n1547, n1548, n1558, n1585, n1586, 
        n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, 
        n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, 
        n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, 
        n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, 
        n1626, n1627, n1636, n1663, n1664, n1665, n1666, n1667, 
        n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
        n1676, n1677, n1678, n1679, n1680, n1681, n1688, n1689, 
        n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, 
        n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, 
        n1706, n1714, n1741, n1742, n1743, n1744, n1745, n1746, 
        n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, 
        n1755, n1756, n1757, n1758, n1759, n1760, n1766, n1767, 
        n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, 
        n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, 
        n1784, n1785, n1792, n1819, n1820, n1821, n1822, n1823, 
        n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, 
        n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, 
        n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, 
        n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, 
        n1860, n1861, n1862, n1863, n1864, n1870, n1897, n1898, 
        n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, 
        n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, 
        n1915, n1916, n1917, n1918, n1922, n1923, n1924, n1925, 
        n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, 
        n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, 
        n1942, n1943, n1948, n1975, n1976, n1977, n1978, n1979, 
        n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, 
        n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, 
        n1996, n1997, n2000, n2001, n2002, n2003, n2004, n2005, 
        n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, 
        n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, 
        n2022, n2026, n2053, n2054, n2055, n2056, n2057, n2058, 
        n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, 
        n2067, n2068, n2069, n2070, n2071, n2073, n2076, n28106, 
        n35568, n5701, n5700, n5699, n5698, n5697, n5696, n5695, 
        n5694, n5693, n5692, n5691, n5690, n5689, n5688, n5687, 
        n5686, n5685, n5684, n5683, n5681, n5680, n5443, n37568, 
        n37536, n62, n5_adj_4946, n21920, n14_adj_4947, n35362, 
        n10_adj_4948, n30752, n21865, n6_adj_4949, n39289, n39285, 
        n34_adj_4950, n31_adj_4951, n22356, n22355, n30_adj_4952, 
        n28, n40110, n20716, n22354, n22353, n22352, n22_adj_4953, 
        n21_adj_4954, n22351, n22350, n22349, n4_adj_4955, n6_adj_4956, 
        n7_adj_4957, n8_adj_4958, n9_adj_4959, n10_adj_4960, n11_adj_4961, 
        n12_adj_4962, n13_adj_4963, n15_adj_4964, n17_adj_4965, n19_adj_4966, 
        n21_adj_4967, n39944, n23_adj_4968, n25_adj_4969, n27, n39942, 
        n29, n30_adj_4970, n31_adj_4971, n33_adj_4972, n35, n35585, 
        n39272, n39271, n31232, n31369, n31231, n31368, n31367, 
        n31366, n31365, n31230, n31229, n31228, n40620, n37256, 
        n28_adj_4973, n27_adj_4974, n26, n25_adj_4975, n134, n135, 
        n136, n137, n138, n139, n140, n141, n142, n143, n144, 
        n145, n146, n147, n148, n149, n150, n151, n152, n153, 
        n154, n155, n156, n157, n158, n159, n160, n161, n162, 
        n163, n164, n165, n22348, n22347, n22346, n22345, n22344, 
        n22343, n22342, n22341, n22340, n22339, n22338, n22337, 
        n22336, n22335, n22334, n22333, n22330, n22326, n22322, 
        n22321, n22320, n22319, n22318, n22498, n22497, n22496, 
        n22495, n22494, n22493, n35254, n31364, n31363, n22492, 
        n22491, n22490, n22489, n22488, n22487, n22486, n22485, 
        n22484, n22483, n22482, n22481, n22480, n22479, n22478, 
        n22477, n22476, n22475, n31362, n22316, n22315, n22314, 
        n22312, n22311, n22310, n22309, n22308, n22307, n22306, 
        n22305, n22304, n22303, n22302, n22300, n35579, n22434, 
        n22433, n22432, n22431, n22430, n22429, n22428, n22427, 
        n22426, n22425, n37470, n2_adj_4976, n3_adj_4977, n4_adj_4978, 
        n5_adj_4979, n6_adj_4980, n7_adj_4981, n8_adj_4982, n9_adj_4983, 
        n10_adj_4984, n11_adj_4985, n12_adj_4986, n13_adj_4987, n14_adj_4988, 
        n15_adj_4989, n16_adj_4990, n17_adj_4991, n18_adj_4992, n19_adj_4993, 
        n20_adj_4994, n21_adj_4995, n22_adj_4996, n23_adj_4997, n24_adj_4998, 
        n25_adj_4999, n4_adj_5000, n31361, n34038, n31227, n31226, 
        n31360, n31816, n31815, n31814, n31813, n31812, n31811, 
        n31810, n31809, n31808, n31807, n31806, n31805, n31804, 
        n31803, n37465, n31802, n31801, n31800, n31799, n31798, 
        n31225, n31797, n31359, n31796, n31795, n31794, n31793, 
        n40108, n30751, n6_adj_5001, n31358, n31357, n31224, n31223, 
        n31356, n31355, n31222, n31221, n31220, n31219, n31218, 
        n13_adj_5002, n30750, n31354, n23_adj_5003, n27_adj_5004, 
        n29_adj_5005, n31353, n30749, n31217, n37, n31216, n39, 
        n43, n45, n49, n35586, n27944, n26_adj_5006, n24_adj_5007, 
        n22_adj_5008, n18_adj_5009, n13920, n31215, n10_adj_5010, 
        n30748, n31352, n31351, n31350, n31214, n31213, n4_adj_5011, 
        n35591, n41168, n22299, n22298, n39214, n31349, n31212, 
        n31348, n16_adj_5012, n31211, n12_adj_5013, n22297, n27086, 
        n38219, n10_adj_5014, n31347, n37680, n20776, n39198, n39196, 
        n30747, n30746, n31346, n22296, n22295, n31210, n22294, 
        n30745, n31345, n31344, n30744, n31209, n7_adj_5015, n36883, 
        n31208, n31343, n31342, n31207, n31206, n31205, n31341, 
        n31204, n31340, n31203, n31339, n38316, n31552, n37535, 
        n31551, n31338, n31337, n31550, n31549, n30743, n31336, 
        n31548, n31547, n31202, n31335, n31546, n31545, n31544, 
        n36364, n31334, n31543, n31542, n31541, n31540, n31539, 
        n22292, n30742, n31333, n31201, n31538, n31537, n31536, 
        n8_adj_5016, n31535, n31534, n31533, n31532, n31332, n31531, 
        n30741, n30740, n7_adj_5017, n31530, n31529, n12_adj_5018, 
        n31528, n31527, n36334, n36332, n11_adj_5019, n31526, n31525, 
        n31524, n31331, n31523, n31200, n31522, n17_adj_5020, n20781, 
        n16_adj_5021, n20726, n5_adj_5022, n28098, n10_adj_5023, n4_adj_5024, 
        n6_adj_5025, n31199, n20731, n31330, n15_adj_5026, n14_adj_5027, 
        n31198, n31329, n31197, n18082, n37463, n6_adj_5028, n5_adj_5029, 
        n37237, n31196, n31328, n28072, n37_adj_5030, n36, n30_adj_5031, 
        n29_adj_5032, n28_adj_5033, n27_adj_5034, n26_adj_5035, n25_adj_5036, 
        n24_adj_5037, n23_adj_5038, n22_adj_5039, n21_adj_5040, n36901;
    
    VCC i2 (.Y(VCC_net));
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.encoder0_position({encoder0_position}), 
            .GND_net(GND_net), .clk32MHz(clk32MHz), .data_o({quadA_debounced, 
            quadB_debounced}), .n38219(n38219), .reg_B({reg_B}), .VCC_net(VCC_net), 
            .ENCODER0_B_c_0(ENCODER0_B_c_0), .n22848(n22848), .n22316(n22316), 
            .ENCODER0_A_c_1(ENCODER0_A_c_1)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(185[15] 190[4])
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF h3_44 (.Q(INLB_c), .C(clk32MHz), .D(hall3));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_58[0]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF h2_43 (.Q(INHB_c), .C(clk32MHz), .D(hall2));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(state_7__N_3881[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    neopixel nx (.GND_net(GND_net), .VCC_net(VCC_net), .clk32MHz(clk32MHz), 
            .\neo_pixel_transmitter.done (\neo_pixel_transmitter.done ), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .start(start), .\state[1] (state[1]), .LED_c(LED_c), .\state_3__N_369[1] (state_3__N_369[1]), 
            .n14(n14), .n36364(n36364), .n21969(n21969), .timer({timer}), 
            .n37680(n37680), .neopxl_color({neopxl_color}), .n22814(n22814), 
            .n22813(n22813), .n22812(n22812), .n22811(n22811), .n22810(n22810), 
            .n22809(n22809), .n22808(n22808), .n22807(n22807), .n22806(n22806), 
            .n22805(n22805), .n22804(n22804), .n22803(n22803), .n22802(n22802), 
            .n22801(n22801), .n22800(n22800), .n22799(n22799), .n22798(n22798), 
            .n22797(n22797), .n22796(n22796), .n22795(n22795), .n22794(n22794), 
            .n22793(n22793), .n22792(n22792), .n22791(n22791), .n22790(n22790), 
            .n22789(n22789), .n22788(n22788), .n22787(n22787), .n22786(n22786), 
            .n22785(n22785), .n22784(n22784), .n22326(n22326), .\neo_pixel_transmitter.done_N_583 (\neo_pixel_transmitter.done_N_583 ), 
            .NEOPXL_c(NEOPXL_c), .n34460(n34460), .n22291(n22291), .n39196(n39196)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(43[10] 49[2])
    SB_LUT4 add_644_4_lut (.I0(duty[2]), .I1(n40620), .I2(n23), .I3(n30741), 
            .O(pwm_setpoint_22__N_11[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_7 (.CI(n31797), 
            .I0(GND_net), .I1(n21_adj_4995), .CO(n31798));
    SB_LUT4 unary_minus_4_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_DFF dir_48 (.Q(INHC_c), .C(clk32MHz), .D(duty[23]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_4996), .I3(n31796), .O(n22_adj_4883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1311_3_lut (.I0(n1923), .I1(n1976), 
            .I2(n1948), .I3(GND_net), .O(n2001));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1271_3_lut (.I0(n1858), .I1(n1911), 
            .I2(n1870), .I3(GND_net), .O(n1936));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1271_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1265_3_lut (.I0(n1852), .I1(n1905), 
            .I2(n1870), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1265_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1266_3_lut (.I0(n1853), .I1(n1906), 
            .I2(n1870), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1266_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1274_3_lut (.I0(n1861), .I1(n1914), 
            .I2(n1870), .I3(GND_net), .O(n1939));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1274_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1269_3_lut (.I0(n1856), .I1(n1909), 
            .I2(n1870), .I3(GND_net), .O(n1934));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1269_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1275_3_lut (.I0(n1862), .I1(n1915), 
            .I2(n1870), .I3(GND_net), .O(n1940));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1275_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1258_3_lut (.I0(n1845), .I1(n1898), 
            .I2(n1870), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1258_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1262_3_lut (.I0(n1849), .I1(n1902), 
            .I2(n1870), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1262_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1270_3_lut (.I0(n1857), .I1(n1910), 
            .I2(n1870), .I3(GND_net), .O(n1935));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1270_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1263_3_lut (.I0(n1850), .I1(n1903), 
            .I2(n1870), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1263_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1259_3_lut (.I0(n1846), .I1(n1899), 
            .I2(n1870), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1259_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1264_3_lut (.I0(n1851), .I1(n1904), 
            .I2(n1870), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1264_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1268_3_lut (.I0(n1855), .I1(n1908), 
            .I2(n1870), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1268_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1261_3_lut (.I0(n1848), .I1(n1901), 
            .I2(n1870), .I3(GND_net), .O(n1926));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1261_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1278_3_lut (.I0(n530), .I1(n1918), 
            .I2(n1870), .I3(GND_net), .O(n1943));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1278_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1277_3_lut (.I0(n1864), .I1(n1917), 
            .I2(n1870), .I3(GND_net), .O(n1942));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1277_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1276_3_lut (.I0(n1863), .I1(n1916), 
            .I2(n1870), .I3(GND_net), .O(n1941));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1276_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3255_i2_3_lut (.I0(encoder0_position[1]), .I1(n24_adj_4881), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n531));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1204_3_lut (.I0(n1766), .I1(n1819), 
            .I2(n1792), .I3(GND_net), .O(n1844));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1204_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1209_3_lut (.I0(n1771), .I1(n1824), 
            .I2(n1792), .I3(GND_net), .O(n1849));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1209_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1205_3_lut (.I0(n1767), .I1(n1820), 
            .I2(n1792), .I3(GND_net), .O(n1845));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1205_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1212_3_lut (.I0(n1774), .I1(n1827), 
            .I2(n1792), .I3(GND_net), .O(n1852));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1212_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1213_3_lut (.I0(n1775), .I1(n1828), 
            .I2(n1792), .I3(GND_net), .O(n1853));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1213_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1215_3_lut (.I0(n1777), .I1(n1830), 
            .I2(n1792), .I3(GND_net), .O(n1855));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1215_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1211_3_lut (.I0(n1773), .I1(n1826), 
            .I2(n1792), .I3(GND_net), .O(n1851));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1211_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1207_3_lut (.I0(n1769), .I1(n1822), 
            .I2(n1792), .I3(GND_net), .O(n1847));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1207_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1208_3_lut (.I0(n1770), .I1(n1823), 
            .I2(n1792), .I3(GND_net), .O(n1848));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1208_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1210_3_lut (.I0(n1772), .I1(n1825), 
            .I2(n1792), .I3(GND_net), .O(n1850));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1210_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1217_3_lut (.I0(n1779), .I1(n1832), 
            .I2(n1792), .I3(GND_net), .O(n1857));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1217_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1219_3_lut (.I0(n1781), .I1(n1834), 
            .I2(n1792), .I3(GND_net), .O(n1859));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1219_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1216_3_lut (.I0(n1778), .I1(n1831), 
            .I2(n1792), .I3(GND_net), .O(n1856));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1216_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1206_3_lut (.I0(n1768), .I1(n1821), 
            .I2(n1792), .I3(GND_net), .O(n1846));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1206_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1220_3_lut (.I0(n1782), .I1(n1835), 
            .I2(n1792), .I3(GND_net), .O(n1860));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1220_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1221_3_lut (.I0(n1783), .I1(n1836), 
            .I2(n1792), .I3(GND_net), .O(n1861));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1221_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1218_3_lut (.I0(n1780), .I1(n1833), 
            .I2(n1792), .I3(GND_net), .O(n1858));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1218_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1156_3_lut (.I0(n1693), .I1(n1746), 
            .I2(n1714), .I3(GND_net), .O(n1771));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1156_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1151_3_lut (.I0(n1688), .I1(n1741), 
            .I2(n1714), .I3(GND_net), .O(n1766));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1151_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1158_3_lut (.I0(n1695), .I1(n1748), 
            .I2(n1714), .I3(GND_net), .O(n1773));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1158_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1155_3_lut (.I0(n1692), .I1(n1745), 
            .I2(n1714), .I3(GND_net), .O(n1770));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1155_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1165_3_lut (.I0(n1702), .I1(n1755), 
            .I2(n1714), .I3(GND_net), .O(n1780));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1165_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1154_3_lut (.I0(n1691), .I1(n1744), 
            .I2(n1714), .I3(GND_net), .O(n1769));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1154_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1161_3_lut (.I0(n1698), .I1(n1751), 
            .I2(n1714), .I3(GND_net), .O(n1776));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1161_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1153_3_lut (.I0(n1690), .I1(n1743), 
            .I2(n1714), .I3(GND_net), .O(n1768));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1153_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1159_3_lut (.I0(n1696), .I1(n1749), 
            .I2(n1714), .I3(GND_net), .O(n1774));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1159_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1162_3_lut (.I0(n1699), .I1(n1752), 
            .I2(n1714), .I3(GND_net), .O(n1777));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1162_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1163_3_lut (.I0(n1700), .I1(n1753), 
            .I2(n1714), .I3(GND_net), .O(n1778));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1163_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1164_3_lut (.I0(n1701), .I1(n1754), 
            .I2(n1714), .I3(GND_net), .O(n1779));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1164_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1160_3_lut (.I0(n1697), .I1(n1750), 
            .I2(n1714), .I3(GND_net), .O(n1775));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1160_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1152_3_lut (.I0(n1689), .I1(n1742), 
            .I2(n1714), .I3(GND_net), .O(n1767));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1152_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1157_3_lut (.I0(n1694), .I1(n1747), 
            .I2(n1714), .I3(GND_net), .O(n1772));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1157_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1168_3_lut (.I0(n1705), .I1(n1758), 
            .I2(n1714), .I3(GND_net), .O(n1783));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1168_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1166_3_lut (.I0(n1703), .I1(n1756), 
            .I2(n1714), .I3(GND_net), .O(n1781));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1166_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1167_3_lut (.I0(n1704), .I1(n1757), 
            .I2(n1714), .I3(GND_net), .O(n1782));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1167_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1102_3_lut (.I0(n1614), .I1(n1667), 
            .I2(n1636), .I3(GND_net), .O(n1692));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1102_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1099_3_lut (.I0(n1611), .I1(n1664), 
            .I2(n1636), .I3(GND_net), .O(n1689));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1099_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1106_3_lut (.I0(n1618), .I1(n1671), 
            .I2(n1636), .I3(GND_net), .O(n1696));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1104_3_lut (.I0(n1616), .I1(n1669), 
            .I2(n1636), .I3(GND_net), .O(n1694));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1100_3_lut (.I0(n1612), .I1(n1665), 
            .I2(n1636), .I3(GND_net), .O(n1690));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1100_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1107_3_lut (.I0(n1619), .I1(n1672), 
            .I2(n1636), .I3(GND_net), .O(n1697));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1103_3_lut (.I0(n1615), .I1(n1668), 
            .I2(n1636), .I3(GND_net), .O(n1693));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1103_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1098_3_lut (.I0(n1610), .I1(n1663), 
            .I2(n1636), .I3(GND_net), .O(n1688));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1098_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1101_3_lut (.I0(n1613), .I1(n1666), 
            .I2(n1636), .I3(GND_net), .O(n1691));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1101_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1108_3_lut (.I0(n1620), .I1(n1673), 
            .I2(n1636), .I3(GND_net), .O(n1698));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1111_3_lut (.I0(n1623), .I1(n1676), 
            .I2(n1636), .I3(GND_net), .O(n1701));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1109_3_lut (.I0(n1621), .I1(n1674), 
            .I2(n1636), .I3(GND_net), .O(n1699));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1110_3_lut (.I0(n1622), .I1(n1675), 
            .I2(n1636), .I3(GND_net), .O(n1700));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1105_3_lut (.I0(n1617), .I1(n1670), 
            .I2(n1636), .I3(GND_net), .O(n1695));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1114_3_lut (.I0(n1626), .I1(n1679), 
            .I2(n1636), .I3(GND_net), .O(n1704));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1112_3_lut (.I0(n1624), .I1(n1677), 
            .I2(n1636), .I3(GND_net), .O(n1702));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1113_3_lut (.I0(n1625), .I1(n1678), 
            .I2(n1636), .I3(GND_net), .O(n1703));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1054_3_lut (.I0(n1541), .I1(n1594), 
            .I2(n1558), .I3(GND_net), .O(n1619));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1056_3_lut (.I0(n1543), .I1(n1596), 
            .I2(n1558), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1048_3_lut (.I0(n1535), .I1(n1588), 
            .I2(n1558), .I3(GND_net), .O(n1613));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1051_3_lut (.I0(n1538), .I1(n1591), 
            .I2(n1558), .I3(GND_net), .O(n1616));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1055_3_lut (.I0(n1542), .I1(n1595), 
            .I2(n1558), .I3(GND_net), .O(n1620));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1055_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1057_3_lut (.I0(n1544), .I1(n1597), 
            .I2(n1558), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1057_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1045_3_lut (.I0(n1532), .I1(n1585), 
            .I2(n1558), .I3(GND_net), .O(n1610));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1060_3_lut (.I0(n1547), .I1(n1600), 
            .I2(n1558), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1058_3_lut (.I0(n1545), .I1(n1598), 
            .I2(n1558), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1059_3_lut (.I0(n1546), .I1(n1599), 
            .I2(n1558), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1050_3_lut (.I0(n1537), .I1(n1590), 
            .I2(n1558), .I3(GND_net), .O(n1615));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1052_3_lut (.I0(n1539), .I1(n1592), 
            .I2(n1558), .I3(GND_net), .O(n1617));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1047_3_lut (.I0(n1534), .I1(n1587), 
            .I2(n1558), .I3(GND_net), .O(n1612));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1049_3_lut (.I0(n1536), .I1(n1589), 
            .I2(n1558), .I3(GND_net), .O(n1614));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1053_3_lut (.I0(n1540), .I1(n1593), 
            .I2(n1558), .I3(GND_net), .O(n1618));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1046_3_lut (.I0(n1533), .I1(n1586), 
            .I2(n1558), .I3(GND_net), .O(n1611));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1001_3_lut (.I0(n1463), .I1(n1516), 
            .I2(n1480), .I3(GND_net), .O(n1541));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i995_3_lut (.I0(n1457), .I1(n1510), 
            .I2(n1480), .I3(GND_net), .O(n1535));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i992_3_lut (.I0(n1454), .I1(n1507), 
            .I2(n1480), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i997_3_lut (.I0(n1459), .I1(n1512), 
            .I2(n1480), .I3(GND_net), .O(n1537));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1000_3_lut (.I0(n1462), .I1(n1515), 
            .I2(n1480), .I3(GND_net), .O(n1540));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i998_3_lut (.I0(n1460), .I1(n1513), 
            .I2(n1480), .I3(GND_net), .O(n1538));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i998_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1002_3_lut (.I0(n1464), .I1(n1517), 
            .I2(n1480), .I3(GND_net), .O(n1542));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1002_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i993_3_lut (.I0(n1455), .I1(n1508), 
            .I2(n1480), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1003_3_lut (.I0(n1465), .I1(n1518), 
            .I2(n1480), .I3(GND_net), .O(n1543));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1003_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i996_3_lut (.I0(n1458), .I1(n1511), 
            .I2(n1480), .I3(GND_net), .O(n1536));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i999_3_lut (.I0(n1461), .I1(n1514), 
            .I2(n1480), .I3(GND_net), .O(n1539));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1007_3_lut (.I0(n1469), .I1(n1522), 
            .I2(n1480), .I3(GND_net), .O(n1547));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1007_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1006_3_lut (.I0(n1468), .I1(n1521), 
            .I2(n1480), .I3(GND_net), .O(n1546));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1006_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3255_i7_3_lut (.I0(encoder0_position[6]), .I1(n19_adj_4886), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n526));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i940_3_lut (.I0(n1377), .I1(n1430), 
            .I2(n1402), .I3(GND_net), .O(n1455));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i940_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i947_3_lut (.I0(n1384), .I1(n1437), 
            .I2(n1402), .I3(GND_net), .O(n1462));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i947_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i950_3_lut (.I0(n1387), .I1(n1440), 
            .I2(n1402), .I3(GND_net), .O(n1465));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i950_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i942_3_lut (.I0(n1379), .I1(n1432), 
            .I2(n1402), .I3(GND_net), .O(n1457));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i942_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i943_3_lut (.I0(n1380), .I1(n1433), 
            .I2(n1402), .I3(GND_net), .O(n1458));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i943_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i939_3_lut (.I0(n1376), .I1(n1429), 
            .I2(n1402), .I3(GND_net), .O(n1454));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i939_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i944_3_lut (.I0(n1381), .I1(n1434), 
            .I2(n1402), .I3(GND_net), .O(n1459));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i944_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_1507__i31 (.Q(delay_counter[31]), .C(CLK_c), 
            .E(n21971), .D(n134), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 encoder0_position_23__I_0_i946_3_lut (.I0(n1383), .I1(n1436), 
            .I2(n1402), .I3(GND_net), .O(n1461));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i946_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i948_3_lut (.I0(n1385), .I1(n1438), 
            .I2(n1402), .I3(GND_net), .O(n1463));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i948_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i945_3_lut (.I0(n1382), .I1(n1435), 
            .I2(n1402), .I3(GND_net), .O(n1460));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i945_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i949_3_lut (.I0(n1386), .I1(n1439), 
            .I2(n1402), .I3(GND_net), .O(n1464));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i949_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i941_3_lut (.I0(n1378), .I1(n1431), 
            .I2(n1402), .I3(GND_net), .O(n1456));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i941_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i892_3_lut (.I0(n1304), .I1(n1357), 
            .I2(n1324), .I3(GND_net), .O(n1382));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i892_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i886_3_lut (.I0(n1298), .I1(n1351), 
            .I2(n1324), .I3(GND_net), .O(n1376));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i886_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i888_3_lut (.I0(n1300), .I1(n1353), 
            .I2(n1324), .I3(GND_net), .O(n1378));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i888_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i894_3_lut (.I0(n1306), .I1(n1359), 
            .I2(n1324), .I3(GND_net), .O(n1384));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i894_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i889_3_lut (.I0(n1301), .I1(n1354), 
            .I2(n1324), .I3(GND_net), .O(n1379));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i889_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i891_3_lut (.I0(n1303), .I1(n1356), 
            .I2(n1324), .I3(GND_net), .O(n1381));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i891_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i895_3_lut (.I0(n1307), .I1(n1360), 
            .I2(n1324), .I3(GND_net), .O(n1385));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i895_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i887_3_lut (.I0(n1299), .I1(n1352), 
            .I2(n1324), .I3(GND_net), .O(n1377));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i887_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i890_3_lut (.I0(n1302), .I1(n1355), 
            .I2(n1324), .I3(GND_net), .O(n1380));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i890_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i893_3_lut (.I0(n1305), .I1(n1358), 
            .I2(n1324), .I3(GND_net), .O(n1383));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i893_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i898_3_lut (.I0(n1310), .I1(n1363), 
            .I2(n1324), .I3(GND_net), .O(n1388));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i898_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14135_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n36883), .I3(GND_net), .O(n22538));   // verilog/coms.v(127[12] 300[6])
    defparam i14135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i896_3_lut (.I0(n1308), .I1(n1361), 
            .I2(n1324), .I3(GND_net), .O(n1386));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i896_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i897_3_lut (.I0(n1309), .I1(n1362), 
            .I2(n1324), .I3(GND_net), .O(n1387));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i897_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i837_3_lut (.I0(n1224), .I1(n1277), 
            .I2(n1246), .I3(GND_net), .O(n1302));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i840_3_lut (.I0(n1227), .I1(n1280), 
            .I2(n1246), .I3(GND_net), .O(n1305));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i839_3_lut (.I0(n1226), .I1(n1279), 
            .I2(n1246), .I3(GND_net), .O(n1304));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i834_3_lut (.I0(n1221), .I1(n1274), 
            .I2(n1246), .I3(GND_net), .O(n1299));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i834_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i836_3_lut (.I0(n1223), .I1(n1276), 
            .I2(n1246), .I3(GND_net), .O(n1301));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i835_3_lut (.I0(n1222), .I1(n1275), 
            .I2(n1246), .I3(GND_net), .O(n1300));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i835_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14136_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n36883), .I3(GND_net), .O(n22539));   // verilog/coms.v(127[12] 300[6])
    defparam i14136_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i838_3_lut (.I0(n1225), .I1(n1278), 
            .I2(n1246), .I3(GND_net), .O(n1303));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14137_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n36883), .I3(GND_net), .O(n22540));   // verilog/coms.v(127[12] 300[6])
    defparam i14137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i833_3_lut (.I0(n1220), .I1(n1273), 
            .I2(n1246), .I3(GND_net), .O(n1298));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i833_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i841_3_lut (.I0(n1228), .I1(n1281), 
            .I2(n1246), .I3(GND_net), .O(n1306));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14138_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n36883), .I3(GND_net), .O(n22541));   // verilog/coms.v(127[12] 300[6])
    defparam i14138_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i844_3_lut (.I0(n1231), .I1(n1284), 
            .I2(n1246), .I3(GND_net), .O(n1309));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i842_3_lut (.I0(n1229), .I1(n1282), 
            .I2(n1246), .I3(GND_net), .O(n1307));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i843_3_lut (.I0(n1230), .I1(n1283), 
            .I2(n1246), .I3(GND_net), .O(n1308));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i780_3_lut (.I0(n1142), .I1(n1195), 
            .I2(n1168), .I3(GND_net), .O(n1220));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i780_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14139_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n36883), .I3(GND_net), .O(n22542));   // verilog/coms.v(127[12] 300[6])
    defparam i14139_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14140_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n36883), .I3(GND_net), .O(n22543));   // verilog/coms.v(127[12] 300[6])
    defparam i14140_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i786_3_lut (.I0(n1148), .I1(n1201), 
            .I2(n1168), .I3(GND_net), .O(n1226));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i786_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i781_3_lut (.I0(n1143), .I1(n1196), 
            .I2(n1168), .I3(GND_net), .O(n1221));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i781_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i787_3_lut (.I0(n1149), .I1(n1202), 
            .I2(n1168), .I3(GND_net), .O(n1227));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i787_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14141_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n36883), .I3(GND_net), .O(n22544));   // verilog/coms.v(127[12] 300[6])
    defparam i14141_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i785_3_lut (.I0(n1147), .I1(n1200), 
            .I2(n1168), .I3(GND_net), .O(n1225));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i785_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i788_3_lut (.I0(n1150), .I1(n1203), 
            .I2(n1168), .I3(GND_net), .O(n1228));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i782_3_lut (.I0(n1144), .I1(n1197), 
            .I2(n1168), .I3(GND_net), .O(n1222));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i782_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i789_3_lut (.I0(n1151), .I1(n1204), 
            .I2(n1168), .I3(GND_net), .O(n1229));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i784_3_lut (.I0(n1146), .I1(n1199), 
            .I2(n1168), .I3(GND_net), .O(n1224));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14142_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n36883), .I3(GND_net), .O(n22545));   // verilog/coms.v(127[12] 300[6])
    defparam i14142_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i783_3_lut (.I0(n1145), .I1(n1198), 
            .I2(n1168), .I3(GND_net), .O(n1223));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i731_3_lut (.I0(n1068), .I1(n1121), 
            .I2(n1090), .I3(GND_net), .O(n1146));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i731_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i729_3_lut (.I0(n1066), .I1(n1119), 
            .I2(n1090), .I3(GND_net), .O(n1144));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i727_3_lut (.I0(n1064), .I1(n1117), 
            .I2(n1090), .I3(GND_net), .O(n1142));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i727_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i732_3_lut (.I0(n1069), .I1(n1122), 
            .I2(n1090), .I3(GND_net), .O(n1147));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i732_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14143_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n36883), .I3(GND_net), .O(n22546));   // verilog/coms.v(127[12] 300[6])
    defparam i14143_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i733_3_lut (.I0(n1070), .I1(n1123), 
            .I2(n1090), .I3(GND_net), .O(n1148));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i733_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i730_3_lut (.I0(n1067), .I1(n1120), 
            .I2(n1090), .I3(GND_net), .O(n1145));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i730_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_1507__i30 (.Q(delay_counter[30]), .C(CLK_c), 
            .E(n21971), .D(n135), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_DFFESR delay_counter_1507__i29 (.Q(delay_counter[29]), .C(CLK_c), 
            .E(n21971), .D(n136), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_DFFESR delay_counter_1507__i28 (.Q(delay_counter[28]), .C(CLK_c), 
            .E(n21971), .D(n137), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 i14144_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n36883), .I3(GND_net), .O(n22547));   // verilog/coms.v(127[12] 300[6])
    defparam i14144_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_1507__i27 (.Q(delay_counter[27]), .C(CLK_c), 
            .E(n21971), .D(n138), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 encoder0_position_23__I_0_i734_3_lut (.I0(n1071), .I1(n1124), 
            .I2(n1090), .I3(GND_net), .O(n1149));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i734_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i728_3_lut (.I0(n1065), .I1(n1118), 
            .I2(n1090), .I3(GND_net), .O(n1143));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i728_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i735_3_lut (.I0(n1072), .I1(n1125), 
            .I2(n1090), .I3(GND_net), .O(n1150));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i735_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i679_3_lut (.I0(n991), .I1(n1044), 
            .I2(n1012), .I3(GND_net), .O(n1069));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i679_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i676_3_lut (.I0(n988), .I1(n1041), 
            .I2(n1012), .I3(GND_net), .O(n1066));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i677_3_lut (.I0(n989), .I1(n1042), 
            .I2(n1012), .I3(GND_net), .O(n1067));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i677_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14145_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n36883), .I3(GND_net), .O(n22548));   // verilog/coms.v(127[12] 300[6])
    defparam i14145_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i682_3_lut (.I0(n994), .I1(n1047), 
            .I2(n1012), .I3(GND_net), .O(n1072));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i682_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_1507__i26 (.Q(delay_counter[26]), .C(CLK_c), 
            .E(n21971), .D(n139), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 encoder0_position_23__I_0_i680_3_lut (.I0(n992), .I1(n1045), 
            .I2(n1012), .I3(GND_net), .O(n1070));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i680_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_1507__i25 (.Q(delay_counter[25]), .C(CLK_c), 
            .E(n21971), .D(n140), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 encoder0_position_23__I_0_i681_3_lut (.I0(n993), .I1(n1046), 
            .I2(n1012), .I3(GND_net), .O(n1071));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i681_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14146_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n36883), .I3(GND_net), .O(n22549));   // verilog/coms.v(127[12] 300[6])
    defparam i14146_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i684_3_lut (.I0(n519), .I1(n1049), 
            .I2(n1012), .I3(GND_net), .O(n1074));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i684_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i683_3_lut (.I0(n995), .I1(n1048), 
            .I2(n1012), .I3(GND_net), .O(n1073));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i683_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i621_3_lut (.I0(n908), .I1(n961), 
            .I2(n934), .I3(GND_net), .O(n986));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i621_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14147_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n36883), .I3(GND_net), .O(n22550));   // verilog/coms.v(127[12] 300[6])
    defparam i14147_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i626_3_lut (.I0(n913), .I1(n966), 
            .I2(n934), .I3(GND_net), .O(n991));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i626_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i624_3_lut (.I0(n911), .I1(n964), 
            .I2(n934), .I3(GND_net), .O(n989));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i624_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i627_3_lut (.I0(n914), .I1(n967), 
            .I2(n934), .I3(GND_net), .O(n992));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i627_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i623_3_lut (.I0(n910), .I1(n963), 
            .I2(n934), .I3(GND_net), .O(n988));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i623_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i622_3_lut (.I0(n909), .I1(n962), 
            .I2(n934), .I3(GND_net), .O(n987));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i622_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_1507__i24 (.Q(delay_counter[24]), .C(CLK_c), 
            .E(n21971), .D(n141), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 encoder0_position_23__I_0_i570_3_lut (.I0(n832), .I1(n885), 
            .I2(n856), .I3(GND_net), .O(n910));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i570_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i569_3_lut (.I0(n831), .I1(n884), 
            .I2(n856), .I3(GND_net), .O(n909));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i569_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i571_3_lut (.I0(n833), .I1(n886), 
            .I2(n856), .I3(GND_net), .O(n911));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i571_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i572_3_lut (.I0(n834), .I1(n887), 
            .I2(n856), .I3(GND_net), .O(n912));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i572_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i568_3_lut (.I0(n830), .I1(n883), 
            .I2(n856), .I3(GND_net), .O(n908));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i568_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i573_3_lut (.I0(n835), .I1(n888), 
            .I2(n856), .I3(GND_net), .O(n913));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14148_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n36883), .I3(GND_net), .O(n22551));   // verilog/coms.v(127[12] 300[6])
    defparam i14148_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_1507__i23 (.Q(delay_counter[23]), .C(CLK_c), 
            .E(n21971), .D(n142), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 encoder0_position_23__I_0_i516_3_lut (.I0(n753), .I1(n806), 
            .I2(n778), .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i516_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i517_3_lut (.I0(n754), .I1(n807), 
            .I2(n778), .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i517_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i520_3_lut (.I0(n757), .I1(n810), 
            .I2(n778), .I3(GND_net), .O(n835));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i520_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14149_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n36883), .I3(GND_net), .O(n22552));   // verilog/coms.v(127[12] 300[6])
    defparam i14149_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i518_3_lut (.I0(n755), .I1(n808), 
            .I2(n778), .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i518_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i519_3_lut (.I0(n756), .I1(n809), 
            .I2(n778), .I3(GND_net), .O(n834));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i519_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i463_3_lut (.I0(n675), .I1(n728), 
            .I2(n700), .I3(GND_net), .O(n753));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i463_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i465_3_lut (.I0(n677), .I1(n730), 
            .I2(n700), .I3(GND_net), .O(n755));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i465_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14150_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n36883), .I3(GND_net), .O(n22553));   // verilog/coms.v(127[12] 300[6])
    defparam i14150_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14151_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n36883), .I3(GND_net), .O(n22554));   // verilog/coms.v(127[12] 300[6])
    defparam i14151_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3856_2_lut (.I0(n2), .I1(encoder0_position[23]), .I2(GND_net), 
            .I3(GND_net), .O(n509));
    defparam i3856_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26327_4_lut (.I0(encoder0_position[22]), .I1(n39289), .I2(encoder0_position[23]), 
            .I3(n3_adj_4904), .O(n675));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i26327_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i26325_3_lut (.I0(encoder0_position[21]), .I1(n36334), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n676));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i26325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3255_i19_3_lut (.I0(encoder0_position[18]), .I1(n7_adj_4898), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n514));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(n514), .I1(n6_adj_4899), .I2(GND_net), .I3(GND_net), 
            .O(n7_adj_4861));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(n4_adj_4903), .I1(n2), .I2(n5_adj_4900), .I3(n7_adj_4861), 
            .O(n4_adj_5000));
    defparam i1_4_lut.LUT_INIT = 16'hc888;
    SB_LUT4 i14152_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n36883), .I3(GND_net), .O(n22555));   // verilog/coms.v(127[12] 300[6])
    defparam i14152_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26357_3_lut (.I0(encoder0_position[19]), .I1(n36368), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n678));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i26357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14153_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n36883), .I3(GND_net), .O(n22556));   // verilog/coms.v(127[12] 300[6])
    defparam i14153_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26321_3_lut (.I0(encoder0_position[20]), .I1(n36330), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n677));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i26321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3255_i18_3_lut (.I0(encoder0_position[17]), .I1(n8_adj_4897), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n515));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19596_4_lut (.I0(n515), .I1(n677), .I2(n678), .I3(n679), 
            .O(n28004));
    defparam i19596_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i14154_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n36883), .I3(GND_net), .O(n22557));   // verilog/coms.v(127[12] 300[6])
    defparam i14154_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30272_4_lut (.I0(n676), .I1(n674), .I2(n675), .I3(n28004), 
            .O(n700));
    defparam i30272_4_lut.LUT_INIT = 16'h1333;
    SB_LUT4 i14155_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n36883), .I3(GND_net), .O(n22558));   // verilog/coms.v(127[12] 300[6])
    defparam i14155_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i26323_3_lut (.I0(encoder0_position[18]), .I1(n36332), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n679));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam i26323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i467_3_lut (.I0(n679), .I1(n732), 
            .I2(n700), .I3(GND_net), .O(n757));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i467_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i466_3_lut (.I0(n678), .I1(n731), 
            .I2(n700), .I3(GND_net), .O(n756));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i466_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i464_3_lut (.I0(n676), .I1(n729), 
            .I2(n700), .I3(GND_net), .O(n754));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i464_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i468_3_lut (.I0(n515), .I1(n733), 
            .I2(n700), .I3(GND_net), .O(n758));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i468_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19004_2_lut (.I0(n516), .I1(n758), .I2(GND_net), .I3(GND_net), 
            .O(n27400));
    defparam i19004_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1659 (.I0(n754), .I1(n27400), .I2(n756), .I3(n757), 
            .O(n4_adj_5011));
    defparam i1_4_lut_adj_1659.LUT_INIT = 16'ha8a0;
    SB_LUT4 i30335_4_lut (.I0(n752), .I1(n755), .I2(n753), .I3(n4_adj_5011), 
            .O(n778));
    defparam i30335_4_lut.LUT_INIT = 16'h0105;
    SB_LUT4 mux_3255_i17_3_lut (.I0(encoder0_position[16]), .I1(n9_adj_4896), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n516));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i522_3_lut (.I0(n516), .I1(n812), 
            .I2(n778), .I3(GND_net), .O(n837));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i521_3_lut (.I0(n758), .I1(n811), 
            .I2(n778), .I3(GND_net), .O(n836));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19426_3_lut (.I0(n517), .I1(n836), .I2(n837), .I3(GND_net), 
            .O(n27830));
    defparam i19426_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut (.I0(n834), .I1(n833), .I2(n27830), .I3(n835), 
            .O(n37256));
    defparam i2_4_lut.LUT_INIT = 16'h8880;
    SB_LUT4 i30348_4_lut (.I0(n37256), .I1(n830), .I2(n832), .I3(n831), 
            .O(n856));
    defparam i30348_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_3255_i16_3_lut (.I0(encoder0_position[15]), .I1(n10_adj_4895), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n517));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i576_3_lut (.I0(n517), .I1(n891), 
            .I2(n856), .I3(GND_net), .O(n916));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i575_3_lut (.I0(n837), .I1(n890), 
            .I2(n856), .I3(GND_net), .O(n915));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i575_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i574_3_lut (.I0(n836), .I1(n889), 
            .I2(n856), .I3(GND_net), .O(n914));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19582_4_lut (.I0(n518), .I1(n914), .I2(n915), .I3(n916), 
            .O(n27990));
    defparam i19582_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1660 (.I0(n913), .I1(n908), .I2(n912), .I3(n27990), 
            .O(n7_adj_4865));
    defparam i2_4_lut_adj_1660.LUT_INIT = 16'heccc;
    SB_LUT4 i30362_4_lut (.I0(n7_adj_4865), .I1(n911), .I2(n909), .I3(n910), 
            .O(n934));
    defparam i30362_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_3255_i15_3_lut (.I0(encoder0_position[14]), .I1(n11_adj_4894), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n518));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i630_3_lut (.I0(n518), .I1(n970), 
            .I2(n934), .I3(GND_net), .O(n995));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i630_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i629_3_lut (.I0(n916), .I1(n969), 
            .I2(n934), .I3(GND_net), .O(n994));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i629_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i628_3_lut (.I0(n915), .I1(n968), 
            .I2(n934), .I3(GND_net), .O(n993));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i628_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3255_i14_3_lut (.I0(encoder0_position[13]), .I1(n12_adj_4893), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n519));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19697_4_lut (.I0(n519), .I1(n993), .I2(n994), .I3(n995), 
            .O(n28106));
    defparam i19697_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_2_lut (.I0(n987), .I1(n988), .I2(GND_net), .I3(GND_net), 
            .O(n6_adj_5028));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1661 (.I0(n992), .I1(n989), .I2(n991), .I3(n28106), 
            .O(n5_adj_5029));
    defparam i1_4_lut_adj_1661.LUT_INIT = 16'heccc;
    SB_LUT4 i30377_4_lut (.I0(n986), .I1(n990), .I2(n5_adj_5029), .I3(n6_adj_5028), 
            .O(n1012));
    defparam i30377_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i625_3_lut (.I0(n912), .I1(n965), 
            .I2(n934), .I3(GND_net), .O(n990));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i625_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i678_3_lut (.I0(n990), .I1(n1043), 
            .I2(n1012), .I3(GND_net), .O(n1068));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i678_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i675_3_lut (.I0(n987), .I1(n1040), 
            .I2(n1012), .I3(GND_net), .O(n1065));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14156_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n36883), .I3(GND_net), .O(n22559));   // verilog/coms.v(127[12] 300[6])
    defparam i14156_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19578_3_lut (.I0(n520), .I1(n1073), .I2(n1074), .I3(GND_net), 
            .O(n27986));
    defparam i19578_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1662 (.I0(n1071), .I1(n1070), .I2(n27986), .I3(n1072), 
            .O(n36901));
    defparam i2_4_lut_adj_1662.LUT_INIT = 16'h8880;
    SB_LUT4 i5_4_lut (.I0(n1065), .I1(n1064), .I2(n36901), .I3(n1068), 
            .O(n12_adj_4860));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30297_4_lut (.I0(n1067), .I1(n12_adj_4860), .I2(n1066), .I3(n1069), 
            .O(n1090));
    defparam i30297_4_lut.LUT_INIT = 16'h0001;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_6 (.CI(n31796), 
            .I0(GND_net), .I1(n22_adj_4996), .CO(n31797));
    SB_LUT4 mux_3255_i13_3_lut (.I0(encoder0_position[12]), .I1(n13_adj_4892), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n520));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i738_3_lut (.I0(n520), .I1(n1128), 
            .I2(n1090), .I3(GND_net), .O(n1153));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i738_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i737_3_lut (.I0(n1074), .I1(n1127), 
            .I2(n1090), .I3(GND_net), .O(n1152));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i737_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i736_3_lut (.I0(n1073), .I1(n1126), 
            .I2(n1090), .I3(GND_net), .O(n1151));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i736_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19689_4_lut (.I0(n521), .I1(n1151), .I2(n1152), .I3(n1153), 
            .O(n28098));
    defparam i19689_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1663 (.I0(n1150), .I1(n1143), .I2(n1149), .I3(n28098), 
            .O(n5_adj_5022));
    defparam i1_4_lut_adj_1663.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1664 (.I0(n5_adj_5022), .I1(n1145), .I2(n1148), 
            .I3(n1147), .O(n6_adj_4872));
    defparam i1_4_lut_adj_1664.LUT_INIT = 16'hfffe;
    SB_LUT4 i30323_4_lut (.I0(n1142), .I1(n1144), .I2(n1146), .I3(n6_adj_4872), 
            .O(n1168));
    defparam i30323_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_3255_i12_3_lut (.I0(encoder0_position[11]), .I1(n14_adj_4891), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n521));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i792_3_lut (.I0(n521), .I1(n1207), 
            .I2(n1168), .I3(GND_net), .O(n1232));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i792_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i791_3_lut (.I0(n1153), .I1(n1206), 
            .I2(n1168), .I3(GND_net), .O(n1231));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1494_3_lut (.I0(n2026), .I1(n5700), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[1]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1494_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i790_3_lut (.I0(n1152), .I1(n1205), 
            .I2(n1168), .I3(GND_net), .O(n1230));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i790_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19685_4_lut (.I0(n522), .I1(n1230), .I2(n1231), .I3(n1232), 
            .O(n28094));
    defparam i19685_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_adj_1665 (.I0(n1223), .I1(n1224), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_5014));
    defparam i1_2_lut_adj_1665.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(n1229), .I1(n1222), .I2(n1228), .I3(n28094), 
            .O(n12_adj_5013));
    defparam i3_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i7_4_lut (.I0(n1225), .I1(n1227), .I2(n1221), .I3(n10_adj_5014), 
            .O(n16_adj_5012));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30455_4_lut (.I0(n1226), .I1(n16_adj_5012), .I2(n12_adj_5013), 
            .I3(n1220), .O(n1246));
    defparam i30455_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1493_3_lut (.I0(n1948), .I1(n5699), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[2]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1493_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1492_3_lut (.I0(n1870), .I1(n5698), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[3]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1492_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 mux_3255_i11_3_lut (.I0(encoder0_position[10]), .I1(n15_adj_4890), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n522));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i846_3_lut (.I0(n522), .I1(n1286), 
            .I2(n1246), .I3(GND_net), .O(n1311));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1491_3_lut (.I0(n1792), .I1(n5697), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[4]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1491_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1490_3_lut (.I0(n1714), .I1(n5696), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[5]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1490_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1489_3_lut (.I0(n1636), .I1(n5695), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[6]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1489_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i845_3_lut (.I0(n1232), .I1(n1285), 
            .I2(n1246), .I3(GND_net), .O(n1310));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1488_3_lut (.I0(n1558), .I1(n5694), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[7]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1488_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 unary_minus_4_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19567_3_lut (.I0(n523), .I1(n1310), .I2(n1311), .I3(GND_net), 
            .O(n27974));
    defparam i19567_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1666 (.I0(n1308), .I1(n1307), .I2(n27974), .I3(n1309), 
            .O(n37465));
    defparam i2_4_lut_adj_1666.LUT_INIT = 16'h8880;
    SB_LUT4 i4_4_lut (.I0(n1306), .I1(n1298), .I2(n37465), .I3(n1303), 
            .O(n10_adj_5023));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1667 (.I0(n1300), .I1(n1301), .I2(n10_adj_5023), 
            .I3(n1299), .O(n6_adj_5001));
    defparam i1_4_lut_adj_1667.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_i1487_3_lut (.I0(n1480), .I1(n5693), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[8]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1487_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i30527_4_lut (.I0(n1304), .I1(n1305), .I2(n1302), .I3(n6_adj_5001), 
            .O(n1324));
    defparam i30527_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_3255_i10_3_lut (.I0(encoder0_position[9]), .I1(n16_adj_4889), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n523));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i900_3_lut (.I0(n523), .I1(n1365), 
            .I2(n1324), .I3(GND_net), .O(n1390));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i900_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1486_3_lut (.I0(n1402), .I1(n5692), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[9]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1486_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i899_3_lut (.I0(n1311), .I1(n1364), 
            .I2(n1324), .I3(GND_net), .O(n1389));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i899_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19563_3_lut (.I0(n524), .I1(n1389), .I2(n1390), .I3(GND_net), 
            .O(n27970));
    defparam i19563_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_23__I_0_i1485_3_lut (.I0(n1324), .I1(n5691), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[10]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1485_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i2_4_lut_adj_1668 (.I0(n1387), .I1(n1386), .I2(n27970), .I3(n1388), 
            .O(n37487));
    defparam i2_4_lut_adj_1668.LUT_INIT = 16'h8880;
    SB_LUT4 i7_4_lut_adj_1669 (.I0(n1383), .I1(n1380), .I2(n1377), .I3(n37487), 
            .O(n18_adj_4863));
    defparam i7_4_lut_adj_1669.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut (.I0(n1385), .I1(n1381), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4864));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_23__I_0_i1484_3_lut (.I0(n1246), .I1(n5690), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[11]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1484_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1483_3_lut (.I0(n1168), .I1(n5689), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[12]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1483_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i9_4_lut (.I0(n1379), .I1(n18_adj_4863), .I2(n1384), .I3(n1378), 
            .O(n20_adj_4862));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30577_4_lut (.I0(n1376), .I1(n20_adj_4862), .I2(n16_adj_4864), 
            .I3(n1382), .O(n1402));
    defparam i30577_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1482_3_lut (.I0(n1090), .I1(n5688), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[13]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1482_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 mux_3255_i9_3_lut (.I0(encoder0_position[8]), .I1(n17_adj_4888), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n524));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1481_3_lut (.I0(n1012), .I1(n5687), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[14]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1481_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i954_3_lut (.I0(n524), .I1(n1444), 
            .I2(n1402), .I3(GND_net), .O(n1469));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i954_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i953_3_lut (.I0(n1390), .I1(n1443), 
            .I2(n1402), .I3(GND_net), .O(n1468));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i953_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i952_3_lut (.I0(n1389), .I1(n1442), 
            .I2(n1402), .I3(GND_net), .O(n1467));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i952_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3255_i8_3_lut (.I0(encoder0_position[7]), .I1(n18_adj_4887), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n525));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19669_4_lut (.I0(n525), .I1(n1467), .I2(n1468), .I3(n1469), 
            .O(n28078));
    defparam i19669_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i8_4_lut (.I0(n1456), .I1(n1464), .I2(n1460), .I3(n1463), 
            .O(n20_adj_4910));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1670 (.I0(n1457), .I1(n1466), .I2(n1465), .I3(n28078), 
            .O(n13_adj_4913));
    defparam i1_4_lut_adj_1670.LUT_INIT = 16'heaaa;
    SB_LUT4 i6_2_lut (.I0(n1461), .I1(n1459), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4911));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut (.I0(n13_adj_4913), .I1(n20_adj_4910), .I2(n1454), 
            .I3(n1458), .O(n22_adj_4909));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14157_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n36883), .I3(GND_net), .O(n22560));   // verilog/coms.v(127[12] 300[6])
    defparam i14157_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30146_4_lut (.I0(n1462), .I1(n22_adj_4909), .I2(n18_adj_4911), 
            .I3(n1455), .O(n1480));
    defparam i30146_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1480_3_lut (.I0(n934), .I1(n5686), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[15]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1480_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i951_3_lut (.I0(n1388), .I1(n1441), 
            .I2(n1402), .I3(GND_net), .O(n1466));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i951_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1479_3_lut (.I0(n856), .I1(n5685), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[16]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1479_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 encoder0_position_23__I_0_i1004_3_lut (.I0(n1466), .I1(n1519), 
            .I2(n1480), .I3(GND_net), .O(n1544));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1004_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i994_3_lut (.I0(n1456), .I1(n1509), 
            .I2(n1480), .I3(GND_net), .O(n1534));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1005_3_lut (.I0(n1467), .I1(n1520), 
            .I2(n1480), .I3(GND_net), .O(n1545));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1005_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14158_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n18082), .I3(GND_net), .O(n22561));   // verilog/coms.v(127[12] 300[6])
    defparam i14158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1478_3_lut (.I0(n778), .I1(n5684), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[17]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1478_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i19663_4_lut (.I0(n526), .I1(n1546), .I2(n1547), .I3(n1548), 
            .O(n28072));
    defparam i19663_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i4_4_lut_adj_1671 (.I0(n1545), .I1(n1534), .I2(n1544), .I3(n28072), 
            .O(n17_adj_4876));
    defparam i4_4_lut_adj_1671.LUT_INIT = 16'heccc;
    SB_LUT4 i8_4_lut_adj_1672 (.I0(n1533), .I1(n1542), .I2(n1538), .I3(n1540), 
            .O(n21_adj_4874));
    defparam i8_4_lut_adj_1672.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(n1539), .I1(n1536), .I2(n1543), .I3(GND_net), 
            .O(n20_adj_4875));
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut (.I0(n21_adj_4874), .I1(n17_adj_4876), .I2(n1537), 
            .I3(n1532), .O(n24_adj_4873));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30180_4_lut (.I0(n1535), .I1(n24_adj_4873), .I2(n20_adj_4875), 
            .I3(n1541), .O(n1558));
    defparam i30180_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1008_3_lut (.I0(n525), .I1(n1523), 
            .I2(n1480), .I3(GND_net), .O(n1548));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1008_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1061_3_lut (.I0(n1548), .I1(n1601), 
            .I2(n1558), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3255_i6_3_lut (.I0(encoder0_position[5]), .I1(n20_adj_4885), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n527));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19537_3_lut (.I0(n527), .I1(n1626), .I2(n1627), .I3(GND_net), 
            .O(n27944));
    defparam i19537_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1673 (.I0(n1624), .I1(n1623), .I2(n27944), .I3(n1625), 
            .O(n37470));
    defparam i2_4_lut_adj_1673.LUT_INIT = 16'h8880;
    SB_LUT4 i4_2_lut (.I0(n1611), .I1(n1618), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_5009));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1674 (.I0(n1614), .I1(n1612), .I2(n1617), .I3(n1615), 
            .O(n24_adj_5007));
    defparam i10_4_lut_adj_1674.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1675 (.I0(n1610), .I1(n1622), .I2(n1620), .I3(n37470), 
            .O(n22_adj_5008));
    defparam i8_4_lut_adj_1675.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n1616), .I1(n24_adj_5007), .I2(n18_adj_5009), 
            .I3(n1613), .O(n26_adj_5006));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30205_4_lut (.I0(n1621), .I1(n26_adj_5006), .I2(n22_adj_5008), 
            .I3(n1619), .O(n1636));
    defparam i30205_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1062_3_lut (.I0(n526), .I1(n1602), 
            .I2(n1558), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1115_3_lut (.I0(n1627), .I1(n1680), 
            .I2(n1636), .I3(GND_net), .O(n1705));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3255_i5_3_lut (.I0(encoder0_position[4]), .I1(n21_adj_4884), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n528));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19535_3_lut (.I0(n528), .I1(n1705), .I2(n1706), .I3(GND_net), 
            .O(n27942));
    defparam i19535_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1676 (.I0(n1703), .I1(n1702), .I2(n27942), .I3(n1704), 
            .O(n37237));
    defparam i2_4_lut_adj_1676.LUT_INIT = 16'h8880;
    SB_LUT4 i5_4_lut_adj_1677 (.I0(n37237), .I1(n1695), .I2(n1700), .I3(n1699), 
            .O(n12_adj_5018));
    defparam i5_4_lut_adj_1677.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_i1477_3_lut (.I0(n700), .I1(n5683), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[18]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1477_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i4_3_lut (.I0(n1701), .I1(n1698), .I2(n1691), .I3(GND_net), 
            .O(n11_adj_5019));
    defparam i4_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_4_lut_adj_1678 (.I0(n1688), .I1(n11_adj_5019), .I2(n1693), 
            .I3(n12_adj_5018), .O(n14_adj_4867));
    defparam i5_4_lut_adj_1678.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(n1697), .I1(n1690), .I2(n1694), .I3(n1696), 
            .O(n15_adj_4866));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30483_4_lut (.I0(n15_adj_4866), .I1(n1689), .I2(n14_adj_4867), 
            .I3(n1692), .O(n1714));
    defparam i30483_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1116_3_lut (.I0(n527), .I1(n1681), 
            .I2(n1636), .I3(GND_net), .O(n1706));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1169_3_lut (.I0(n1706), .I1(n1759), 
            .I2(n1714), .I3(GND_net), .O(n1784));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1169_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3255_i4_3_lut (.I0(encoder0_position[3]), .I1(n22_adj_4883), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n529));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19531_3_lut (.I0(n529), .I1(n1784), .I2(n1785), .I3(GND_net), 
            .O(n27938));
    defparam i19531_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_4_lut_adj_1679 (.I0(n1782), .I1(n1781), .I2(n27938), .I3(n1783), 
            .O(n37463));
    defparam i2_4_lut_adj_1679.LUT_INIT = 16'h8880;
    SB_LUT4 i12_4_lut_adj_1680 (.I0(n1772), .I1(n1767), .I2(n1775), .I3(n1779), 
            .O(n28_adj_4973));
    defparam i12_4_lut_adj_1680.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1681 (.I0(n1770), .I1(n1773), .I2(n1766), .I3(n1771), 
            .O(n26));
    defparam i10_4_lut_adj_1681.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1682 (.I0(n1778), .I1(n1777), .I2(n1774), .I3(n1768), 
            .O(n27_adj_4974));
    defparam i11_4_lut_adj_1682.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1683 (.I0(n37463), .I1(n1776), .I2(n1769), .I3(n1780), 
            .O(n25_adj_4975));
    defparam i9_4_lut_adj_1683.LUT_INIT = 16'hfffe;
    SB_LUT4 i30508_4_lut (.I0(n25_adj_4975), .I1(n27_adj_4974), .I2(n26), 
            .I3(n28_adj_4973), .O(n1792));
    defparam i30508_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1170_3_lut (.I0(n528), .I1(n1760), 
            .I2(n1714), .I3(GND_net), .O(n1785));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1170_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1224_3_lut (.I0(n529), .I1(n1839), 
            .I2(n1792), .I3(GND_net), .O(n1864));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1224_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1223_3_lut (.I0(n1785), .I1(n1838), 
            .I2(n1792), .I3(GND_net), .O(n1863));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1223_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1222_3_lut (.I0(n1784), .I1(n1837), 
            .I2(n1792), .I3(GND_net), .O(n1862));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1222_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3255_i3_3_lut (.I0(encoder0_position[2]), .I1(n23_adj_4882), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n530));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19645_4_lut (.I0(n530), .I1(n1862), .I2(n1863), .I3(n1864), 
            .O(n28054));
    defparam i19645_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1684 (.I0(n1858), .I1(n1861), .I2(n1860), .I3(n28054), 
            .O(n4_adj_5024));
    defparam i1_4_lut_adj_1684.LUT_INIT = 16'heaaa;
    SB_LUT4 i3_2_lut (.I0(n1846), .I1(n1856), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_4871));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut_adj_1685 (.I0(n1859), .I1(n10_adj_4871), .I2(n1857), 
            .I3(n4_adj_5024), .O(n12_adj_4869));
    defparam i5_4_lut_adj_1685.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_4_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_3_lut_adj_1686 (.I0(n1850), .I1(n1848), .I2(n1854), .I3(GND_net), 
            .O(n11_adj_4870));
    defparam i4_3_lut_adj_1686.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_4_lut_adj_1687 (.I0(n1847), .I1(n1851), .I2(n11_adj_4870), 
            .I3(n12_adj_4869), .O(n14_adj_5027));
    defparam i5_4_lut_adj_1687.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1688 (.I0(n1855), .I1(n1853), .I2(n1852), .I3(n1845), 
            .O(n15_adj_5026));
    defparam i6_4_lut_adj_1688.LUT_INIT = 16'hfffe;
    SB_LUT4 i30556_4_lut (.I0(n15_adj_5026), .I1(n1849), .I2(n14_adj_5027), 
            .I3(n1844), .O(n1870));
    defparam i30556_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1214_3_lut (.I0(n1776), .I1(n1829), 
            .I2(n1792), .I3(GND_net), .O(n1854));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1214_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1267_3_lut (.I0(n1854), .I1(n1907), 
            .I2(n1870), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1267_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1272_3_lut (.I0(n1859), .I1(n1912), 
            .I2(n1870), .I3(GND_net), .O(n1937));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1272_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1273_3_lut (.I0(n1860), .I1(n1913), 
            .I2(n1870), .I3(GND_net), .O(n1938));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1273_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1260_3_lut (.I0(n1847), .I1(n1900), 
            .I2(n1870), .I3(GND_net), .O(n1925));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1260_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i10_4_lut_adj_1689 (.I0(n1925), .I1(n1938), .I2(n1937), .I3(n1932), 
            .O(n28));
    defparam i10_4_lut_adj_1689.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(n1926), .I1(n1933), .I2(n1929), .I3(n1924), 
            .O(n31_adj_4951));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19641_4_lut (.I0(n531), .I1(n1941), .I2(n1942), .I3(n1943), 
            .O(n28050));
    defparam i19641_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i4_2_lut_adj_1690 (.I0(n1928), .I1(n1935), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4953));
    defparam i4_2_lut_adj_1690.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1691 (.I0(n1931), .I1(n1930), .I2(n1922), .I3(n1936), 
            .O(n30_adj_4952));
    defparam i12_4_lut_adj_1691.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n31_adj_4951), .I1(n1927), .I2(n28), .I3(n1923), 
            .O(n34_adj_4950));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14159_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n18082), .I3(GND_net), .O(n22562));   // verilog/coms.v(127[12] 300[6])
    defparam i14159_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1692 (.I0(n1940), .I1(n1934), .I2(n1939), .I3(n28050), 
            .O(n21_adj_4954));
    defparam i3_4_lut_adj_1692.LUT_INIT = 16'heccc;
    SB_LUT4 i30404_4_lut (.I0(n21_adj_4954), .I1(n34_adj_4950), .I2(n30_adj_4952), 
            .I3(n22_adj_4953), .O(n1948));
    defparam i30404_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_23__I_0_i1257_3_lut (.I0(n1844), .I1(n1897), 
            .I2(n1870), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1257_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1310_3_lut (.I0(n1922), .I1(n1975), 
            .I2(n1948), .I3(GND_net), .O(n2000));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i13_1_lut (.I0(encoder0_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4932));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13889_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n21865), .I3(GND_net), .O(n22292));   // verilog/coms.v(127[12] 300[6])
    defparam i13889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14160_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n18082), .I3(GND_net), .O(n22563));   // verilog/coms.v(127[12] 300[6])
    defparam i14160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14161_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n18082), .I3(GND_net), .O(n22564));   // verilog/coms.v(127[12] 300[6])
    defparam i14161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14162_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n18082), .I3(GND_net), .O(n22565));   // verilog/coms.v(127[12] 300[6])
    defparam i14162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14163_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n18082), .I3(GND_net), .O(n22566));   // verilog/coms.v(127[12] 300[6])
    defparam i14163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_65_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[10]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_65_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[11]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14164_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n18082), .I3(GND_net), .O(n22567));   // verilog/coms.v(127[12] 300[6])
    defparam i14164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i14_1_lut (.I0(encoder0_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4931));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14165_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n18082), .I3(GND_net), .O(n22568));   // verilog/coms.v(127[12] 300[6])
    defparam i14165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_65_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[12]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14166_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n18082), .I3(GND_net), .O(n22569));   // verilog/coms.v(127[12] 300[6])
    defparam i14166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_65_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[13]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14167_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n18082), .I3(GND_net), .O(n22570));   // verilog/coms.v(127[12] 300[6])
    defparam i14167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i15_1_lut (.I0(encoder0_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4930));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14168_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n18082), .I3(GND_net), .O(n22571));   // verilog/coms.v(127[12] 300[6])
    defparam i14168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_65_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[14]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14169_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n18082), .I3(GND_net), .O(n22572));   // verilog/coms.v(127[12] 300[6])
    defparam i14169_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_4997), .I3(n31795), .O(n23_adj_4882)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14170_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n18082), .I3(GND_net), .O(n22573));   // verilog/coms.v(127[12] 300[6])
    defparam i14170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14171_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n18082), .I3(GND_net), .O(n22574));   // verilog/coms.v(127[12] 300[6])
    defparam i14171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14172_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n18082), .I3(GND_net), .O(n22575));   // verilog/coms.v(127[12] 300[6])
    defparam i14172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i16_1_lut (.I0(encoder0_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4929));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14173_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n18082), .I3(GND_net), .O(n22576));   // verilog/coms.v(127[12] 300[6])
    defparam i14173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14174_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n18082), .I3(GND_net), .O(n22577));   // verilog/coms.v(127[12] 300[6])
    defparam i14174_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14175_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n18082), .I3(GND_net), .O(n22578));   // verilog/coms.v(127[12] 300[6])
    defparam i14175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14176_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n18082), .I3(GND_net), .O(n22579));   // verilog/coms.v(127[12] 300[6])
    defparam i14176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14177_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n18082), .I3(GND_net), .O(n22580));   // verilog/coms.v(127[12] 300[6])
    defparam i14177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14178_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n18082), .I3(GND_net), .O(n22581));   // verilog/coms.v(127[12] 300[6])
    defparam i14178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14179_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n18082), .I3(GND_net), .O(n22582));   // verilog/coms.v(127[12] 300[6])
    defparam i14179_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1373_3_lut (.I0(n2010), .I1(n2063), 
            .I2(n2026), .I3(GND_net), .O(n29_adj_5005));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14180_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n18082), .I3(GND_net), .O(n22583));   // verilog/coms.v(127[12] 300[6])
    defparam i14180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1374_3_lut (.I0(n2011), .I1(n2064), 
            .I2(n2026), .I3(GND_net), .O(n27_adj_5004));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1365_3_lut (.I0(n2002), .I1(n2055), 
            .I2(n2026), .I3(GND_net), .O(n45));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1365_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14181_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n18082), .I3(GND_net), .O(n22584));   // verilog/coms.v(127[12] 300[6])
    defparam i14181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1381_3_lut (.I0(n2018), .I1(n2071), 
            .I2(n2026), .I3(GND_net), .O(n13_adj_5002));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14182_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n18082), .I3(GND_net), .O(n22585));   // verilog/coms.v(127[12] 300[6])
    defparam i14182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14183_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n18082), .I3(GND_net), .O(n22586));   // verilog/coms.v(127[12] 300[6])
    defparam i14183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_65_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[15]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_i1368_3_lut (.I0(n2005), .I1(n2058), 
            .I2(n2026), .I3(GND_net), .O(n39));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1368_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16_4_lut_adj_1693 (.I0(n2020), .I1(n39214), .I2(n2026), .I3(n2019), 
            .O(n5_adj_4946));
    defparam i16_4_lut_adj_1693.LUT_INIT = 16'hac0c;
    SB_LUT4 i29535_3_lut (.I0(n532), .I1(n2021), .I2(n2022), .I3(GND_net), 
            .O(n39271));
    defparam i29535_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mux_65_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[16]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_23__I_0_i1363_3_lut (.I0(n2000), .I1(n2053), 
            .I2(n2026), .I3(GND_net), .O(n49));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1363_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1366_3_lut (.I0(n2003), .I1(n2056), 
            .I2(n2026), .I3(GND_net), .O(n43));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1366_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1694 (.I0(n39271), .I1(n5_adj_4946), .I2(n39272), 
            .I3(n2026), .O(n34038));
    defparam i1_4_lut_adj_1694.LUT_INIT = 16'h88c0;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i17_1_lut (.I0(encoder0_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4928));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29541_2_lut (.I0(start), .I1(n14), .I2(GND_net), .I3(GND_net), 
            .O(n39198));   // verilog/neopixel.v(35[12] 117[6])
    defparam i29541_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i4_4_lut_adj_1695 (.I0(n2016), .I1(n29_adj_5005), .I2(n2069), 
            .I3(n2026), .O(n24_adj_5037));
    defparam i4_4_lut_adj_1695.LUT_INIT = 16'heefc;
    SB_LUT4 i2_4_lut_adj_1696 (.I0(n34038), .I1(n2001), .I2(n2054), .I3(n2026), 
            .O(n22_adj_5039));
    defparam i2_4_lut_adj_1696.LUT_INIT = 16'heefa;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i18_1_lut (.I0(encoder0_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4927));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i19_1_lut (.I0(encoder0_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4926));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_4_lut_adj_1697 (.I0(n2007), .I1(n49), .I2(n2060), .I3(n2026), 
            .O(n23_adj_5038));
    defparam i3_4_lut_adj_1697.LUT_INIT = 16'heefc;
    SB_LUT4 i31_4_lut (.I0(n39198), .I1(n39196), .I2(state[1]), .I3(\neo_pixel_transmitter.done ), 
            .O(n34460));   // verilog/neopixel.v(35[12] 117[6])
    defparam i31_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i1_4_lut_adj_1698 (.I0(n2014), .I1(n43), .I2(n2067), .I3(n2026), 
            .O(n21_adj_5040));
    defparam i1_4_lut_adj_1698.LUT_INIT = 16'heefc;
    SB_LUT4 i13891_4_lut (.I0(state_7__N_3881[3]), .I1(data[7]), .I2(n27086), 
            .I3(n20731), .O(n22294));   // verilog/i2c_controller.v(89[8] 155[6])
    defparam i13891_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_23__I_0_i1369_3_lut (.I0(n2006), .I1(n2059), 
            .I2(n2026), .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1369_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13892_4_lut (.I0(state_7__N_3881[3]), .I1(data[6]), .I2(n27086), 
            .I3(n20726), .O(n22295));   // verilog/i2c_controller.v(89[8] 155[6])
    defparam i13892_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_23__I_0_i1376_3_lut (.I0(n2013), .I1(n2066), 
            .I2(n2026), .I3(GND_net), .O(n23_adj_5003));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13893_4_lut (.I0(state_7__N_3881[3]), .I1(data[5]), .I2(n4_adj_4945), 
            .I3(n20731), .O(n22296));   // verilog/i2c_controller.v(89[8] 155[6])
    defparam i13893_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i8_4_lut_adj_1699 (.I0(n2008), .I1(n27_adj_5004), .I2(n2061), 
            .I3(n2026), .O(n28_adj_5033));
    defparam i8_4_lut_adj_1699.LUT_INIT = 16'heefc;
    SB_LUT4 i6_4_lut_adj_1700 (.I0(n2004), .I1(n45), .I2(n2057), .I3(n2026), 
            .O(n26_adj_5035));
    defparam i6_4_lut_adj_1700.LUT_INIT = 16'heefc;
    SB_LUT4 i7_4_lut_adj_1701 (.I0(n2012), .I1(n13_adj_5002), .I2(n2065), 
            .I3(n2026), .O(n27_adj_5034));
    defparam i7_4_lut_adj_1701.LUT_INIT = 16'heefc;
    SB_LUT4 mux_65_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[17]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i5_4_lut_adj_1702 (.I0(n2017), .I1(n23_adj_5003), .I2(n2070), 
            .I3(n2026), .O(n25_adj_5036));
    defparam i5_4_lut_adj_1702.LUT_INIT = 16'heefc;
    SB_LUT4 i10_4_lut_adj_1703 (.I0(n2009), .I1(n39), .I2(n2062), .I3(n2026), 
            .O(n30_adj_5031));
    defparam i10_4_lut_adj_1703.LUT_INIT = 16'heefc;
    SB_LUT4 i16_4_lut_adj_1704 (.I0(n21_adj_5040), .I1(n23_adj_5038), .I2(n22_adj_5039), 
            .I3(n24_adj_5037), .O(n36));
    defparam i16_4_lut_adj_1704.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1705 (.I0(n2015), .I1(n37), .I2(n2068), .I3(n2026), 
            .O(n29_adj_5032));
    defparam i9_4_lut_adj_1705.LUT_INIT = 16'heefc;
    SB_LUT4 i17_4_lut (.I0(n25_adj_5036), .I1(n27_adj_5034), .I2(n26_adj_5035), 
            .I3(n28_adj_5033), .O(n37_adj_5030));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13894_4_lut (.I0(state_7__N_3881[3]), .I1(data[4]), .I2(n4_adj_4945), 
            .I3(n20726), .O(n22297));   // verilog/i2c_controller.v(89[8] 155[6])
    defparam i13894_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30433_4_lut (.I0(n37_adj_5030), .I1(n29_adj_5032), .I2(n36), 
            .I3(n30_adj_5031), .O(n28040));
    defparam i30433_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i13895_4_lut (.I0(state_7__N_3881[3]), .I1(data[3]), .I2(n4_adj_4877), 
            .I3(n20731), .O(n22298));   // verilog/i2c_controller.v(89[8] 155[6])
    defparam i13895_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i20_1_lut (.I0(encoder0_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4925));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13896_4_lut (.I0(state_7__N_3881[3]), .I1(data[2]), .I2(n4_adj_4877), 
            .I3(n20726), .O(n22299));   // verilog/i2c_controller.v(89[8] 155[6])
    defparam i13896_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_65_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[18]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13897_4_lut (.I0(state_7__N_3881[3]), .I1(data[1]), .I2(n10_adj_5010), 
            .I3(n20731), .O(n22300));   // verilog/i2c_controller.v(89[8] 155[6])
    defparam i13897_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14184_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n18082), .I3(GND_net), .O(n22587));   // verilog/coms.v(127[12] 300[6])
    defparam i14184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14185_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n18082), .I3(GND_net), .O(n22588));   // verilog/coms.v(127[12] 300[6])
    defparam i14185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1706 (.I0(n2002), .I1(n2011), .I2(n2008), .I3(n2001), 
            .O(n30));
    defparam i11_4_lut_adj_1706.LUT_INIT = 16'hfffe;
    SB_LUT4 i19519_3_lut (.I0(n532), .I1(n2021), .I2(n2022), .I3(GND_net), 
            .O(n27926));
    defparam i19519_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i14186_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n18082), .I3(GND_net), .O(n22589));   // verilog/coms.v(127[12] 300[6])
    defparam i14186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14187_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n18082), .I3(GND_net), .O(n22590));   // verilog/coms.v(127[12] 300[6])
    defparam i14187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1707 (.I0(n2019), .I1(n2018), .I2(n27926), .I3(n2020), 
            .O(n37048));
    defparam i2_4_lut_adj_1707.LUT_INIT = 16'h8880;
    SB_LUT4 i15_4_lut (.I0(n2003), .I1(n30), .I2(n2015), .I3(n2014), 
            .O(n34));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14188_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n18082), .I3(GND_net), .O(n22591));   // verilog/coms.v(127[12] 300[6])
    defparam i14188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14189_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n18082), .I3(GND_net), .O(n22592));   // verilog/coms.v(127[12] 300[6])
    defparam i14189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14190_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n18082), .I3(GND_net), .O(n22593));   // verilog/coms.v(127[12] 300[6])
    defparam i14190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_4_lut_adj_1708 (.I0(n2000), .I1(n2016), .I2(n2010), .I3(n2006), 
            .O(n32));
    defparam i13_4_lut_adj_1708.LUT_INIT = 16'hfffe;
    SB_DFFESR delay_counter_1507__i22 (.Q(delay_counter[22]), .C(CLK_c), 
            .E(n21971), .D(n143), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_5 (.CI(n31795), 
            .I0(GND_net), .I1(n23_adj_4997), .CO(n31796));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_4998), .I3(n31794), .O(n24_adj_4881)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_4 (.CI(n31794), 
            .I0(GND_net), .I1(n24_adj_4998), .CO(n31795));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_4999), .I3(n31793), .O(n25_adj_4880)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14_4_lut (.I0(n2009), .I1(n2004), .I2(n2013), .I3(n2007), 
            .O(n33));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1709 (.I0(n2017), .I1(n2005), .I2(n2012), .I3(n37048), 
            .O(n31));
    defparam i12_4_lut_adj_1709.LUT_INIT = 16'hfffe;
    SB_LUT4 i30429_4_lut (.I0(n31), .I1(n33), .I2(n32), .I3(n34), .O(n2026));
    defparam i30429_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i13899_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n26980), 
            .I3(n20781), .O(n22302));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13899_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4976));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i21_1_lut (.I0(encoder0_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4924));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_65_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[19]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13900_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n26980), 
            .I3(n20776), .O(n22303));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13900_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 mux_65_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[20]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13901_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_4921), 
            .I3(n20781), .O(n22304));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13901_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13902_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_4921), 
            .I3(n20776), .O(n22305));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13902_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_4_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13903_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_4920), 
            .I3(n20781), .O(n22306));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13903_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 mux_65_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[21]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13904_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_4920), 
            .I3(n20776), .O(n22307));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13904_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14191_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n18082), .I3(GND_net), .O(n22594));   // verilog/coms.v(127[12] 300[6])
    defparam i14191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14192_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n18082), .I3(GND_net), .O(n22595));   // verilog/coms.v(127[12] 300[6])
    defparam i14192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i23_1_lut (.I0(encoder0_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4923));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14193_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n18082), .I3(GND_net), .O(n22596));   // verilog/coms.v(127[12] 300[6])
    defparam i14193_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_1507__i21 (.Q(delay_counter[21]), .C(CLK_c), 
            .E(n21971), .D(n144), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 mux_65_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[22]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14194_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n18082), .I3(GND_net), .O(n22597));   // verilog/coms.v(127[12] 300[6])
    defparam i14194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14195_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n18082), .I3(GND_net), .O(n22598));   // verilog/coms.v(127[12] 300[6])
    defparam i14195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14196_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n18082), .I3(GND_net), .O(n22599));   // verilog/coms.v(127[12] 300[6])
    defparam i14196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14197_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n18082), .I3(GND_net), .O(n22600));   // verilog/coms.v(127[12] 300[6])
    defparam i14197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14198_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n18082), .I3(GND_net), .O(n22601));   // verilog/coms.v(127[12] 300[6])
    defparam i14198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1710 (.I0(control_mode[3]), .I1(control_mode[5]), 
            .I2(control_mode[4]), .I3(control_mode[7]), .O(n10_adj_4859));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam i4_4_lut_adj_1710.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(control_mode[6]), .I1(n10_adj_4859), .I2(control_mode[2]), 
            .I3(GND_net), .O(n20716));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i14199_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n18082), .I3(GND_net), .O(n22602));   // verilog/coms.v(127[12] 300[6])
    defparam i14199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1711 (.I0(n20608), .I1(control_mode[1]), .I2(GND_net), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(167[5:22])
    defparam i1_2_lut_adj_1711.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_3_lut (.I0(control_mode[0]), .I1(control_mode[1]), .I2(n20716), 
            .I3(GND_net), .O(n15_adj_4917));   // verilog/TinyFPGA_B.v(166[5:22])
    defparam i2_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i14200_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n18082), .I3(GND_net), .O(n22603));   // verilog/coms.v(127[12] 300[6])
    defparam i14200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14201_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n18082), .I3(GND_net), .O(n22604));   // verilog/coms.v(127[12] 300[6])
    defparam i14201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_65_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[23]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_4_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14202_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n18082), .I3(GND_net), .O(n22605));   // verilog/coms.v(127[12] 300[6])
    defparam i14202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14203_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n18082), .I3(GND_net), .O(n22606));   // verilog/coms.v(127[12] 300[6])
    defparam i14203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14204_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n18082), .I3(GND_net), .O(n22607));   // verilog/coms.v(127[12] 300[6])
    defparam i14204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14205_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n18082), .I3(GND_net), .O(n22608));   // verilog/coms.v(127[12] 300[6])
    defparam i14205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14206_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n18082), 
            .I3(GND_net), .O(n22609));   // verilog/coms.v(127[12] 300[6])
    defparam i14206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14207_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n18082), 
            .I3(GND_net), .O(n22610));   // verilog/coms.v(127[12] 300[6])
    defparam i14207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14208_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n18082), 
            .I3(GND_net), .O(n22611));   // verilog/coms.v(127[12] 300[6])
    defparam i14208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14209_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n18082), 
            .I3(GND_net), .O(n22612));   // verilog/coms.v(127[12] 300[6])
    defparam i14209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14210_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n18082), 
            .I3(GND_net), .O(n22613));   // verilog/coms.v(127[12] 300[6])
    defparam i14210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14211_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n18082), 
            .I3(GND_net), .O(n22614));   // verilog/coms.v(127[12] 300[6])
    defparam i14211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14212_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n18082), 
            .I3(GND_net), .O(n22615));   // verilog/coms.v(127[12] 300[6])
    defparam i14212_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14213_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n18082), 
            .I3(GND_net), .O(n22616));   // verilog/coms.v(127[12] 300[6])
    defparam i14213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14214_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n18082), 
            .I3(GND_net), .O(n22617));   // verilog/coms.v(127[12] 300[6])
    defparam i14214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14215_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n18082), 
            .I3(GND_net), .O(n22618));   // verilog/coms.v(127[12] 300[6])
    defparam i14215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14216_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n18082), 
            .I3(GND_net), .O(n22619));   // verilog/coms.v(127[12] 300[6])
    defparam i14216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14217_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n18082), 
            .I3(GND_net), .O(n22620));   // verilog/coms.v(127[12] 300[6])
    defparam i14217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14218_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n18082), 
            .I3(GND_net), .O(n22621));   // verilog/coms.v(127[12] 300[6])
    defparam i14218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14219_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n18082), 
            .I3(GND_net), .O(n22622));   // verilog/coms.v(127[12] 300[6])
    defparam i14219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14220_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n18082), 
            .I3(GND_net), .O(n22623));   // verilog/coms.v(127[12] 300[6])
    defparam i14220_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14221_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n18082), 
            .I3(GND_net), .O(n22624));   // verilog/coms.v(127[12] 300[6])
    defparam i14221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_583 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13905_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_4914), 
            .I3(n20781), .O(n22308));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13905_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14222_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n18082), 
            .I3(GND_net), .O(n22625));   // verilog/coms.v(127[12] 300[6])
    defparam i14222_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14223_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n18082), 
            .I3(GND_net), .O(n22626));   // verilog/coms.v(127[12] 300[6])
    defparam i14223_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14224_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n18082), 
            .I3(GND_net), .O(n22627));   // verilog/coms.v(127[12] 300[6])
    defparam i14224_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14225_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n18082), 
            .I3(GND_net), .O(n22628));   // verilog/coms.v(127[12] 300[6])
    defparam i14225_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14226_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n18082), 
            .I3(GND_net), .O(n22629));   // verilog/coms.v(127[12] 300[6])
    defparam i14226_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_3 (.CI(n31793), 
            .I0(GND_net), .I1(n25_adj_4999), .CO(n31794));
    SB_LUT4 i14227_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n18082), 
            .I3(GND_net), .O(n22630));   // verilog/coms.v(127[12] 300[6])
    defparam i14227_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14228_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n18082), 
            .I3(GND_net), .O(n22631));   // verilog/coms.v(127[12] 300[6])
    defparam i14228_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14229_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n18082), 
            .I3(GND_net), .O(n22632));   // verilog/coms.v(127[12] 300[6])
    defparam i14229_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14230_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n18082), .I3(GND_net), .O(n22633));   // verilog/coms.v(127[12] 300[6])
    defparam i14230_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14231_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n18082), .I3(GND_net), .O(n22634));   // verilog/coms.v(127[12] 300[6])
    defparam i14231_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14232_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n18082), .I3(GND_net), .O(n22635));   // verilog/coms.v(127[12] 300[6])
    defparam i14232_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14233_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n18082), .I3(GND_net), .O(n22636));   // verilog/coms.v(127[12] 300[6])
    defparam i14233_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14234_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n18082), .I3(GND_net), .O(n22637));   // verilog/coms.v(127[12] 300[6])
    defparam i14234_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14235_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n18082), .I3(GND_net), .O(n22638));   // verilog/coms.v(127[12] 300[6])
    defparam i14235_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14236_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n18082), .I3(GND_net), .O(n22639));   // verilog/coms.v(127[12] 300[6])
    defparam i14236_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14237_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n18082), .I3(GND_net), .O(n22640));   // verilog/coms.v(127[12] 300[6])
    defparam i14237_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14238_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n18082), .I3(GND_net), .O(n22641));   // verilog/coms.v(127[12] 300[6])
    defparam i14238_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14239_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n18082), .I3(GND_net), .O(n22642));   // verilog/coms.v(127[12] 300[6])
    defparam i14239_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14240_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n18082), .I3(GND_net), .O(n22643));   // verilog/coms.v(127[12] 300[6])
    defparam i14240_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14241_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n18082), .I3(GND_net), .O(n22644));   // verilog/coms.v(127[12] 300[6])
    defparam i14241_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14242_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n18082), .I3(GND_net), .O(n22645));   // verilog/coms.v(127[12] 300[6])
    defparam i14242_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(VCC_net), .CO(n31793));
    SB_LUT4 i14243_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n18082), .I3(GND_net), .O(n22646));   // verilog/coms.v(127[12] 300[6])
    defparam i14243_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14244_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n18082), .I3(GND_net), .O(n22647));   // verilog/coms.v(127[12] 300[6])
    defparam i14244_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14245_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n18082), .I3(GND_net), .O(n22648));   // verilog/coms.v(127[12] 300[6])
    defparam i14245_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14246_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n18082), .I3(GND_net), .O(n22649));   // verilog/coms.v(127[12] 300[6])
    defparam i14246_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14247_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n18082), .I3(GND_net), .O(n22650));   // verilog/coms.v(127[12] 300[6])
    defparam i14247_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14248_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n18082), .I3(GND_net), .O(n22651));   // verilog/coms.v(127[12] 300[6])
    defparam i14248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14249_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n18082), .I3(GND_net), .O(n22652));   // verilog/coms.v(127[12] 300[6])
    defparam i14249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14250_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n18082), .I3(GND_net), .O(n22653));   // verilog/coms.v(127[12] 300[6])
    defparam i14250_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14251_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n18082), .I3(GND_net), .O(n22654));   // verilog/coms.v(127[12] 300[6])
    defparam i14251_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14252_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n18082), .I3(GND_net), .O(n22655));   // verilog/coms.v(127[12] 300[6])
    defparam i14252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13906_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22309));   // verilog/coms.v(127[12] 300[6])
    defparam i13906_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13907_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n21865), 
            .I3(GND_net), .O(n22310));   // verilog/coms.v(127[12] 300[6])
    defparam i13907_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13908_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n21865), 
            .I3(GND_net), .O(n22311));   // verilog/coms.v(127[12] 300[6])
    defparam i13908_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13909_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n36883), .I3(GND_net), .O(n22312));   // verilog/coms.v(127[12] 300[6])
    defparam i13909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13911_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n21865), .I3(GND_net), .O(n22314));   // verilog/coms.v(127[12] 300[6])
    defparam i13911_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13912_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n21865), .I3(GND_net), .O(n22315));   // verilog/coms.v(127[12] 300[6])
    defparam i13912_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13913_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n38219), 
            .I3(GND_net), .O(n22316));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_3255_i1_3_lut (.I0(encoder0_position[0]), .I1(n25_adj_4880), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n532));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1712 (.I0(n15_adj_4901), .I1(data_ready), .I2(state_adj_5082[1]), 
            .I3(state_adj_5082[0]), .O(n35362));   // verilog/eeprom.v(25[8] 57[4])
    defparam i1_4_lut_adj_1712.LUT_INIT = 16'hccd0;
    SB_LUT4 i13915_4_lut (.I0(rw), .I1(state_adj_5082[0]), .I2(state_adj_5082[1]), 
            .I3(n3461), .O(n22318));   // verilog/eeprom.v(25[8] 57[4])
    defparam i13915_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i13916_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5088[1]), .I2(n13920), 
            .I3(n4_adj_4868), .O(n22319));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13916_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 i13917_3_lut (.I0(quadB_debounced_adj_4906), .I1(reg_B_adj_5099[0]), 
            .I2(n37217), .I3(GND_net), .O(n22320));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13917_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_644_4 (.CI(n30741), .I0(n40620), .I1(n23), .CO(n30742));
    SB_LUT4 i13918_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(state_7__N_3865[0]), 
            .I3(n15_adj_4901), .O(n22321));   // verilog/i2c_controller.v(89[8] 155[6])
    defparam i13918_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 encoder0_position_23__I_0_i1332_3_lut (.I0(n531), .I1(n1997), 
            .I2(n1948), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1332_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13919_3_lut (.I0(ID[0]), .I1(data[0]), .I2(data_ready), .I3(GND_net), 
            .O(n22322));   // verilog/TinyFPGA_B.v(233[10] 247[6])
    defparam i13919_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[0]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 i2_3_lut_adj_1713 (.I0(n62), .I1(n21971), .I2(delay_counter[31]), 
            .I3(GND_net), .O(n37894));
    defparam i2_3_lut_adj_1713.LUT_INIT = 16'h0808;
    SB_LUT4 encoder0_position_23__I_0_i1495_3_lut (.I0(n28040), .I1(n5701), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(encoder0_position_scaled_23__N_34[0]));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1495_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 i13923_4_lut (.I0(n36364), .I1(state[1]), .I2(state_3__N_369[1]), 
            .I3(n21969), .O(n22326));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13923_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i13927_4_lut (.I0(state_7__N_3881[3]), .I1(data[0]), .I2(n10_adj_5010), 
            .I3(n20726), .O(n22330));   // verilog/i2c_controller.v(89[8] 155[6])
    defparam i13927_4_lut.LUT_INIT = 16'hccca;
    SB_DFFESR delay_counter_1507__i20 (.Q(delay_counter[20]), .C(CLK_c), 
            .E(n21971), .D(n145), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_DFFESR delay_counter_1507__i19 (.Q(delay_counter[19]), .C(CLK_c), 
            .E(n21971), .D(n146), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 add_644_3_lut (.I0(duty[1]), .I1(n40620), .I2(n24), .I3(n30740), 
            .O(pwm_setpoint_22__N_11[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i13930_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n21865), .I3(GND_net), .O(n22333));   // verilog/coms.v(127[12] 300[6])
    defparam i13930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13931_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n21865), .I3(GND_net), .O(n22334));   // verilog/coms.v(127[12] 300[6])
    defparam i13931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13932_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n21865), .I3(GND_net), .O(n22335));   // verilog/coms.v(127[12] 300[6])
    defparam i13932_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_1507__i18 (.Q(delay_counter[18]), .C(CLK_c), 
            .E(n21971), .D(n147), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 i13933_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n21865), .I3(GND_net), .O(n22336));   // verilog/coms.v(127[12] 300[6])
    defparam i13933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13934_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n21865), .I3(GND_net), .O(n22337));   // verilog/coms.v(127[12] 300[6])
    defparam i13934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13935_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n21865), .I3(GND_net), .O(n22338));   // verilog/coms.v(127[12] 300[6])
    defparam i13935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_644_3 (.CI(n30740), .I0(n40620), .I1(n24), .CO(n30741));
    SB_DFF h1_42 (.Q(INLA_c), .C(clk32MHz), .D(hall1));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFFESR delay_counter_1507__i17 (.Q(delay_counter[17]), .C(CLK_c), 
            .E(n21971), .D(n148), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 unary_minus_4_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i13936_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n21865), .I3(GND_net), .O(n22339));   // verilog/coms.v(127[12] 300[6])
    defparam i13936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder1_position[23]), 
            .I2(n3_adj_4923), .I3(n31028), .O(displacement_23__N_58[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_1507__i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n21971), 
            .D(n165), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 encoder1_position_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder1_position[22]), 
            .I2(n3_adj_4923), .I3(n31027), .O(displacement_23__N_58[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_63_i1_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[0]), 
            .I3(encoder0_position_scaled[0]), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_63_i2_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[1]), 
            .I3(encoder0_position_scaled[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_63_i3_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[2]), 
            .I3(encoder0_position_scaled[2]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14253_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n18082), .I3(GND_net), .O(n22656));   // verilog/coms.v(127[12] 300[6])
    defparam i14253_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14254_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n18082), .I3(GND_net), .O(n22657));   // verilog/coms.v(127[12] 300[6])
    defparam i14254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_63_i4_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[3]), 
            .I3(encoder0_position_scaled[3]), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i4_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14255_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n18082), .I3(GND_net), .O(n22658));   // verilog/coms.v(127[12] 300[6])
    defparam i14255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14256_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n18082), .I3(GND_net), .O(n22659));   // verilog/coms.v(127[12] 300[6])
    defparam i14256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_63_i5_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[4]), 
            .I3(encoder0_position_scaled[4]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_DFFESR delay_counter_1507__i16 (.Q(delay_counter[16]), .C(CLK_c), 
            .E(n21971), .D(n149), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 add_644_2_lut (.I0(duty[0]), .I1(n40620), .I2(n25), .I3(VCC_net), 
            .O(pwm_setpoint_22__N_11[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i14257_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n18082), .I3(GND_net), .O(n22660));   // verilog/coms.v(127[12] 300[6])
    defparam i14257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_63_i6_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[5]), 
            .I3(encoder0_position_scaled[5]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14258_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n18082), .I3(GND_net), .O(n22661));   // verilog/coms.v(127[12] 300[6])
    defparam i14258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14259_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n18082), .I3(GND_net), .O(n22662));   // verilog/coms.v(127[12] 300[6])
    defparam i14259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14260_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n18082), .I3(GND_net), .O(n22663));   // verilog/coms.v(127[12] 300[6])
    defparam i14260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14261_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n18082), .I3(GND_net), .O(n22664));   // verilog/coms.v(127[12] 300[6])
    defparam i14261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14262_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n18082), .I3(GND_net), .O(n22665));   // verilog/coms.v(127[12] 300[6])
    defparam i14262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_63_i7_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[6]), 
            .I3(encoder0_position_scaled[6]), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i7_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14263_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n18082), .I3(GND_net), .O(n22666));   // verilog/coms.v(127[12] 300[6])
    defparam i14263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_63_i8_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[7]), 
            .I3(encoder0_position_scaled[7]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14264_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n18082), .I3(GND_net), .O(n22667));   // verilog/coms.v(127[12] 300[6])
    defparam i14264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14265_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n18082), .I3(GND_net), .O(n22668));   // verilog/coms.v(127[12] 300[6])
    defparam i14265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14266_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n18082), .I3(GND_net), .O(n22669));   // verilog/coms.v(127[12] 300[6])
    defparam i14266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14267_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n18082), .I3(GND_net), .O(n22670));   // verilog/coms.v(127[12] 300[6])
    defparam i14267_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_24 (.CI(n31027), .I0(encoder1_position[22]), 
            .I1(n3_adj_4923), .CO(n31028));
    SB_LUT4 i14268_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n18082), .I3(GND_net), .O(n22671));   // verilog/coms.v(127[12] 300[6])
    defparam i14268_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder1_position[21]), 
            .I2(n3_adj_4923), .I3(n31026), .O(displacement_23__N_58[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14269_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n18082), .I3(GND_net), .O(n22672));   // verilog/coms.v(127[12] 300[6])
    defparam i14269_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14270_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n18082), .I3(GND_net), .O(n22673));   // verilog/coms.v(127[12] 300[6])
    defparam i14270_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14271_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n18082), .I3(GND_net), .O(n22674));   // verilog/coms.v(127[12] 300[6])
    defparam i14271_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14272_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n18082), .I3(GND_net), .O(n22675));   // verilog/coms.v(127[12] 300[6])
    defparam i14272_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_63_i9_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[8]), 
            .I3(encoder0_position_scaled[8]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY encoder1_position_23__I_0_add_2_23 (.CI(n31026), .I0(encoder1_position[21]), 
            .I1(n3_adj_4923), .CO(n31027));
    SB_CARRY add_644_2 (.CI(VCC_net), .I0(n40620), .I1(n25), .CO(n30740));
    SB_LUT4 encoder1_position_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder1_position[20]), 
            .I2(n5_adj_4924), .I3(n31025), .O(displacement_23__N_58[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i1_1_lut (.I0(encoder0_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4944));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_63_i10_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[9]), 
            .I3(encoder0_position_scaled[9]), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_CARRY encoder1_position_23__I_0_add_2_22 (.CI(n31025), .I0(encoder1_position[20]), 
            .I1(n5_adj_4924), .CO(n31026));
    SB_LUT4 encoder1_position_23__I_0_inv_0_i2_1_lut (.I0(encoder0_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4943));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i3_1_lut (.I0(encoder0_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4942));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i4_1_lut (.I0(encoder0_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4941));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_65_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[0]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_63_i11_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[10]), 
            .I3(encoder0_position_scaled[10]), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i5_1_lut (.I0(encoder0_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4940));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_63_i12_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[11]), 
            .I3(encoder0_position_scaled[11]), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_65_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[1]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder1_position_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder1_position[19]), 
            .I2(n6_adj_4925), .I3(n31024), .O(displacement_23__N_58[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_63_i13_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[12]), 
            .I3(encoder0_position_scaled[12]), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i6_1_lut (.I0(encoder0_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4939));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1331_3_lut (.I0(n1943), .I1(n1996), 
            .I2(n1948), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1331_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1330_3_lut (.I0(n1942), .I1(n1995), 
            .I2(n1948), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1330_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1329_3_lut (.I0(n1941), .I1(n1994), 
            .I2(n1948), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1329_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1328_3_lut (.I0(n1940), .I1(n1993), 
            .I2(n1948), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1328_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_65_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[2]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder1_position_23__I_0_add_2_21 (.CI(n31024), .I0(encoder1_position[19]), 
            .I1(n6_adj_4925), .CO(n31025));
    SB_LUT4 mux_63_i14_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[13]), 
            .I3(encoder0_position_scaled[13]), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i7_1_lut (.I0(encoder0_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4938));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_65_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[3]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_63_i15_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[14]), 
            .I3(encoder0_position_scaled[14]), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder1_position_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder1_position[18]), 
            .I2(n7_adj_4926), .I3(n31023), .O(displacement_23__N_58[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i8_1_lut (.I0(encoder0_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4937));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_63_i16_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[15]), 
            .I3(encoder0_position_scaled[15]), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_23__I_0_i1327_3_lut (.I0(n1939), .I1(n1992), 
            .I2(n1948), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1327_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_63_i17_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[16]), 
            .I3(encoder0_position_scaled[16]), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i17_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_23__I_0_i1326_3_lut (.I0(n1938), .I1(n1991), 
            .I2(n1948), .I3(GND_net), .O(n2016));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1326_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder1_position_23__I_0_add_2_20 (.CI(n31023), .I0(encoder1_position[18]), 
            .I1(n7_adj_4926), .CO(n31024));
    SB_LUT4 encoder1_position_23__I_0_inv_0_i9_1_lut (.I0(encoder0_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4936));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_63_i18_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[17]), 
            .I3(encoder0_position_scaled[17]), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i10_1_lut (.I0(encoder0_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4935));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_65_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[4]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14273_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n18082), .I3(GND_net), .O(n22676));   // verilog/coms.v(127[12] 300[6])
    defparam i14273_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_65_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[5]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14274_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n18082), .I3(GND_net), .O(n22677));   // verilog/coms.v(127[12] 300[6])
    defparam i14274_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14275_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n18082), .I3(GND_net), .O(n22678));   // verilog/coms.v(127[12] 300[6])
    defparam i14275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder1_position[17]), 
            .I2(n8_adj_4927), .I3(n31022), .O(displacement_23__N_58[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14276_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n18082), .I3(GND_net), .O(n22679));   // verilog/coms.v(127[12] 300[6])
    defparam i14276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14277_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n18082), .I3(GND_net), .O(n22680));   // verilog/coms.v(127[12] 300[6])
    defparam i14277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1325_3_lut (.I0(n1937), .I1(n1990), 
            .I2(n1948), .I3(GND_net), .O(n2015));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1325_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14278_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position_scaled[7]), 
            .I2(n18082), .I3(GND_net), .O(n22681));   // verilog/coms.v(127[12] 300[6])
    defparam i14278_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_19 (.CI(n31022), .I0(encoder1_position[17]), 
            .I1(n8_adj_4927), .CO(n31023));
    SB_LUT4 encoder0_position_23__I_0_i1324_3_lut (.I0(n1936), .I1(n1989), 
            .I2(n1948), .I3(GND_net), .O(n2014));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1324_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1323_3_lut (.I0(n1935), .I1(n1988), 
            .I2(n1948), .I3(GND_net), .O(n2013));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1323_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder1_position[16]), 
            .I2(n9_adj_4928), .I3(n31021), .O(displacement_23__N_58[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_i1322_3_lut (.I0(n1934), .I1(n1987), 
            .I2(n1948), .I3(GND_net), .O(n2012));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1322_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14279_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position_scaled[6]), 
            .I2(n18082), .I3(GND_net), .O(n22682));   // verilog/coms.v(127[12] 300[6])
    defparam i14279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1321_3_lut (.I0(n1933), .I1(n1986), 
            .I2(n1948), .I3(GND_net), .O(n2011));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_65_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[6]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 unary_minus_4_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4856));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14280_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position_scaled[5]), 
            .I2(n18082), .I3(GND_net), .O(n22683));   // verilog/coms.v(127[12] 300[6])
    defparam i14280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14281_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position_scaled[4]), 
            .I2(n18082), .I3(GND_net), .O(n22684));   // verilog/coms.v(127[12] 300[6])
    defparam i14281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14282_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position_scaled[3]), 
            .I2(n18082), .I3(GND_net), .O(n22685));   // verilog/coms.v(127[12] 300[6])
    defparam i14282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_63_i19_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[18]), 
            .I3(encoder0_position_scaled[18]), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_65_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[7]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14283_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position_scaled[2]), 
            .I2(n18082), .I3(GND_net), .O(n22686));   // verilog/coms.v(127[12] 300[6])
    defparam i14283_3_lut.LUT_INIT = 16'hcaca;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_23__I_0_i1320_3_lut (.I0(n1932), .I1(n1985), 
            .I2(n1948), .I3(GND_net), .O(n2010));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14284_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position_scaled[1]), 
            .I2(n18082), .I3(GND_net), .O(n22687));   // verilog/coms.v(127[12] 300[6])
    defparam i14284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30262_1_lut (.I0(n700), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40291));
    defparam i30262_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i11_1_lut (.I0(encoder0_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4934));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_65_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[8]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14285_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position_scaled[0]), 
            .I2(n18082), .I3(GND_net), .O(n22688));   // verilog/coms.v(127[12] 300[6])
    defparam i14285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14286_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position_scaled[15]), 
            .I2(n18082), .I3(GND_net), .O(n22689));   // verilog/coms.v(127[12] 300[6])
    defparam i14286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30324_1_lut (.I0(n778), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40353));
    defparam i30324_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14287_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position_scaled[14]), 
            .I2(n18082), .I3(GND_net), .O(n22690));   // verilog/coms.v(127[12] 300[6])
    defparam i14287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1319_3_lut (.I0(n1931), .I1(n1984), 
            .I2(n1948), .I3(GND_net), .O(n2009));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1318_3_lut (.I0(n1930), .I1(n1983), 
            .I2(n1948), .I3(GND_net), .O(n2008));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder1_position_23__I_0_inv_0_i12_1_lut (.I0(encoder0_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4933));   // verilog/TinyFPGA_B.v(202[21:65])
    defparam encoder1_position_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14288_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position_scaled[13]), 
            .I2(n18082), .I3(GND_net), .O(n22691));   // verilog/coms.v(127[12] 300[6])
    defparam i14288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1317_3_lut (.I0(n1929), .I1(n1982), 
            .I2(n1948), .I3(GND_net), .O(n2007));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14289_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position_scaled[12]), 
            .I2(n18082), .I3(GND_net), .O(n22692));   // verilog/coms.v(127[12] 300[6])
    defparam i14289_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14290_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position_scaled[11]), 
            .I2(n18082), .I3(GND_net), .O(n22693));   // verilog/coms.v(127[12] 300[6])
    defparam i14290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_65_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15_adj_4917), .I3(n15), .O(motor_state_23__N_82[9]));   // verilog/TinyFPGA_B.v(166[5] 168[10])
    defparam mux_65_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14291_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position_scaled[10]), 
            .I2(n18082), .I3(GND_net), .O(n22694));   // verilog/coms.v(127[12] 300[6])
    defparam i14291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14292_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position_scaled[9]), 
            .I2(n18082), .I3(GND_net), .O(n22695));   // verilog/coms.v(127[12] 300[6])
    defparam i14292_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14293_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position_scaled[8]), 
            .I2(n18082), .I3(GND_net), .O(n22696));   // verilog/coms.v(127[12] 300[6])
    defparam i14293_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_18 (.CI(n31021), .I0(encoder1_position[16]), 
            .I1(n9_adj_4928), .CO(n31022));
    SB_LUT4 mux_63_i20_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[19]), 
            .I3(encoder0_position_scaled[19]), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_63_i21_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[20]), 
            .I3(encoder0_position_scaled[20]), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder1_position_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder1_position[15]), 
            .I2(n10_adj_4929), .I3(n31020), .O(displacement_23__N_58[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_17 (.CI(n31020), .I0(encoder1_position[15]), 
            .I1(n10_adj_4929), .CO(n31021));
    SB_LUT4 encoder1_position_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder1_position[14]), 
            .I2(n11_adj_4930), .I3(n31019), .O(displacement_23__N_58[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_16 (.CI(n31019), .I0(encoder1_position[14]), 
            .I1(n11_adj_4930), .CO(n31020));
    SB_LUT4 i14294_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position_scaled[22]), 
            .I2(n18082), .I3(GND_net), .O(n22697));   // verilog/coms.v(127[12] 300[6])
    defparam i14294_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_63_i22_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[21]), 
            .I3(encoder0_position_scaled[22]), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_63_i23_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[22]), 
            .I3(encoder0_position_scaled[22]), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14295_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position_scaled[22]), 
            .I2(n18082), .I3(GND_net), .O(n22698));   // verilog/coms.v(127[12] 300[6])
    defparam i14295_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14296_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position_scaled[22]), 
            .I2(n18082), .I3(GND_net), .O(n22699));   // verilog/coms.v(127[12] 300[6])
    defparam i14296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14297_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position_scaled[20]), 
            .I2(n18082), .I3(GND_net), .O(n22700));   // verilog/coms.v(127[12] 300[6])
    defparam i14297_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_63_i24_3_lut_4_lut (.I0(n20608), .I1(control_mode[1]), .I2(motor_state_23__N_82[23]), 
            .I3(encoder0_position_scaled[22]), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam mux_63_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i14298_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position_scaled[19]), 
            .I2(n18082), .I3(GND_net), .O(n22701));   // verilog/coms.v(127[12] 300[6])
    defparam i14298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder1_position[13]), 
            .I2(n12_adj_4931), .I3(n31018), .O(displacement_23__N_58[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14299_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position_scaled[18]), 
            .I2(n18082), .I3(GND_net), .O(n22702));   // verilog/coms.v(127[12] 300[6])
    defparam i14299_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_15 (.CI(n31018), .I0(encoder1_position[13]), 
            .I1(n12_adj_4931), .CO(n31019));
    SB_LUT4 i14300_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position_scaled[17]), 
            .I2(n18082), .I3(GND_net), .O(n22703));   // verilog/coms.v(127[12] 300[6])
    defparam i14300_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder1_position[12]), 
            .I2(n13_adj_4932), .I3(n31017), .O(displacement_23__N_58[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14301_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position_scaled[16]), 
            .I2(n18082), .I3(GND_net), .O(n22704));   // verilog/coms.v(127[12] 300[6])
    defparam i14301_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14302_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n18082), .I3(GND_net), .O(n22705));   // verilog/coms.v(127[12] 300[6])
    defparam i14302_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14303_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n18082), .I3(GND_net), .O(n22706));   // verilog/coms.v(127[12] 300[6])
    defparam i14303_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14304_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n18082), .I3(GND_net), .O(n22707));   // verilog/coms.v(127[12] 300[6])
    defparam i14304_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_26_lut (.I0(GND_net), .I1(n2000), 
            .I2(VCC_net), .I3(n31395), .O(n2053)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1361_25_lut (.I0(GND_net), .I1(n2001), 
            .I2(VCC_net), .I3(n31394), .O(n2054)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14305_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n18082), .I3(GND_net), .O(n22708));   // verilog/coms.v(127[12] 300[6])
    defparam i14305_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1361_25 (.CI(n31394), .I0(n2001), 
            .I1(VCC_net), .CO(n31395));
    SB_LUT4 encoder0_position_23__I_0_add_1361_24_lut (.I0(GND_net), .I1(n2002), 
            .I2(VCC_net), .I3(n31393), .O(n2055)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14306_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n18082), .I3(GND_net), .O(n22709));   // verilog/coms.v(127[12] 300[6])
    defparam i14306_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1361_24 (.CI(n31393), .I0(n2002), 
            .I1(VCC_net), .CO(n31394));
    SB_LUT4 i14307_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n18082), .I3(GND_net), .O(n22710));   // verilog/coms.v(127[12] 300[6])
    defparam i14307_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14308_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n18082), .I3(GND_net), .O(n22711));   // verilog/coms.v(127[12] 300[6])
    defparam i14308_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14309_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n18082), .I3(GND_net), .O(n22712));   // verilog/coms.v(127[12] 300[6])
    defparam i14309_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_14 (.CI(n31017), .I0(encoder1_position[12]), 
            .I1(n13_adj_4932), .CO(n31018));
    SB_LUT4 i14310_3_lut (.I0(\data_out_frame[4] [7]), .I1(ID[7]), .I2(n18082), 
            .I3(GND_net), .O(n22713));   // verilog/coms.v(127[12] 300[6])
    defparam i14310_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14311_3_lut (.I0(\data_out_frame[4] [6]), .I1(ID[6]), .I2(n18082), 
            .I3(GND_net), .O(n22714));   // verilog/coms.v(127[12] 300[6])
    defparam i14311_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14312_3_lut (.I0(\data_out_frame[4] [5]), .I1(ID[5]), .I2(n18082), 
            .I3(GND_net), .O(n22715));   // verilog/coms.v(127[12] 300[6])
    defparam i14312_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_23_lut (.I0(GND_net), .I1(n2003), 
            .I2(VCC_net), .I3(n31392), .O(n2056)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14313_3_lut (.I0(\data_out_frame[4] [4]), .I1(ID[4]), .I2(n18082), 
            .I3(GND_net), .O(n22716));   // verilog/coms.v(127[12] 300[6])
    defparam i14313_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14314_3_lut (.I0(\data_out_frame[4] [3]), .I1(ID[3]), .I2(n18082), 
            .I3(GND_net), .O(n22717));   // verilog/coms.v(127[12] 300[6])
    defparam i14314_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14315_3_lut (.I0(\data_out_frame[4] [2]), .I1(ID[2]), .I2(n18082), 
            .I3(GND_net), .O(n22718));   // verilog/coms.v(127[12] 300[6])
    defparam i14315_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1361_23 (.CI(n31392), .I0(n2003), 
            .I1(VCC_net), .CO(n31393));
    SB_LUT4 i14316_3_lut (.I0(\data_out_frame[4] [1]), .I1(ID[1]), .I2(n18082), 
            .I3(GND_net), .O(n22719));   // verilog/coms.v(127[12] 300[6])
    defparam i14316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_22_lut (.I0(GND_net), .I1(n2004), 
            .I2(VCC_net), .I3(n31391), .O(n2057)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_22 (.CI(n31391), .I0(n2004), 
            .I1(VCC_net), .CO(n31392));
    SB_LUT4 encoder0_position_23__I_0_add_1361_21_lut (.I0(GND_net), .I1(n2005), 
            .I2(VCC_net), .I3(n31390), .O(n2058)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_21 (.CI(n31390), .I0(n2005), 
            .I1(VCC_net), .CO(n31391));
    SB_LUT4 encoder0_position_23__I_0_add_1361_20_lut (.I0(GND_net), .I1(n2006), 
            .I2(VCC_net), .I3(n31389), .O(n2059)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_20 (.CI(n31389), .I0(n2006), 
            .I1(VCC_net), .CO(n31390));
    SB_LUT4 i14317_3_lut (.I0(\data_out_frame[4] [0]), .I1(ID[0]), .I2(n18082), 
            .I3(GND_net), .O(n22720));   // verilog/coms.v(127[12] 300[6])
    defparam i14317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14318_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n21865), 
            .I3(GND_net), .O(n22721));   // verilog/coms.v(127[12] 300[6])
    defparam i14318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_19_lut (.I0(GND_net), .I1(n2007), 
            .I2(VCC_net), .I3(n31388), .O(n2060)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_19 (.CI(n31388), .I0(n2007), 
            .I1(VCC_net), .CO(n31389));
    SB_LUT4 encoder1_position_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder1_position[11]), 
            .I2(n14_adj_4933), .I3(n31016), .O(displacement_23__N_58[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_23__I_0_add_1361_18_lut (.I0(GND_net), .I1(n2008), 
            .I2(VCC_net), .I3(n31387), .O(n2061)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14321_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n21865), 
            .I3(GND_net), .O(n22724));   // verilog/coms.v(127[12] 300[6])
    defparam i14321_3_lut.LUT_INIT = 16'hcaca;
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder1_position_23__I_0_add_2_13 (.CI(n31016), .I0(encoder1_position[11]), 
            .I1(n14_adj_4933), .CO(n31017));
    SB_LUT4 i14322_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n21865), 
            .I3(GND_net), .O(n22725));   // verilog/coms.v(127[12] 300[6])
    defparam i14322_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1361_18 (.CI(n31387), .I0(n2008), 
            .I1(VCC_net), .CO(n31388));
    SB_LUT4 encoder0_position_23__I_0_add_1361_17_lut (.I0(GND_net), .I1(n2009), 
            .I2(VCC_net), .I3(n31386), .O(n2062)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_17 (.CI(n31386), .I0(n2009), 
            .I1(VCC_net), .CO(n31387));
    SB_LUT4 encoder1_position_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder1_position[10]), 
            .I2(n15_adj_4934), .I3(n31015), .O(displacement_23__N_58[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1361_16_lut (.I0(GND_net), .I1(n2010), 
            .I2(VCC_net), .I3(n31385), .O(n2063)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_16 (.CI(n31385), .I0(n2010), 
            .I1(VCC_net), .CO(n31386));
    SB_LUT4 encoder0_position_23__I_0_add_1361_15_lut (.I0(GND_net), .I1(n2011), 
            .I2(VCC_net), .I3(n31384), .O(n2064)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_4_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4855));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_add_1361_15 (.CI(n31384), .I0(n2011), 
            .I1(VCC_net), .CO(n31385));
    SB_LUT4 i14323_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n21865), 
            .I3(GND_net), .O(n22726));   // verilog/coms.v(127[12] 300[6])
    defparam i14323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14324_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n21865), 
            .I3(GND_net), .O(n22727));   // verilog/coms.v(127[12] 300[6])
    defparam i14324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_14_lut (.I0(GND_net), .I1(n2012), 
            .I2(VCC_net), .I3(n31383), .O(n2065)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_14 (.CI(n31383), .I0(n2012), 
            .I1(VCC_net), .CO(n31384));
    SB_LUT4 encoder0_position_23__I_0_add_1361_13_lut (.I0(GND_net), .I1(n2013), 
            .I2(VCC_net), .I3(n31382), .O(n2066)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_13 (.CI(n31382), .I0(n2013), 
            .I1(VCC_net), .CO(n31383));
    SB_LUT4 encoder0_position_23__I_0_add_1361_12_lut (.I0(GND_net), .I1(n2014), 
            .I2(VCC_net), .I3(n31381), .O(n2067)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_12 (.CI(n31381), .I0(n2014), 
            .I1(VCC_net), .CO(n31382));
    SB_LUT4 encoder0_position_23__I_0_add_1361_11_lut (.I0(GND_net), .I1(n2015), 
            .I2(VCC_net), .I3(n31380), .O(n2068)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_11 (.CI(n31380), .I0(n2015), 
            .I1(VCC_net), .CO(n31381));
    SB_LUT4 i14325_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n21865), 
            .I3(GND_net), .O(n22728));   // verilog/coms.v(127[12] 300[6])
    defparam i14325_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_12 (.CI(n31015), .I0(encoder1_position[10]), 
            .I1(n15_adj_4934), .CO(n31016));
    SB_LUT4 encoder1_position_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder1_position[9]), 
            .I2(n16_adj_4935), .I3(n31014), .O(displacement_23__N_58[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_11 (.CI(n31014), .I0(encoder1_position[9]), 
            .I1(n16_adj_4935), .CO(n31015));
    SB_LUT4 encoder1_position_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder1_position[8]), 
            .I2(n17_adj_4936), .I3(n31013), .O(displacement_23__N_58[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_10 (.CI(n31013), .I0(encoder1_position[8]), 
            .I1(n17_adj_4936), .CO(n31014));
    SB_LUT4 encoder0_position_23__I_0_add_1361_10_lut (.I0(GND_net), .I1(n2016), 
            .I2(VCC_net), .I3(n31379), .O(n2069)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14326_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n21865), 
            .I3(GND_net), .O(n22729));   // verilog/coms.v(127[12] 300[6])
    defparam i14326_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1361_10 (.CI(n31379), .I0(n2016), 
            .I1(VCC_net), .CO(n31380));
    SB_LUT4 encoder0_position_23__I_0_add_1361_9_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n31378), .O(n2070)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder1_position_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder1_position[7]), 
            .I2(n18_adj_4937), .I3(n31012), .O(displacement_23__N_58[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_9 (.CI(n31012), .I0(encoder1_position[7]), 
            .I1(n18_adj_4937), .CO(n31013));
    SB_LUT4 encoder1_position_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder1_position[6]), 
            .I2(n19_adj_4938), .I3(n31011), .O(displacement_23__N_58[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_9 (.CI(n31378), .I0(n2017), 
            .I1(VCC_net), .CO(n31379));
    SB_LUT4 i14327_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n21865), 
            .I3(GND_net), .O(n22730));   // verilog/coms.v(127[12] 300[6])
    defparam i14327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_8_lut (.I0(GND_net), .I1(n2018), 
            .I2(GND_net), .I3(n31377), .O(n2071)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_8 (.CI(n31377), .I0(n2018), 
            .I1(GND_net), .CO(n31378));
    SB_LUT4 i14328_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n21865), 
            .I3(GND_net), .O(n22731));   // verilog/coms.v(127[12] 300[6])
    defparam i14328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1361_7_lut (.I0(n2073), .I1(n2019), 
            .I2(GND_net), .I3(n31376), .O(n39214)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i14329_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n21865), 
            .I3(GND_net), .O(n22732));   // verilog/coms.v(127[12] 300[6])
    defparam i14329_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1361_7 (.CI(n31376), .I0(n2019), 
            .I1(GND_net), .CO(n31377));
    SB_LUT4 encoder0_position_23__I_0_add_1361_6_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n31375), .O(n2073)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14330_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n21865), 
            .I3(GND_net), .O(n22733));   // verilog/coms.v(127[12] 300[6])
    defparam i14330_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1361_6 (.CI(n31375), .I0(n2020), 
            .I1(VCC_net), .CO(n31376));
    SB_LUT4 encoder0_position_23__I_0_add_1361_5_lut (.I0(n6_adj_4949), .I1(n2021), 
            .I2(GND_net), .I3(n31374), .O(n39272)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_5_lut.LUT_INIT = 16'hebbe;
    SB_CARRY encoder1_position_23__I_0_add_2_8 (.CI(n31011), .I0(encoder1_position[6]), 
            .I1(n19_adj_4938), .CO(n31012));
    SB_LUT4 encoder1_position_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder1_position[5]), 
            .I2(n20_adj_4939), .I3(n31010), .O(displacement_23__N_58[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_7 (.CI(n31010), .I0(encoder1_position[5]), 
            .I1(n20_adj_4939), .CO(n31011));
    SB_LUT4 encoder1_position_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder1_position[4]), 
            .I2(n21_adj_4940), .I3(n31009), .O(displacement_23__N_58[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder1_position_23__I_0_add_2_6 (.CI(n31009), .I0(encoder1_position[4]), 
            .I1(n21_adj_4940), .CO(n31010));
    SB_LUT4 encoder1_position_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder1_position[3]), 
            .I2(n22_adj_4941), .I3(n31008), .O(displacement_23__N_58[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1361_5 (.CI(n31374), .I0(n2021), 
            .I1(GND_net), .CO(n31375));
    SB_CARRY encoder1_position_23__I_0_add_2_5 (.CI(n31008), .I0(encoder1_position[3]), 
            .I1(n22_adj_4941), .CO(n31009));
    SB_LUT4 i14331_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n21865), 
            .I3(GND_net), .O(n22734));   // verilog/coms.v(127[12] 300[6])
    defparam i14331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14332_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n21865), 
            .I3(GND_net), .O(n22735));   // verilog/coms.v(127[12] 300[6])
    defparam i14332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder1_position_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder1_position[2]), 
            .I2(n23_adj_4942), .I3(n31007), .O(displacement_23__N_58[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14333_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n21865), 
            .I3(GND_net), .O(n22736));   // verilog/coms.v(127[12] 300[6])
    defparam i14333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14334_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n21865), 
            .I3(GND_net), .O(n22737));   // verilog/coms.v(127[12] 300[6])
    defparam i14334_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_4 (.CI(n31007), .I0(encoder1_position[2]), 
            .I1(n23_adj_4942), .CO(n31008));
    SB_LUT4 encoder1_position_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder1_position[1]), 
            .I2(n24_adj_4943), .I3(n31006), .O(displacement_23__N_58[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_1507_add_4_33_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[31]), .I3(n31552), .O(n134)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_1507_add_4_32_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[30]), .I3(n31551), .O(n135)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14335_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n21865), 
            .I3(GND_net), .O(n22738));   // verilog/coms.v(127[12] 300[6])
    defparam i14335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14336_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n21865), 
            .I3(GND_net), .O(n22739));   // verilog/coms.v(127[12] 300[6])
    defparam i14336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14337_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n21865), 
            .I3(GND_net), .O(n22740));   // verilog/coms.v(127[12] 300[6])
    defparam i14337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14338_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n21865), 
            .I3(GND_net), .O(n22741));   // verilog/coms.v(127[12] 300[6])
    defparam i14338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14339_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n21865), 
            .I3(GND_net), .O(n22742));   // verilog/coms.v(127[12] 300[6])
    defparam i14339_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder1_position_23__I_0_add_2_3 (.CI(n31006), .I0(encoder1_position[1]), 
            .I1(n24_adj_4943), .CO(n31007));
    SB_LUT4 encoder1_position_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder1_position[0]), 
            .I2(n25_adj_4944), .I3(VCC_net), .O(displacement_23__N_58[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder1_position_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1361_4_lut (.I0(n2076), .I1(n2022), 
            .I2(VCC_net), .I3(n31373), .O(n6_adj_4949)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder1_position_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder1_position[0]), 
            .I1(n25_adj_4944), .CO(n31006));
    SB_LUT4 i14340_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n21865), 
            .I3(GND_net), .O(n22743));   // verilog/coms.v(127[12] 300[6])
    defparam i14340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14341_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n21865), 
            .I3(GND_net), .O(n22744));   // verilog/coms.v(127[12] 300[6])
    defparam i14341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14342_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n21865), 
            .I3(GND_net), .O(n22745));   // verilog/coms.v(127[12] 300[6])
    defparam i14342_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1361_4 (.CI(n31373), .I0(n2022), 
            .I1(VCC_net), .CO(n31374));
    SB_LUT4 encoder0_position_23__I_0_add_1361_3_lut (.I0(GND_net), .I1(n532), 
            .I2(GND_net), .I3(n31372), .O(n2076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1361_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14343_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n21865), 
            .I3(GND_net), .O(n22746));   // verilog/coms.v(127[12] 300[6])
    defparam i14343_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1361_3 (.CI(n31372), .I0(n532), 
            .I1(GND_net), .CO(n31373));
    SB_CARRY encoder0_position_23__I_0_add_1361_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(VCC_net), .CO(n31372));
    SB_LUT4 add_1839_23_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n31371), .O(n5680)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1839_22_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n31370), .O(n5681)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14344_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n21865), 
            .I3(GND_net), .O(n22747));   // verilog/coms.v(127[12] 300[6])
    defparam i14344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14345_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n21865), 
            .I3(GND_net), .O(n22748));   // verilog/coms.v(127[12] 300[6])
    defparam i14345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14346_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n21865), 
            .I3(GND_net), .O(n22749));   // verilog/coms.v(127[12] 300[6])
    defparam i14346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14347_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n21865), 
            .I3(GND_net), .O(n22750));   // verilog/coms.v(127[12] 300[6])
    defparam i14347_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY delay_counter_1507_add_4_32 (.CI(n31551), .I0(GND_net), .I1(delay_counter[30]), 
            .CO(n31552));
    SB_LUT4 delay_counter_1507_add_4_31_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[29]), .I3(n31550), .O(n136)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1507_add_4_31 (.CI(n31550), .I0(GND_net), .I1(delay_counter[29]), 
            .CO(n31551));
    SB_CARRY add_1839_22 (.CI(n31370), .I0(GND_net), .I1(VCC_net), .CO(n31371));
    SB_LUT4 add_1839_21_lut (.I0(encoder0_position[23]), .I1(GND_net), .I2(n619), 
            .I3(n31369), .O(encoder0_position_scaled_23__N_34[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_1839_21 (.CI(n31369), .I0(GND_net), .I1(n619), .CO(n31370));
    SB_LUT4 delay_counter_1507_add_4_30_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[28]), .I3(n31549), .O(n137)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1507_add_4_30 (.CI(n31549), .I0(GND_net), .I1(delay_counter[28]), 
            .CO(n31550));
    SB_LUT4 add_1839_20_lut (.I0(GND_net), .I1(GND_net), .I2(n700), .I3(n31368), 
            .O(n5683)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1839_20 (.CI(n31368), .I0(GND_net), .I1(n700), .CO(n31369));
    SB_LUT4 i14348_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n21865), 
            .I3(GND_net), .O(n22751));   // verilog/coms.v(127[12] 300[6])
    defparam i14348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14349_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n21865), 
            .I3(GND_net), .O(n22752));   // verilog/coms.v(127[12] 300[6])
    defparam i14349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 delay_counter_1507_add_4_29_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[27]), .I3(n31548), .O(n138)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1839_19_lut (.I0(GND_net), .I1(GND_net), .I2(n778), .I3(n31367), 
            .O(n5684)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1839_19 (.CI(n31367), .I0(GND_net), .I1(n778), .CO(n31368));
    SB_LUT4 add_1839_18_lut (.I0(GND_net), .I1(GND_net), .I2(n856), .I3(n31366), 
            .O(n5685)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1507_add_4_29 (.CI(n31548), .I0(GND_net), .I1(delay_counter[27]), 
            .CO(n31549));
    SB_LUT4 i14350_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22753));   // verilog/coms.v(127[12] 300[6])
    defparam i14350_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1839_18 (.CI(n31366), .I0(GND_net), .I1(n856), .CO(n31367));
    SB_LUT4 delay_counter_1507_add_4_28_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[26]), .I3(n31547), .O(n139)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1839_17_lut (.I0(GND_net), .I1(GND_net), .I2(n934), .I3(n31365), 
            .O(n5686)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1839_17 (.CI(n31365), .I0(GND_net), .I1(n934), .CO(n31366));
    SB_CARRY delay_counter_1507_add_4_28 (.CI(n31547), .I0(GND_net), .I1(delay_counter[26]), 
            .CO(n31548));
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_10));   // verilog/TinyFPGA_B.v(143[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14008_3_lut (.I0(\data_in_frame[15] [7]), .I1(rx_data[7]), 
            .I2(n35561), .I3(GND_net), .O(n22411));   // verilog/coms.v(127[12] 300[6])
    defparam i14008_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14351_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22754));   // verilog/coms.v(127[12] 300[6])
    defparam i14351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14352_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22755));   // verilog/coms.v(127[12] 300[6])
    defparam i14352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14353_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22756));   // verilog/coms.v(127[12] 300[6])
    defparam i14353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14354_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22757));   // verilog/coms.v(127[12] 300[6])
    defparam i14354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 delay_counter_1507_add_4_27_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[25]), .I3(n31546), .O(n140)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1839_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1012), .I3(n31364), 
            .O(n5687)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1839_16 (.CI(n31364), .I0(GND_net), .I1(n1012), .CO(n31365));
    SB_LUT4 add_1839_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1090), .I3(n31363), 
            .O(n5688)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1839_15 (.CI(n31363), .I0(GND_net), .I1(n1090), .CO(n31364));
    SB_LUT4 add_1839_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1168), .I3(n31362), 
            .O(n5689)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14355_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22758));   // verilog/coms.v(127[12] 300[6])
    defparam i14355_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1839_14 (.CI(n31362), .I0(GND_net), .I1(n1168), .CO(n31363));
    SB_LUT4 i14356_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22759));   // verilog/coms.v(127[12] 300[6])
    defparam i14356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14357_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22760));   // verilog/coms.v(127[12] 300[6])
    defparam i14357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14358_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22761));   // verilog/coms.v(127[12] 300[6])
    defparam i14358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14359_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22762));   // verilog/coms.v(127[12] 300[6])
    defparam i14359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1316_3_lut (.I0(n1928), .I1(n1981), 
            .I2(n1948), .I3(GND_net), .O(n2006));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1316_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30363_1_lut (.I0(n1012), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40392));
    defparam i30363_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_i1315_3_lut (.I0(n1927), .I1(n1980), 
            .I2(n1948), .I3(GND_net), .O(n2005));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_i1314_3_lut (.I0(n1926), .I1(n1979), 
            .I2(n1948), .I3(GND_net), .O(n2004));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1314_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14360_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22763));   // verilog/coms.v(127[12] 300[6])
    defparam i14360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_i1313_3_lut (.I0(n1925), .I1(n1978), 
            .I2(n1948), .I3(GND_net), .O(n2003));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1313_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14361_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22764));   // verilog/coms.v(127[12] 300[6])
    defparam i14361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14362_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22765));   // verilog/coms.v(127[12] 300[6])
    defparam i14362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14363_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22766));   // verilog/coms.v(127[12] 300[6])
    defparam i14363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1839_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1246), .I3(n31361), 
            .O(n5690)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14364_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22767));   // verilog/coms.v(127[12] 300[6])
    defparam i14364_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1839_13 (.CI(n31361), .I0(GND_net), .I1(n1246), .CO(n31362));
    SB_LUT4 i14365_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22768));   // verilog/coms.v(127[12] 300[6])
    defparam i14365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14366_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22769));   // verilog/coms.v(127[12] 300[6])
    defparam i14366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14367_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22770));   // verilog/coms.v(127[12] 300[6])
    defparam i14367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14368_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22771));   // verilog/coms.v(127[12] 300[6])
    defparam i14368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14369_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22772));   // verilog/coms.v(127[12] 300[6])
    defparam i14369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14370_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22773));   // verilog/coms.v(127[12] 300[6])
    defparam i14370_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_58[23]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_58[22]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_58[21]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_58[20]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_58[19]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_58[18]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_58[17]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_58[16]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_58[15]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_58[14]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_58[13]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_58[12]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_58[11]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_58[10]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_58[9]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_58[8]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_58[7]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_58[6]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_58[5]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_58[4]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_58[3]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_58[2]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_58[1]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4995));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_1839_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1324), .I3(n31360), 
            .O(n5691)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14371_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22774));   // verilog/coms.v(127[12] 300[6])
    defparam i14371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14372_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22775));   // verilog/coms.v(127[12] 300[6])
    defparam i14372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14373_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22776));   // verilog/coms.v(127[12] 300[6])
    defparam i14373_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_1839_12 (.CI(n31360), .I0(GND_net), .I1(n1324), .CO(n31361));
    SB_LUT4 i14374_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22777));   // verilog/coms.v(127[12] 300[6])
    defparam i14374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1839_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1402), .I3(n31359), 
            .O(n5692)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1839_11 (.CI(n31359), .I0(GND_net), .I1(n1402), .CO(n31360));
    SB_LUT4 add_1839_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1480), .I3(n31358), 
            .O(n5693)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14375_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22778));   // verilog/coms.v(127[12] 300[6])
    defparam i14375_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14376_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22779));   // verilog/coms.v(127[12] 300[6])
    defparam i14376_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14377_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22780));   // verilog/coms.v(127[12] 300[6])
    defparam i14377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14378_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22781));   // verilog/coms.v(127[12] 300[6])
    defparam i14378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14379_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22782));   // verilog/coms.v(127[12] 300[6])
    defparam i14379_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14380_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n22783));   // verilog/coms.v(127[12] 300[6])
    defparam i14380_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY delay_counter_1507_add_4_27 (.CI(n31546), .I0(GND_net), .I1(delay_counter[25]), 
            .CO(n31547));
    SB_LUT4 delay_counter_1507_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[24]), .I3(n31545), .O(n141)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1839_10 (.CI(n31358), .I0(GND_net), .I1(n1480), .CO(n31359));
    SB_LUT4 i14381_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n37680), .I3(GND_net), .O(n22784));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14381_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY delay_counter_1507_add_4_26 (.CI(n31545), .I0(GND_net), .I1(delay_counter[24]), 
            .CO(n31546));
    SB_LUT4 i14382_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n37680), .I3(GND_net), .O(n22785));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1839_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1558), .I3(n31357), 
            .O(n5694)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1839_9 (.CI(n31357), .I0(GND_net), .I1(n1558), .CO(n31358));
    SB_LUT4 i14383_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n37680), .I3(GND_net), .O(n22786));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1839_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1636), .I3(n31356), 
            .O(n5695)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
            .C(clk32MHz), .D(n5680), .R(n2_adj_4976));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_LUT4 i6_4_lut_adj_1714 (.I0(delay_counter[0]), .I1(delay_counter[6]), 
            .I2(delay_counter[9]), .I3(delay_counter[3]), .O(n16_adj_5021));
    defparam i6_4_lut_adj_1714.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1715 (.I0(delay_counter[4]), .I1(delay_counter[8]), 
            .I2(delay_counter[7]), .I3(delay_counter[1]), .O(n17_adj_5020));
    defparam i7_4_lut_adj_1715.LUT_INIT = 16'hfffe;
    SB_LUT4 delay_counter_1507_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[23]), .I3(n31544), .O(n142)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1839_8 (.CI(n31356), .I0(GND_net), .I1(n1636), .CO(n31357));
    SB_LUT4 add_1839_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1714), .I3(n31355), 
            .O(n5696)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1507_add_4_25 (.CI(n31544), .I0(GND_net), .I1(delay_counter[23]), 
            .CO(n31545));
    SB_CARRY add_1839_7 (.CI(n31355), .I0(GND_net), .I1(n1714), .CO(n31356));
    SB_LUT4 add_1839_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1792), .I3(n31354), 
            .O(n5697)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1839_6 (.CI(n31354), .I0(GND_net), .I1(n1792), .CO(n31355));
    SB_LUT4 i14384_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n37680), .I3(GND_net), .O(n22787));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 delay_counter_1507_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[22]), .I3(n31543), .O(n143)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1839_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1870), .I3(n31353), 
            .O(n5698)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1839_5 (.CI(n31353), .I0(GND_net), .I1(n1870), .CO(n31354));
    SB_CARRY delay_counter_1507_add_4_24 (.CI(n31543), .I0(GND_net), .I1(delay_counter[22]), 
            .CO(n31544));
    SB_LUT4 add_1839_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1948), .I3(n31352), 
            .O(n5699)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1839_4 (.CI(n31352), .I0(GND_net), .I1(n1948), .CO(n31353));
    SB_LUT4 add_1839_3_lut (.I0(GND_net), .I1(GND_net), .I2(n2026), .I3(n31351), 
            .O(n5700)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1839_3 (.CI(n31351), .I0(GND_net), .I1(n2026), .CO(n31352));
    SB_LUT4 i14385_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n37680), .I3(GND_net), .O(n22788));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 delay_counter_1507_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[21]), .I3(n31542), .O(n144)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9_4_lut_adj_1716 (.I0(n17_adj_5020), .I1(delay_counter[5]), 
            .I2(n16_adj_5021), .I3(delay_counter[2]), .O(n37568));
    defparam i9_4_lut_adj_1716.LUT_INIT = 16'hfffe;
    SB_LUT4 i14386_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n37680), .I3(GND_net), .O(n22789));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1839_2_lut (.I0(GND_net), .I1(GND_net), .I2(n28040), .I3(VCC_net), 
            .O(n5701)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1839_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14387_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n37680), .I3(GND_net), .O(n22790));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14387_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY delay_counter_1507_add_4_23 (.CI(n31542), .I0(GND_net), .I1(delay_counter[21]), 
            .CO(n31543));
    SB_CARRY add_1839_2 (.CI(VCC_net), .I0(GND_net), .I1(n28040), .CO(n31351));
    SB_LUT4 i2_4_lut_adj_1717 (.I0(n37568), .I1(delay_counter[12]), .I2(delay_counter[10]), 
            .I3(delay_counter[11]), .O(n37536));
    defparam i2_4_lut_adj_1717.LUT_INIT = 16'hffec;
    SB_LUT4 encoder0_position_23__I_0_add_1308_24_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n31350), .O(n1975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_3_lut (.I0(delay_counter[14]), .I1(delay_counter[15]), .I2(delay_counter[17]), 
            .I3(GND_net), .O(n8_adj_5016));
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_1718 (.I0(delay_counter[16]), .I1(n8_adj_5016), 
            .I2(n37536), .I3(delay_counter[13]), .O(n37529));
    defparam i4_4_lut_adj_1718.LUT_INIT = 16'hfeee;
    SB_LUT4 encoder0_position_23__I_0_add_1308_23_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n31349), .O(n1976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14388_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n37680), .I3(GND_net), .O(n22791));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 delay_counter_1507_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[20]), .I3(n31541), .O(n145)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_23 (.CI(n31349), .I0(n1923), 
            .I1(VCC_net), .CO(n31350));
    SB_LUT4 encoder0_position_23__I_0_add_1308_22_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n31348), .O(n1977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_1719 (.I0(delay_counter[22]), .I1(n37529), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5017));
    defparam i2_4_lut_adj_1719.LUT_INIT = 16'ha8a0;
    SB_LUT4 i2_2_lut_adj_1720 (.I0(delay_counter[28]), .I1(delay_counter[29]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4948));
    defparam i2_2_lut_adj_1720.LUT_INIT = 16'heeee;
    SB_CARRY encoder0_position_23__I_0_add_1308_22 (.CI(n31348), .I0(n1924), 
            .I1(VCC_net), .CO(n31349));
    SB_CARRY delay_counter_1507_add_4_22 (.CI(n31541), .I0(GND_net), .I1(delay_counter[20]), 
            .CO(n31542));
    SB_LUT4 i14389_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n37680), .I3(GND_net), .O(n22792));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14389_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1308_21_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n31347), .O(n1978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_1507_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[19]), .I3(n31540), .O(n146)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14390_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n37680), .I3(GND_net), .O(n22793));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14390_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i6_4_lut_adj_1721 (.I0(delay_counter[24]), .I1(delay_counter[30]), 
            .I2(delay_counter[26]), .I3(delay_counter[27]), .O(n14_adj_4947));
    defparam i6_4_lut_adj_1721.LUT_INIT = 16'hfffe;
    SB_LUT4 i14391_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n37680), .I3(GND_net), .O(n22794));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14391_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1308_21 (.CI(n31347), .I0(n1925), 
            .I1(VCC_net), .CO(n31348));
    SB_LUT4 encoder0_position_23__I_0_add_1308_20_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n31346), .O(n1979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut_adj_1722 (.I0(n7_adj_5017), .I1(delay_counter[20]), 
            .I2(delay_counter[21]), .I3(delay_counter[23]), .O(n37535));
    defparam i4_4_lut_adj_1722.LUT_INIT = 16'h8000;
    SB_LUT4 i14392_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n37680), .I3(GND_net), .O(n22795));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14392_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14393_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n37680), .I3(GND_net), .O(n22796));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14393_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1308_20 (.CI(n31346), .I0(n1926), 
            .I1(VCC_net), .CO(n31347));
    SB_LUT4 i14394_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n37680), .I3(GND_net), .O(n22797));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14394_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14395_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n37680), .I3(GND_net), .O(n22798));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14395_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14396_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n37680), .I3(GND_net), .O(n22799));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14396_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1308_19_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n31345), .O(n1980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14397_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n37680), .I3(GND_net), .O(n22800));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14397_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1308_19 (.CI(n31345), .I0(n1927), 
            .I1(VCC_net), .CO(n31346));
    SB_CARRY delay_counter_1507_add_4_21 (.CI(n31540), .I0(GND_net), .I1(delay_counter[19]), 
            .CO(n31541));
    SB_LUT4 encoder0_position_23__I_0_add_1308_18_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n31344), .O(n1981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_18 (.CI(n31344), .I0(n1928), 
            .I1(VCC_net), .CO(n31345));
    SB_LUT4 delay_counter_1507_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[18]), .I3(n31539), .O(n147)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1308_17_lut (.I0(GND_net), .I1(n1929), 
            .I2(VCC_net), .I3(n31343), .O(n1982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_17 (.CI(n31343), .I0(n1929), 
            .I1(VCC_net), .CO(n31344));
    SB_LUT4 encoder0_position_23__I_0_add_1308_16_lut (.I0(GND_net), .I1(n1930), 
            .I2(VCC_net), .I3(n31342), .O(n1983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_16 (.CI(n31342), .I0(n1930), 
            .I1(VCC_net), .CO(n31343));
    SB_LUT4 encoder0_position_23__I_0_add_1308_15_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n31341), .O(n1984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1507_add_4_20 (.CI(n31539), .I0(GND_net), .I1(delay_counter[18]), 
            .CO(n31540));
    SB_LUT4 delay_counter_1507_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[17]), .I3(n31538), .O(n148)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_15 (.CI(n31341), .I0(n1931), 
            .I1(VCC_net), .CO(n31342));
    SB_LUT4 encoder0_position_23__I_0_add_1308_14_lut (.I0(GND_net), .I1(n1932), 
            .I2(VCC_net), .I3(n31340), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1507_add_4_19 (.CI(n31538), .I0(GND_net), .I1(delay_counter[17]), 
            .CO(n31539));
    SB_CARRY encoder0_position_23__I_0_add_1308_14 (.CI(n31340), .I0(n1932), 
            .I1(VCC_net), .CO(n31341));
    SB_LUT4 encoder0_position_23__I_0_add_1308_13_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n31339), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14398_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n37680), .I3(GND_net), .O(n22801));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14398_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1308_13 (.CI(n31339), .I0(n1933), 
            .I1(VCC_net), .CO(n31340));
    SB_LUT4 encoder0_position_23__I_0_add_1308_12_lut (.I0(GND_net), .I1(n1934), 
            .I2(VCC_net), .I3(n31338), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_12 (.CI(n31338), .I0(n1934), 
            .I1(VCC_net), .CO(n31339));
    SB_LUT4 encoder0_position_23__I_0_add_1308_11_lut (.I0(GND_net), .I1(n1935), 
            .I2(VCC_net), .I3(n31337), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14399_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n37680), .I3(GND_net), .O(n22802));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14399_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1308_11 (.CI(n31337), .I0(n1935), 
            .I1(VCC_net), .CO(n31338));
    SB_LUT4 encoder0_position_23__I_0_add_1308_10_lut (.I0(GND_net), .I1(n1936), 
            .I2(VCC_net), .I3(n31336), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_10 (.CI(n31336), .I0(n1936), 
            .I1(VCC_net), .CO(n31337));
    SB_LUT4 encoder0_position_23__I_0_add_1308_9_lut (.I0(GND_net), .I1(n1937), 
            .I2(VCC_net), .I3(n31335), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_9 (.CI(n31335), .I0(n1937), 
            .I1(VCC_net), .CO(n31336));
    SB_LUT4 encoder0_position_23__I_0_add_1308_8_lut (.I0(GND_net), .I1(n1938), 
            .I2(VCC_net), .I3(n31334), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_8 (.CI(n31334), .I0(n1938), 
            .I1(VCC_net), .CO(n31335));
    SB_LUT4 encoder0_position_23__I_0_add_1308_7_lut (.I0(GND_net), .I1(n1939), 
            .I2(GND_net), .I3(n31333), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_7 (.CI(n31333), .I0(n1939), 
            .I1(GND_net), .CO(n31334));
    SB_LUT4 encoder0_position_23__I_0_add_1308_6_lut (.I0(GND_net), .I1(n1940), 
            .I2(GND_net), .I3(n31332), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_6 (.CI(n31332), .I0(n1940), 
            .I1(GND_net), .CO(n31333));
    SB_LUT4 encoder0_position_23__I_0_add_1308_5_lut (.I0(GND_net), .I1(n1941), 
            .I2(VCC_net), .I3(n31331), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_5 (.CI(n31331), .I0(n1941), 
            .I1(VCC_net), .CO(n31332));
    SB_LUT4 encoder0_position_23__I_0_add_1308_4_lut (.I0(GND_net), .I1(n1942), 
            .I2(GND_net), .I3(n31330), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_4 (.CI(n31330), .I0(n1942), 
            .I1(GND_net), .CO(n31331));
    SB_LUT4 delay_counter_1507_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[16]), .I3(n31537), .O(n149)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1308_3_lut (.I0(GND_net), .I1(n1943), 
            .I2(VCC_net), .I3(n31329), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1308_3 (.CI(n31329), .I0(n1943), 
            .I1(VCC_net), .CO(n31330));
    SB_LUT4 i14400_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n37680), .I3(GND_net), .O(n22803));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14400_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1308_2_lut (.I0(GND_net), .I1(n531), 
            .I2(GND_net), .I3(VCC_net), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1308_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
            .C(clk32MHz), .D(n5681), .R(n2_adj_4976));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_LUT4 i14401_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n37680), .I3(GND_net), .O(n22804));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14401_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1308_2 (.CI(VCC_net), .I0(n531), 
            .I1(GND_net), .CO(n31329));
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[19]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[18]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_LUT4 i14402_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n37680), .I3(GND_net), .O(n22805));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14402_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14403_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n37680), .I3(GND_net), .O(n22806));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14403_3_lut.LUT_INIT = 16'hacac;
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[17]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_LUT4 encoder0_position_23__I_0_add_1255_23_lut (.I0(GND_net), .I1(n1844), 
            .I2(VCC_net), .I3(n31328), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_23_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[16]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[15]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[14]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[13]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[12]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[11]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(clk32MHz), .D(encoder0_position_scaled_23__N_34[10]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[9]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[8]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[7]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[6]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[5]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[4]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[3]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[2]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[1]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[22]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[21]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[20]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[19]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[18]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[17]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[16]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[15]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[14]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[13]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[12]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[11]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[10]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[9]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[8]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[7]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[6]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[5]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[4]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[3]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[2]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk32MHz), .D(pwm_setpoint_22__N_11[1]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 i14404_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n37680), .I3(GND_net), .O(n22807));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14404_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_1507__i15 (.Q(delay_counter[15]), .C(CLK_c), 
            .E(n21971), .D(n150), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_CARRY delay_counter_1507_add_4_18 (.CI(n31537), .I0(GND_net), .I1(delay_counter[16]), 
            .CO(n31538));
    SB_LUT4 encoder0_position_23__I_0_add_1255_22_lut (.I0(GND_net), .I1(n1845), 
            .I2(VCC_net), .I3(n31327), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_22 (.CI(n31327), .I0(n1845), 
            .I1(VCC_net), .CO(n31328));
    SB_LUT4 encoder0_position_23__I_0_add_1255_21_lut (.I0(GND_net), .I1(n1846), 
            .I2(VCC_net), .I3(n31326), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_21 (.CI(n31326), .I0(n1846), 
            .I1(VCC_net), .CO(n31327));
    SB_LUT4 encoder0_position_23__I_0_add_1255_20_lut (.I0(GND_net), .I1(n1847), 
            .I2(VCC_net), .I3(n31325), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_20 (.CI(n31325), .I0(n1847), 
            .I1(VCC_net), .CO(n31326));
    SB_LUT4 encoder0_position_23__I_0_add_1255_19_lut (.I0(GND_net), .I1(n1848), 
            .I2(VCC_net), .I3(n31324), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_19 (.CI(n31324), .I0(n1848), 
            .I1(VCC_net), .CO(n31325));
    SB_LUT4 encoder0_position_23__I_0_add_1255_18_lut (.I0(GND_net), .I1(n1849), 
            .I2(VCC_net), .I3(n31323), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_18 (.CI(n31323), .I0(n1849), 
            .I1(VCC_net), .CO(n31324));
    SB_LUT4 i14020_3_lut (.I0(\data_in_frame[14] [3]), .I1(rx_data[3]), 
            .I2(n35562), .I3(GND_net), .O(n22423));   // verilog/coms.v(127[12] 300[6])
    defparam i14020_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1255_17_lut (.I0(GND_net), .I1(n1850), 
            .I2(VCC_net), .I3(n31322), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_17 (.CI(n31322), .I0(n1850), 
            .I1(VCC_net), .CO(n31323));
    SB_LUT4 encoder0_position_23__I_0_add_1255_16_lut (.I0(GND_net), .I1(n1851), 
            .I2(VCC_net), .I3(n31321), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_16 (.CI(n31321), .I0(n1851), 
            .I1(VCC_net), .CO(n31322));
    SB_LUT4 encoder0_position_23__I_0_add_1255_15_lut (.I0(GND_net), .I1(n1852), 
            .I2(VCC_net), .I3(n31320), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_15 (.CI(n31320), .I0(n1852), 
            .I1(VCC_net), .CO(n31321));
    SB_LUT4 delay_counter_1507_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[15]), .I3(n31536), .O(n150)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1255_14_lut (.I0(GND_net), .I1(n1853), 
            .I2(VCC_net), .I3(n31319), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_14 (.CI(n31319), .I0(n1853), 
            .I1(VCC_net), .CO(n31320));
    SB_LUT4 i14405_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n37680), .I3(GND_net), .O(n22808));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14405_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1255_13_lut (.I0(GND_net), .I1(n1854), 
            .I2(VCC_net), .I3(n31318), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1507_add_4_17 (.CI(n31536), .I0(GND_net), .I1(delay_counter[15]), 
            .CO(n31537));
    SB_CARRY encoder0_position_23__I_0_add_1255_13 (.CI(n31318), .I0(n1854), 
            .I1(VCC_net), .CO(n31319));
    SB_LUT4 i14406_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n37680), .I3(GND_net), .O(n22809));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14406_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1255_12_lut (.I0(GND_net), .I1(n1855), 
            .I2(VCC_net), .I3(n31317), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_12 (.CI(n31317), .I0(n1855), 
            .I1(VCC_net), .CO(n31318));
    SB_LUT4 i14407_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n37680), .I3(GND_net), .O(n22810));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14407_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14408_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n37680), .I3(GND_net), .O(n22811));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14408_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14409_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n37680), .I3(GND_net), .O(n22812));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14409_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1255_11_lut (.I0(GND_net), .I1(n1856), 
            .I2(VCC_net), .I3(n31316), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14410_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n37680), .I3(GND_net), .O(n22813));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14410_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1255_11 (.CI(n31316), .I0(n1856), 
            .I1(VCC_net), .CO(n31317));
    SB_LUT4 delay_counter_1507_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[14]), .I3(n31535), .O(n151)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1255_10_lut (.I0(GND_net), .I1(n1857), 
            .I2(VCC_net), .I3(n31315), .O(n1910)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_10 (.CI(n31315), .I0(n1857), 
            .I1(VCC_net), .CO(n31316));
    SB_LUT4 encoder0_position_23__I_0_add_1255_9_lut (.I0(GND_net), .I1(n1858), 
            .I2(VCC_net), .I3(n31314), .O(n1911)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_9 (.CI(n31314), .I0(n1858), 
            .I1(VCC_net), .CO(n31315));
    SB_CARRY delay_counter_1507_add_4_16 (.CI(n31535), .I0(GND_net), .I1(delay_counter[14]), 
            .CO(n31536));
    SB_LUT4 delay_counter_1507_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[13]), .I3(n31534), .O(n152)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1255_8_lut (.I0(GND_net), .I1(n1859), 
            .I2(VCC_net), .I3(n31313), .O(n1912)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_8 (.CI(n31313), .I0(n1859), 
            .I1(VCC_net), .CO(n31314));
    SB_LUT4 encoder0_position_23__I_0_add_1255_7_lut (.I0(GND_net), .I1(n1860), 
            .I2(GND_net), .I3(n31312), .O(n1913)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_7 (.CI(n31312), .I0(n1860), 
            .I1(GND_net), .CO(n31313));
    SB_CARRY delay_counter_1507_add_4_15 (.CI(n31534), .I0(GND_net), .I1(delay_counter[13]), 
            .CO(n31535));
    SB_LUT4 encoder0_position_23__I_0_add_1255_6_lut (.I0(GND_net), .I1(n1861), 
            .I2(GND_net), .I3(n31311), .O(n1914)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_1507_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[12]), .I3(n31533), .O(n153)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1507_add_4_14 (.CI(n31533), .I0(GND_net), .I1(delay_counter[12]), 
            .CO(n31534));
    SB_CARRY encoder0_position_23__I_0_add_1255_6 (.CI(n31311), .I0(n1861), 
            .I1(GND_net), .CO(n31312));
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_23__I_0_add_1255_5_lut (.I0(GND_net), .I1(n1862), 
            .I2(VCC_net), .I3(n31310), .O(n1915)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_5_lut.LUT_INIT = 16'hC33C;
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 delay_counter_1507_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[11]), .I3(n31532), .O(n154)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_5 (.CI(n31310), .I0(n1862), 
            .I1(VCC_net), .CO(n31311));
    SB_LUT4 encoder0_position_23__I_0_add_1255_4_lut (.I0(GND_net), .I1(n1863), 
            .I2(GND_net), .I3(n31309), .O(n1916)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_1507__i14 (.Q(delay_counter[14]), .C(CLK_c), 
            .E(n21971), .D(n151), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_CARRY encoder0_position_23__I_0_add_1255_4 (.CI(n31309), .I0(n1863), 
            .I1(GND_net), .CO(n31310));
    SB_LUT4 encoder0_position_23__I_0_add_1255_3_lut (.I0(GND_net), .I1(n1864), 
            .I2(VCC_net), .I3(n31308), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_3 (.CI(n31308), .I0(n1864), 
            .I1(VCC_net), .CO(n31309));
    SB_LUT4 encoder0_position_23__I_0_add_1255_2_lut (.I0(GND_net), .I1(n530), 
            .I2(GND_net), .I3(VCC_net), .O(n1918)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1255_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1255_2 (.CI(VCC_net), .I0(n530), 
            .I1(GND_net), .CO(n31308));
    SB_LUT4 i14411_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n37680), .I3(GND_net), .O(n22814));   // verilog/neopixel.v(35[12] 117[6])
    defparam i14411_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY delay_counter_1507_add_4_13 (.CI(n31532), .I0(GND_net), .I1(delay_counter[11]), 
            .CO(n31533));
    SB_LUT4 encoder0_position_23__I_0_add_1202_22_lut (.I0(GND_net), .I1(n1766), 
            .I2(VCC_net), .I3(n31307), .O(n1819)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1202_21_lut (.I0(GND_net), .I1(n1767), 
            .I2(VCC_net), .I3(n31306), .O(n1820)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_21 (.CI(n31306), .I0(n1767), 
            .I1(VCC_net), .CO(n31307));
    SB_LUT4 encoder0_position_23__I_0_add_1202_20_lut (.I0(GND_net), .I1(n1768), 
            .I2(VCC_net), .I3(n31305), .O(n1821)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_20 (.CI(n31305), .I0(n1768), 
            .I1(VCC_net), .CO(n31306));
    SB_LUT4 delay_counter_1507_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[10]), .I3(n31531), .O(n155)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1202_19_lut (.I0(GND_net), .I1(n1769), 
            .I2(VCC_net), .I3(n31304), .O(n1822)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_19 (.CI(n31304), .I0(n1769), 
            .I1(VCC_net), .CO(n31305));
    SB_CARRY delay_counter_1507_add_4_12 (.CI(n31531), .I0(GND_net), .I1(delay_counter[10]), 
            .CO(n31532));
    SB_LUT4 encoder0_position_23__I_0_add_1202_18_lut (.I0(GND_net), .I1(n1770), 
            .I2(VCC_net), .I3(n31303), .O(n1823)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_1507_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[9]), .I3(n31530), .O(n156)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1507_add_4_11 (.CI(n31530), .I0(GND_net), .I1(delay_counter[9]), 
            .CO(n31531));
    SB_CARRY encoder0_position_23__I_0_add_1202_18 (.CI(n31303), .I0(n1770), 
            .I1(VCC_net), .CO(n31304));
    SB_LUT4 encoder0_position_23__I_0_add_1202_17_lut (.I0(GND_net), .I1(n1771), 
            .I2(VCC_net), .I3(n31302), .O(n1824)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_17 (.CI(n31302), .I0(n1771), 
            .I1(VCC_net), .CO(n31303));
    SB_LUT4 i14009_3_lut (.I0(\data_in_frame[15] [6]), .I1(rx_data[6]), 
            .I2(n35561), .I3(GND_net), .O(n22412));   // verilog/coms.v(127[12] 300[6])
    defparam i14009_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14010_3_lut (.I0(\data_in_frame[15] [5]), .I1(rx_data[5]), 
            .I2(n35561), .I3(GND_net), .O(n22413));   // verilog/coms.v(127[12] 300[6])
    defparam i14010_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1202_16_lut (.I0(GND_net), .I1(n1772), 
            .I2(VCC_net), .I3(n31301), .O(n1825)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_16 (.CI(n31301), .I0(n1772), 
            .I1(VCC_net), .CO(n31302));
    SB_LUT4 encoder0_position_23__I_0_add_1202_15_lut (.I0(GND_net), .I1(n1773), 
            .I2(VCC_net), .I3(n31300), .O(n1826)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_1507_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[8]), .I3(n31529), .O(n157)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_15 (.CI(n31300), .I0(n1773), 
            .I1(VCC_net), .CO(n31301));
    SB_LUT4 encoder0_position_23__I_0_add_1202_14_lut (.I0(GND_net), .I1(n1774), 
            .I2(VCC_net), .I3(n31299), .O(n1827)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_14 (.CI(n31299), .I0(n1774), 
            .I1(VCC_net), .CO(n31300));
    SB_CARRY delay_counter_1507_add_4_10 (.CI(n31529), .I0(GND_net), .I1(delay_counter[8]), 
            .CO(n31530));
    SB_LUT4 encoder0_position_23__I_0_add_1202_13_lut (.I0(GND_net), .I1(n1775), 
            .I2(VCC_net), .I3(n31298), .O(n1828)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_1507_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[7]), .I3(n31528), .O(n158)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_13 (.CI(n31298), .I0(n1775), 
            .I1(VCC_net), .CO(n31299));
    SB_CARRY delay_counter_1507_add_4_9 (.CI(n31528), .I0(GND_net), .I1(delay_counter[7]), 
            .CO(n31529));
    SB_LUT4 encoder0_position_23__I_0_add_1202_12_lut (.I0(GND_net), .I1(n1776), 
            .I2(VCC_net), .I3(n31297), .O(n1829)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_12 (.CI(n31297), .I0(n1776), 
            .I1(VCC_net), .CO(n31298));
    SB_LUT4 delay_counter_1507_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[6]), .I3(n31527), .O(n159)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14415_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n21865), .I3(GND_net), .O(n22818));   // verilog/coms.v(127[12] 300[6])
    defparam i14415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4999));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4998));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_add_1202_11_lut (.I0(GND_net), .I1(n1777), 
            .I2(VCC_net), .I3(n31296), .O(n1830)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_11 (.CI(n31296), .I0(n1777), 
            .I1(VCC_net), .CO(n31297));
    SB_LUT4 encoder0_position_23__I_0_add_1202_10_lut (.I0(GND_net), .I1(n1778), 
            .I2(VCC_net), .I3(n31295), .O(n1831)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14416_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n21865), .I3(GND_net), .O(n22819));   // verilog/coms.v(127[12] 300[6])
    defparam i14416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14011_3_lut (.I0(\data_in_frame[15] [4]), .I1(rx_data[4]), 
            .I2(n35561), .I3(GND_net), .O(n22414));   // verilog/coms.v(127[12] 300[6])
    defparam i14011_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14012_3_lut (.I0(\data_in_frame[15] [3]), .I1(rx_data[3]), 
            .I2(n35561), .I3(GND_net), .O(n22415));   // verilog/coms.v(127[12] 300[6])
    defparam i14012_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1202_10 (.CI(n31295), .I0(n1778), 
            .I1(VCC_net), .CO(n31296));
    SB_LUT4 encoder0_position_23__I_0_add_1202_9_lut (.I0(GND_net), .I1(n1779), 
            .I2(VCC_net), .I3(n31294), .O(n1832)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14417_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n21865), .I3(GND_net), .O(n22820));   // verilog/coms.v(127[12] 300[6])
    defparam i14417_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1202_9 (.CI(n31294), .I0(n1779), 
            .I1(VCC_net), .CO(n31295));
    SB_CARRY delay_counter_1507_add_4_8 (.CI(n31527), .I0(GND_net), .I1(delay_counter[6]), 
            .CO(n31528));
    SB_LUT4 encoder0_position_23__I_0_add_1202_8_lut (.I0(GND_net), .I1(n1780), 
            .I2(VCC_net), .I3(n31293), .O(n1833)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_8 (.CI(n31293), .I0(n1780), 
            .I1(VCC_net), .CO(n31294));
    SB_LUT4 i14418_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n21865), .I3(GND_net), .O(n22821));   // verilog/coms.v(127[12] 300[6])
    defparam i14418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1202_7_lut (.I0(GND_net), .I1(n1781), 
            .I2(GND_net), .I3(n31292), .O(n1834)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_7 (.CI(n31292), .I0(n1781), 
            .I1(GND_net), .CO(n31293));
    SB_LUT4 encoder0_position_23__I_0_add_1202_6_lut (.I0(GND_net), .I1(n1782), 
            .I2(GND_net), .I3(n31291), .O(n1835)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_1507_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[5]), .I3(n31526), .O(n160)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_6 (.CI(n31291), .I0(n1782), 
            .I1(GND_net), .CO(n31292));
    SB_LUT4 encoder0_position_23__I_0_add_1202_5_lut (.I0(GND_net), .I1(n1783), 
            .I2(VCC_net), .I3(n31290), .O(n1836)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1507_add_4_7 (.CI(n31526), .I0(GND_net), .I1(delay_counter[5]), 
            .CO(n31527));
    SB_CARRY encoder0_position_23__I_0_add_1202_5 (.CI(n31290), .I0(n1783), 
            .I1(VCC_net), .CO(n31291));
    SB_LUT4 delay_counter_1507_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[4]), .I3(n31525), .O(n161)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1507_add_4_6 (.CI(n31525), .I0(GND_net), .I1(delay_counter[4]), 
            .CO(n31526));
    SB_LUT4 encoder0_position_23__I_0_add_1202_4_lut (.I0(GND_net), .I1(n1784), 
            .I2(GND_net), .I3(n31289), .O(n1837)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14013_3_lut (.I0(\data_in_frame[15] [2]), .I1(rx_data[2]), 
            .I2(n35561), .I3(GND_net), .O(n22416));   // verilog/coms.v(127[12] 300[6])
    defparam i14013_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4997));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14014_3_lut (.I0(\data_in_frame[15] [1]), .I1(rx_data[1]), 
            .I2(n35561), .I3(GND_net), .O(n22417));   // verilog/coms.v(127[12] 300[6])
    defparam i14014_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1202_4 (.CI(n31289), .I0(n1784), 
            .I1(GND_net), .CO(n31290));
    SB_LUT4 encoder0_position_23__I_0_add_1202_3_lut (.I0(GND_net), .I1(n1785), 
            .I2(VCC_net), .I3(n31288), .O(n1838)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14015_3_lut (.I0(\data_in_frame[15] [0]), .I1(rx_data[0]), 
            .I2(n35561), .I3(GND_net), .O(n22418));   // verilog/coms.v(127[12] 300[6])
    defparam i14015_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1202_3 (.CI(n31288), .I0(n1785), 
            .I1(VCC_net), .CO(n31289));
    SB_LUT4 encoder0_position_23__I_0_add_1202_2_lut (.I0(GND_net), .I1(n529), 
            .I2(GND_net), .I3(VCC_net), .O(n1839)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1202_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14016_3_lut (.I0(\data_in_frame[14] [7]), .I1(rx_data[7]), 
            .I2(n35562), .I3(GND_net), .O(n22419));   // verilog/coms.v(127[12] 300[6])
    defparam i14016_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 delay_counter_1507_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[3]), .I3(n31524), .O(n162)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1202_2 (.CI(VCC_net), .I0(n529), 
            .I1(GND_net), .CO(n31288));
    SB_CARRY delay_counter_1507_add_4_5 (.CI(n31524), .I0(GND_net), .I1(delay_counter[3]), 
            .CO(n31525));
    SB_LUT4 encoder0_position_23__I_0_add_1149_21_lut (.I0(GND_net), .I1(n1688), 
            .I2(VCC_net), .I3(n31287), .O(n1741)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_1507_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[2]), .I3(n31523), .O(n163)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1149_20_lut (.I0(GND_net), .I1(n1689), 
            .I2(VCC_net), .I3(n31286), .O(n1742)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY delay_counter_1507_add_4_4 (.CI(n31523), .I0(GND_net), .I1(delay_counter[2]), 
            .CO(n31524));
    SB_CARRY encoder0_position_23__I_0_add_1149_20 (.CI(n31286), .I0(n1689), 
            .I1(VCC_net), .CO(n31287));
    SB_LUT4 encoder0_position_23__I_0_add_1149_19_lut (.I0(GND_net), .I1(n1690), 
            .I2(VCC_net), .I3(n31285), .O(n1743)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_19 (.CI(n31285), .I0(n1690), 
            .I1(VCC_net), .CO(n31286));
    SB_LUT4 encoder0_position_23__I_0_add_1149_18_lut (.I0(GND_net), .I1(n1691), 
            .I2(VCC_net), .I3(n31284), .O(n1744)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_18 (.CI(n31284), .I0(n1691), 
            .I1(VCC_net), .CO(n31285));
    SB_LUT4 encoder0_position_23__I_0_add_1149_17_lut (.I0(GND_net), .I1(n1692), 
            .I2(VCC_net), .I3(n31283), .O(n1745)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 delay_counter_1507_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[1]), .I3(n31522), .O(n164)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_17 (.CI(n31283), .I0(n1692), 
            .I1(VCC_net), .CO(n31284));
    SB_LUT4 i14419_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n21865), .I3(GND_net), .O(n22822));   // verilog/coms.v(127[12] 300[6])
    defparam i14419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1149_16_lut (.I0(GND_net), .I1(n1693), 
            .I2(VCC_net), .I3(n31282), .O(n1746)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_16 (.CI(n31282), .I0(n1693), 
            .I1(VCC_net), .CO(n31283));
    SB_LUT4 i14420_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n21865), .I3(GND_net), .O(n22823));   // verilog/coms.v(127[12] 300[6])
    defparam i14420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1149_15_lut (.I0(GND_net), .I1(n1694), 
            .I2(VCC_net), .I3(n31281), .O(n1747)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_15 (.CI(n31281), .I0(n1694), 
            .I1(VCC_net), .CO(n31282));
    SB_CARRY delay_counter_1507_add_4_3 (.CI(n31522), .I0(GND_net), .I1(delay_counter[1]), 
            .CO(n31523));
    SB_LUT4 encoder0_position_23__I_0_add_1149_14_lut (.I0(GND_net), .I1(n1695), 
            .I2(VCC_net), .I3(n31280), .O(n1748)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14017_3_lut (.I0(\data_in_frame[14] [6]), .I1(rx_data[6]), 
            .I2(n35562), .I3(GND_net), .O(n22420));   // verilog/coms.v(127[12] 300[6])
    defparam i14017_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_23__I_0_add_1149_14 (.CI(n31280), .I0(n1695), 
            .I1(VCC_net), .CO(n31281));
    SB_LUT4 encoder0_position_23__I_0_add_1149_13_lut (.I0(GND_net), .I1(n1696), 
            .I2(VCC_net), .I3(n31279), .O(n1749)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_13 (.CI(n31279), .I0(n1696), 
            .I1(VCC_net), .CO(n31280));
    SB_LUT4 encoder0_position_23__I_0_add_1149_12_lut (.I0(GND_net), .I1(n1697), 
            .I2(VCC_net), .I3(n31278), .O(n1750)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14421_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n21865), .I3(GND_net), .O(n22824));   // verilog/coms.v(127[12] 300[6])
    defparam i14421_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1149_12 (.CI(n31278), .I0(n1697), 
            .I1(VCC_net), .CO(n31279));
    SB_LUT4 i14422_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n21865), .I3(GND_net), .O(n22825));   // verilog/coms.v(127[12] 300[6])
    defparam i14422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 delay_counter_1507_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(delay_counter[0]), .I3(VCC_net), .O(n165)) /* synthesis syn_instantiated=1 */ ;
    defparam delay_counter_1507_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1149_11_lut (.I0(GND_net), .I1(n1698), 
            .I2(VCC_net), .I3(n31277), .O(n1751)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_11 (.CI(n31277), .I0(n1698), 
            .I1(VCC_net), .CO(n31278));
    SB_CARRY delay_counter_1507_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(delay_counter[0]), 
            .CO(n31522));
    SB_LUT4 encoder0_position_23__I_0_add_1149_10_lut (.I0(GND_net), .I1(n1699), 
            .I2(VCC_net), .I3(n31276), .O(n1752)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_10 (.CI(n31276), .I0(n1699), 
            .I1(VCC_net), .CO(n31277));
    SB_LUT4 encoder0_position_23__I_0_add_1149_9_lut (.I0(GND_net), .I1(n1700), 
            .I2(VCC_net), .I3(n31275), .O(n1753)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_9 (.CI(n31275), .I0(n1700), 
            .I1(VCC_net), .CO(n31276));
    SB_LUT4 encoder0_position_23__I_0_add_1149_8_lut (.I0(GND_net), .I1(n1701), 
            .I2(VCC_net), .I3(n31274), .O(n1754)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_8 (.CI(n31274), .I0(n1701), 
            .I1(VCC_net), .CO(n31275));
    SB_LUT4 i14423_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n21865), .I3(GND_net), .O(n22826));   // verilog/coms.v(127[12] 300[6])
    defparam i14423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1149_7_lut (.I0(GND_net), .I1(n1702), 
            .I2(GND_net), .I3(n31273), .O(n1755)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_7 (.CI(n31273), .I0(n1702), 
            .I1(GND_net), .CO(n31274));
    SB_LUT4 i14424_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n21865), .I3(GND_net), .O(n22827));   // verilog/coms.v(127[12] 300[6])
    defparam i14424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1149_6_lut (.I0(GND_net), .I1(n1703), 
            .I2(GND_net), .I3(n31272), .O(n1756)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_6 (.CI(n31272), .I0(n1703), 
            .I1(GND_net), .CO(n31273));
    SB_LUT4 encoder0_position_23__I_0_add_1149_5_lut (.I0(GND_net), .I1(n1704), 
            .I2(VCC_net), .I3(n31271), .O(n1757)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_5 (.CI(n31271), .I0(n1704), 
            .I1(VCC_net), .CO(n31272));
    SB_LUT4 encoder0_position_23__I_0_add_1149_4_lut (.I0(GND_net), .I1(n1705), 
            .I2(GND_net), .I3(n31270), .O(n1758)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14425_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n21865), .I3(GND_net), .O(n22828));   // verilog/coms.v(127[12] 300[6])
    defparam i14425_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1149_4 (.CI(n31270), .I0(n1705), 
            .I1(GND_net), .CO(n31271));
    SB_LUT4 encoder0_position_23__I_0_add_1149_3_lut (.I0(GND_net), .I1(n1706), 
            .I2(VCC_net), .I3(n31269), .O(n1759)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14426_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n21865), .I3(GND_net), .O(n22829));   // verilog/coms.v(127[12] 300[6])
    defparam i14426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14427_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n21865), .I3(GND_net), .O(n22830));   // verilog/coms.v(127[12] 300[6])
    defparam i14427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14428_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n21865), .I3(GND_net), .O(n22831));   // verilog/coms.v(127[12] 300[6])
    defparam i14428_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1149_3 (.CI(n31269), .I0(n1706), 
            .I1(VCC_net), .CO(n31270));
    SB_LUT4 encoder0_position_23__I_0_add_1149_2_lut (.I0(GND_net), .I1(n528), 
            .I2(GND_net), .I3(VCC_net), .O(n1760)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1149_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1149_2 (.CI(VCC_net), .I0(n528), 
            .I1(GND_net), .CO(n31269));
    SB_LUT4 encoder0_position_23__I_0_add_1096_20_lut (.I0(GND_net), .I1(n1610), 
            .I2(VCC_net), .I3(n31268), .O(n1663)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1096_19_lut (.I0(GND_net), .I1(n1611), 
            .I2(VCC_net), .I3(n31267), .O(n1664)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_19 (.CI(n31267), .I0(n1611), 
            .I1(VCC_net), .CO(n31268));
    SB_LUT4 encoder0_position_23__I_0_add_1096_18_lut (.I0(GND_net), .I1(n1612), 
            .I2(VCC_net), .I3(n31266), .O(n1665)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_18 (.CI(n31266), .I0(n1612), 
            .I1(VCC_net), .CO(n31267));
    SB_LUT4 i14429_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n21865), .I3(GND_net), .O(n22832));   // verilog/coms.v(127[12] 300[6])
    defparam i14429_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1096_17_lut (.I0(GND_net), .I1(n1613), 
            .I2(VCC_net), .I3(n31265), .O(n1666)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_17 (.CI(n31265), .I0(n1613), 
            .I1(VCC_net), .CO(n31266));
    SB_LUT4 encoder0_position_23__I_0_add_1096_16_lut (.I0(GND_net), .I1(n1614), 
            .I2(VCC_net), .I3(n31264), .O(n1667)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_16 (.CI(n31264), .I0(n1614), 
            .I1(VCC_net), .CO(n31265));
    SB_LUT4 encoder0_position_23__I_0_add_1096_15_lut (.I0(GND_net), .I1(n1615), 
            .I2(VCC_net), .I3(n31263), .O(n1668)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_15 (.CI(n31263), .I0(n1615), 
            .I1(VCC_net), .CO(n31264));
    SB_LUT4 encoder0_position_23__I_0_add_1096_14_lut (.I0(GND_net), .I1(n1616), 
            .I2(VCC_net), .I3(n31262), .O(n1669)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_14 (.CI(n31262), .I0(n1616), 
            .I1(VCC_net), .CO(n31263));
    SB_LUT4 encoder0_position_23__I_0_add_1096_13_lut (.I0(GND_net), .I1(n1617), 
            .I2(VCC_net), .I3(n31261), .O(n1670)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_13 (.CI(n31261), .I0(n1617), 
            .I1(VCC_net), .CO(n31262));
    SB_LUT4 i14430_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n21865), .I3(GND_net), .O(n22833));   // verilog/coms.v(127[12] 300[6])
    defparam i14430_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1096_12_lut (.I0(GND_net), .I1(n1618), 
            .I2(VCC_net), .I3(n31260), .O(n1671)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14431_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n21865), .I3(GND_net), .O(n22834));   // verilog/coms.v(127[12] 300[6])
    defparam i14431_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1096_12 (.CI(n31260), .I0(n1618), 
            .I1(VCC_net), .CO(n31261));
    SB_LUT4 i14432_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n21865), .I3(GND_net), .O(n22835));   // verilog/coms.v(127[12] 300[6])
    defparam i14432_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14433_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n21865), .I3(GND_net), .O(n22836));   // verilog/coms.v(127[12] 300[6])
    defparam i14433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1096_11_lut (.I0(GND_net), .I1(n1619), 
            .I2(VCC_net), .I3(n31259), .O(n1672)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_11 (.CI(n31259), .I0(n1619), 
            .I1(VCC_net), .CO(n31260));
    SB_LUT4 encoder0_position_23__I_0_add_1096_10_lut (.I0(GND_net), .I1(n1620), 
            .I2(VCC_net), .I3(n31258), .O(n1673)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_10 (.CI(n31258), .I0(n1620), 
            .I1(VCC_net), .CO(n31259));
    SB_LUT4 i14434_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n21865), .I3(GND_net), .O(n22837));   // verilog/coms.v(127[12] 300[6])
    defparam i14434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1096_9_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n31257), .O(n1674)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_9 (.CI(n31257), .I0(n1621), 
            .I1(VCC_net), .CO(n31258));
    SB_LUT4 encoder0_position_23__I_0_add_1096_8_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n31256), .O(n1675)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_8 (.CI(n31256), .I0(n1622), 
            .I1(VCC_net), .CO(n31257));
    SB_LUT4 encoder0_position_23__I_0_add_1096_7_lut (.I0(GND_net), .I1(n1623), 
            .I2(GND_net), .I3(n31255), .O(n1676)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14435_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n21865), .I3(GND_net), .O(n22838));   // verilog/coms.v(127[12] 300[6])
    defparam i14435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14436_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n21865), .I3(GND_net), .O(n22839));   // verilog/coms.v(127[12] 300[6])
    defparam i14436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14437_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n21865), .I3(GND_net), .O(n22840));   // verilog/coms.v(127[12] 300[6])
    defparam i14437_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1096_7 (.CI(n31255), .I0(n1623), 
            .I1(GND_net), .CO(n31256));
    SB_LUT4 encoder0_position_23__I_0_add_1096_6_lut (.I0(GND_net), .I1(n1624), 
            .I2(GND_net), .I3(n31254), .O(n1677)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_6 (.CI(n31254), .I0(n1624), 
            .I1(GND_net), .CO(n31255));
    SB_LUT4 encoder0_position_23__I_0_add_1096_5_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n31253), .O(n1678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_5 (.CI(n31253), .I0(n1625), 
            .I1(VCC_net), .CO(n31254));
    SB_LUT4 add_644_24_lut (.I0(duty[22]), .I1(n40620), .I2(n3), .I3(n30761), 
            .O(pwm_setpoint_22__N_11[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i14444_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_4914), 
            .I3(n20776), .O(n22847));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14444_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14445_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n38219), 
            .I3(GND_net), .O(n22848));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i14445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i7_4_lut_adj_1723 (.I0(n37535), .I1(n14_adj_4947), .I2(n10_adj_4948), 
            .I3(delay_counter[25]), .O(n62));
    defparam i7_4_lut_adj_1723.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_add_1096_4_lut (.I0(GND_net), .I1(n1626), 
            .I2(GND_net), .I3(n31252), .O(n1679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_4 (.CI(n31252), .I0(n1626), 
            .I1(GND_net), .CO(n31253));
    SB_LUT4 i2_3_lut_adj_1724 (.I0(delay_counter[31]), .I1(n21971), .I2(n62), 
            .I3(GND_net), .O(n22157));   // verilog/TinyFPGA_B.v(237[10:34])
    defparam i2_3_lut_adj_1724.LUT_INIT = 16'h4040;
    SB_LUT4 encoder0_position_23__I_0_add_1096_3_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n31251), .O(n1680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_3 (.CI(n31251), .I0(n1627), 
            .I1(VCC_net), .CO(n31252));
    SB_LUT4 i2_2_lut_adj_1725 (.I0(ID[1]), .I1(ID[2]), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_4858));   // verilog/TinyFPGA_B.v(235[8:13])
    defparam i2_2_lut_adj_1725.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1726 (.I0(ID[7]), .I1(ID[4]), .I2(ID[5]), .I3(ID[6]), 
            .O(n14_adj_4857));   // verilog/TinyFPGA_B.v(235[8:13])
    defparam i6_4_lut_adj_1726.LUT_INIT = 16'hfffe;
    SB_LUT4 i30093_4_lut (.I0(ID[0]), .I1(n14_adj_4857), .I2(n10_adj_4858), 
            .I3(ID[3]), .O(n21971));   // verilog/TinyFPGA_B.v(235[8:13])
    defparam i30093_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i14446_3_lut (.I0(quadA_debounced_adj_4905), .I1(reg_B_adj_5099[1]), 
            .I2(n37217), .I3(GND_net), .O(n22849));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i14446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1096_2_lut (.I0(GND_net), .I1(n527), 
            .I2(GND_net), .I3(VCC_net), .O(n1681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1096_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1096_2 (.CI(VCC_net), .I0(n527), 
            .I1(GND_net), .CO(n31251));
    SB_LUT4 encoder0_position_23__I_0_add_1043_19_lut (.I0(GND_net), .I1(n1532), 
            .I2(VCC_net), .I3(n31250), .O(n1585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_1043_18_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n31249), .O(n1586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_18 (.CI(n31249), .I0(n1533), 
            .I1(VCC_net), .CO(n31250));
    SB_LUT4 i14447_3_lut (.I0(ID[1]), .I1(data[1]), .I2(data_ready), .I3(GND_net), 
            .O(n22850));   // verilog/TinyFPGA_B.v(233[10] 247[6])
    defparam i14447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1043_17_lut (.I0(GND_net), .I1(n1534), 
            .I2(VCC_net), .I3(n31248), .O(n1587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_17 (.CI(n31248), .I0(n1534), 
            .I1(VCC_net), .CO(n31249));
    SB_LUT4 i14448_3_lut (.I0(ID[2]), .I1(data[2]), .I2(data_ready), .I3(GND_net), 
            .O(n22851));   // verilog/TinyFPGA_B.v(233[10] 247[6])
    defparam i14448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1043_16_lut (.I0(GND_net), .I1(n1535), 
            .I2(VCC_net), .I3(n31247), .O(n1588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_16 (.CI(n31247), .I0(n1535), 
            .I1(VCC_net), .CO(n31248));
    SB_LUT4 i14449_3_lut (.I0(ID[3]), .I1(data[3]), .I2(data_ready), .I3(GND_net), 
            .O(n22852));   // verilog/TinyFPGA_B.v(233[10] 247[6])
    defparam i14449_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14450_3_lut (.I0(ID[4]), .I1(data[4]), .I2(data_ready), .I3(GND_net), 
            .O(n22853));   // verilog/TinyFPGA_B.v(233[10] 247[6])
    defparam i14450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14451_3_lut (.I0(ID[5]), .I1(data[5]), .I2(data_ready), .I3(GND_net), 
            .O(n22854));   // verilog/TinyFPGA_B.v(233[10] 247[6])
    defparam i14451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1043_15_lut (.I0(GND_net), .I1(n1536), 
            .I2(VCC_net), .I3(n31246), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_15 (.CI(n31246), .I0(n1536), 
            .I1(VCC_net), .CO(n31247));
    SB_LUT4 encoder0_position_23__I_0_add_1043_14_lut (.I0(GND_net), .I1(n1537), 
            .I2(VCC_net), .I3(n31245), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_14 (.CI(n31245), .I0(n1537), 
            .I1(VCC_net), .CO(n31246));
    SB_LUT4 encoder0_position_23__I_0_add_1043_13_lut (.I0(GND_net), .I1(n1538), 
            .I2(VCC_net), .I3(n31244), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_13 (.CI(n31244), .I0(n1538), 
            .I1(VCC_net), .CO(n31245));
    SB_LUT4 i14452_3_lut (.I0(ID[6]), .I1(data[6]), .I2(data_ready), .I3(GND_net), 
            .O(n22855));   // verilog/TinyFPGA_B.v(233[10] 247[6])
    defparam i14452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_1043_12_lut (.I0(GND_net), .I1(n1539), 
            .I2(VCC_net), .I3(n31243), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_12 (.CI(n31243), .I0(n1539), 
            .I1(VCC_net), .CO(n31244));
    SB_LUT4 encoder0_position_23__I_0_add_1043_11_lut (.I0(GND_net), .I1(n1540), 
            .I2(VCC_net), .I3(n31242), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_11 (.CI(n31242), .I0(n1540), 
            .I1(VCC_net), .CO(n31243));
    SB_LUT4 encoder0_position_23__I_0_add_1043_10_lut (.I0(GND_net), .I1(n1541), 
            .I2(VCC_net), .I3(n31241), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_10 (.CI(n31241), .I0(n1541), 
            .I1(VCC_net), .CO(n31242));
    SB_LUT4 encoder0_position_23__I_0_add_1043_9_lut (.I0(GND_net), .I1(n1542), 
            .I2(VCC_net), .I3(n31240), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_9 (.CI(n31240), .I0(n1542), 
            .I1(VCC_net), .CO(n31241));
    SB_LUT4 encoder0_position_23__I_0_add_1043_8_lut (.I0(GND_net), .I1(n1543), 
            .I2(VCC_net), .I3(n31239), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14453_3_lut (.I0(ID[7]), .I1(data[7]), .I2(data_ready), .I3(GND_net), 
            .O(n22856));   // verilog/TinyFPGA_B.v(233[10] 247[6])
    defparam i14453_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_1043_8 (.CI(n31239), .I0(n1543), 
            .I1(VCC_net), .CO(n31240));
    SB_LUT4 encoder0_position_23__I_0_add_1043_7_lut (.I0(GND_net), .I1(n1544), 
            .I2(GND_net), .I3(n31238), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_7 (.CI(n31238), .I0(n1544), 
            .I1(GND_net), .CO(n31239));
    SB_LUT4 encoder0_position_23__I_0_add_1043_6_lut (.I0(GND_net), .I1(n1545), 
            .I2(GND_net), .I3(n31237), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_6 (.CI(n31237), .I0(n1545), 
            .I1(GND_net), .CO(n31238));
    SB_LUT4 encoder0_position_23__I_0_add_1043_5_lut (.I0(GND_net), .I1(n1546), 
            .I2(VCC_net), .I3(n31236), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_5 (.CI(n31236), .I0(n1546), 
            .I1(VCC_net), .CO(n31237));
    SB_LUT4 i14018_3_lut (.I0(\data_in_frame[14] [5]), .I1(rx_data[5]), 
            .I2(n35562), .I3(GND_net), .O(n22421));   // verilog/coms.v(127[12] 300[6])
    defparam i14018_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_add_1043_4_lut (.I0(GND_net), .I1(n1547), 
            .I2(GND_net), .I3(n31235), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_644_23_lut (.I0(duty[21]), .I1(n40620), .I2(n4), .I3(n30760), 
            .O(pwm_setpoint_22__N_11[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_add_1043_4 (.CI(n31235), .I0(n1547), 
            .I1(GND_net), .CO(n31236));
    SB_LUT4 encoder0_position_23__I_0_add_1043_3_lut (.I0(GND_net), .I1(n1548), 
            .I2(VCC_net), .I3(n31234), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_1043_3 (.CI(n31234), .I0(n1548), 
            .I1(VCC_net), .CO(n31235));
    SB_CARRY add_644_23 (.CI(n30760), .I0(n40620), .I1(n4), .CO(n30761));
    SB_LUT4 encoder0_position_23__I_0_add_1043_2_lut (.I0(GND_net), .I1(n526), 
            .I2(GND_net), .I3(VCC_net), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_1043_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_644_22_lut (.I0(duty[20]), .I1(n40620), .I2(n5), .I3(n30759), 
            .O(pwm_setpoint_22__N_11[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_add_1043_2 (.CI(VCC_net), .I0(n526), 
            .I1(GND_net), .CO(n31234));
    SB_LUT4 i14440_3_lut (.I0(n22193), .I1(r_Bit_Index[0]), .I2(n22012), 
            .I3(GND_net), .O(n22843));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14440_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i14414_3_lut (.I0(n22195), .I1(r_Bit_Index_adj_5090[0]), .I2(n21920), 
            .I3(GND_net), .O(n22817));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i14414_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 i1_4_lut_adj_1727 (.I0(n27098), .I1(n35591), .I2(state_adj_5082[0]), 
            .I3(read), .O(n35254));   // verilog/eeprom.v(25[8] 57[4])
    defparam i1_4_lut_adj_1727.LUT_INIT = 16'h8280;
    SB_LUT4 encoder0_position_23__I_0_add_990_18_lut (.I0(GND_net), .I1(n1454), 
            .I2(VCC_net), .I3(n31233), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_644_22 (.CI(n30759), .I0(n40620), .I1(n5), .CO(n30760));
    SB_LUT4 encoder0_position_23__I_0_add_990_17_lut (.I0(GND_net), .I1(n1455), 
            .I2(VCC_net), .I3(n31232), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_644_21_lut (.I0(duty[19]), .I1(n40620), .I2(n6), .I3(n30758), 
            .O(pwm_setpoint_22__N_11[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_add_990_17 (.CI(n31232), .I0(n1455), 
            .I1(VCC_net), .CO(n31233));
    SB_LUT4 encoder0_position_23__I_0_add_990_16_lut (.I0(GND_net), .I1(n1456), 
            .I2(VCC_net), .I3(n31231), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_16 (.CI(n31231), .I0(n1456), 
            .I1(VCC_net), .CO(n31232));
    SB_CARRY add_644_21 (.CI(n30758), .I0(n40620), .I1(n6), .CO(n30759));
    SB_LUT4 encoder0_position_23__I_0_add_990_15_lut (.I0(GND_net), .I1(n1457), 
            .I2(VCC_net), .I3(n31230), .O(n1510)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_15 (.CI(n31230), .I0(n1457), 
            .I1(VCC_net), .CO(n31231));
    SB_LUT4 encoder0_position_23__I_0_add_990_14_lut (.I0(GND_net), .I1(n1458), 
            .I2(VCC_net), .I3(n31229), .O(n1511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_14 (.CI(n31229), .I0(n1458), 
            .I1(VCC_net), .CO(n31230));
    SB_LUT4 encoder0_position_23__I_0_add_990_13_lut (.I0(GND_net), .I1(n1459), 
            .I2(VCC_net), .I3(n31228), .O(n1512)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_13 (.CI(n31228), .I0(n1459), 
            .I1(VCC_net), .CO(n31229));
    SB_LUT4 encoder0_position_23__I_0_add_990_12_lut (.I0(GND_net), .I1(n1460), 
            .I2(VCC_net), .I3(n31227), .O(n1513)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_644_20_lut (.I0(duty[18]), .I1(n40620), .I2(n7), .I3(n30757), 
            .O(pwm_setpoint_22__N_11[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_add_990_12 (.CI(n31227), .I0(n1460), 
            .I1(VCC_net), .CO(n31228));
    SB_LUT4 encoder0_position_23__I_0_add_990_11_lut (.I0(GND_net), .I1(n1461), 
            .I2(VCC_net), .I3(n31226), .O(n1514)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_11 (.CI(n31226), .I0(n1461), 
            .I1(VCC_net), .CO(n31227));
    SB_LUT4 encoder0_position_23__I_0_add_990_10_lut (.I0(GND_net), .I1(n1462), 
            .I2(VCC_net), .I3(n31225), .O(n1515)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_716_i6_3_lut_3_lut (.I0(pwm_setpoint[2]), .I1(pwm_setpoint[3]), 
            .I2(pwm_counter[3]), .I3(GND_net), .O(n6_adj_4956));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_716_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10_adj_4960));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29293_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n39321));
    defparam i29293_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_716_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12_adj_4962));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_716_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8_adj_4958));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_23__I_0_add_990_10 (.CI(n31225), .I0(n1462), 
            .I1(VCC_net), .CO(n31226));
    SB_DFFESR delay_counter_1507__i13 (.Q(delay_counter[13]), .C(CLK_c), 
            .E(n21971), .D(n152), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 encoder0_position_23__I_0_add_990_9_lut (.I0(GND_net), .I1(n1463), 
            .I2(VCC_net), .I3(n31224), .O(n1516)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29307_2_lut_4_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[4]), .I3(pwm_setpoint[4]), .O(n39335));
    defparam i29307_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i26426_4_lut (.I0(n7_adj_5015), .I1(state_adj_5082[0]), .I2(n6_adj_5025), 
            .I3(state_adj_5111[0]), .O(n36440));
    defparam i26426_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i1_3_lut (.I0(state_adj_5082[1]), .I1(read), .I2(n35591), 
            .I3(GND_net), .O(n12_adj_4878));   // verilog/eeprom.v(25[8] 57[4])
    defparam i1_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 i1_4_lut_adj_1728 (.I0(n27098), .I1(n12_adj_4878), .I2(state_adj_5082[0]), 
            .I3(n35591), .O(n35272));   // verilog/eeprom.v(25[8] 57[4])
    defparam i1_4_lut_adj_1728.LUT_INIT = 16'h88a8;
    SB_CARRY encoder0_position_23__I_0_add_990_9 (.CI(n31224), .I0(n1463), 
            .I1(VCC_net), .CO(n31225));
    SB_LUT4 encoder0_position_23__I_0_add_990_8_lut (.I0(GND_net), .I1(n1464), 
            .I2(VCC_net), .I3(n31223), .O(n1517)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_8 (.CI(n31223), .I0(n1464), 
            .I1(VCC_net), .CO(n31224));
    SB_LUT4 encoder0_position_23__I_0_add_990_7_lut (.I0(GND_net), .I1(n1465), 
            .I2(GND_net), .I3(n31222), .O(n1518)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_7 (.CI(n31222), .I0(n1465), 
            .I1(GND_net), .CO(n31223));
    SB_LUT4 encoder0_position_23__I_0_add_990_6_lut (.I0(GND_net), .I1(n1466), 
            .I2(GND_net), .I3(n31221), .O(n1519)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_6 (.CI(n31221), .I0(n1466), 
            .I1(GND_net), .CO(n31222));
    SB_LUT4 encoder0_position_23__I_0_add_990_5_lut (.I0(GND_net), .I1(n1467), 
            .I2(VCC_net), .I3(n31220), .O(n1520)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_5 (.CI(n31220), .I0(n1467), 
            .I1(VCC_net), .CO(n31221));
    SB_LUT4 encoder0_position_23__I_0_add_990_4_lut (.I0(GND_net), .I1(n1468), 
            .I2(GND_net), .I3(n31219), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_4 (.CI(n31219), .I0(n1468), 
            .I1(GND_net), .CO(n31220));
    SB_CARRY add_644_20 (.CI(n30757), .I0(n40620), .I1(n7), .CO(n30758));
    SB_LUT4 encoder0_position_23__I_0_add_990_3_lut (.I0(GND_net), .I1(n1469), 
            .I2(VCC_net), .I3(n31218), .O(n1522)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_3 (.CI(n31218), .I0(n1469), 
            .I1(VCC_net), .CO(n31219));
    SB_LUT4 add_644_19_lut (.I0(duty[17]), .I1(n40620), .I2(n8), .I3(n30756), 
            .O(pwm_setpoint_22__N_11[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_990_2_lut (.I0(GND_net), .I1(n525), 
            .I2(GND_net), .I3(VCC_net), .O(n1523)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_990_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_990_2 (.CI(VCC_net), .I0(n525), 
            .I1(GND_net), .CO(n31218));
    SB_LUT4 encoder0_position_23__I_0_add_937_17_lut (.I0(GND_net), .I1(n1376), 
            .I2(VCC_net), .I3(n31217), .O(n1429)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_937_16_lut (.I0(GND_net), .I1(n1377), 
            .I2(VCC_net), .I3(n31216), .O(n1430)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_644_19 (.CI(n30756), .I0(n40620), .I1(n8), .CO(n30757));
    SB_CARRY encoder0_position_23__I_0_add_937_16 (.CI(n31216), .I0(n1377), 
            .I1(VCC_net), .CO(n31217));
    SB_LUT4 encoder0_position_23__I_0_add_937_15_lut (.I0(GND_net), .I1(n1378), 
            .I2(VCC_net), .I3(n31215), .O(n1431)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_15 (.CI(n31215), .I0(n1378), 
            .I1(VCC_net), .CO(n31216));
    SB_LUT4 encoder0_position_23__I_0_add_937_14_lut (.I0(GND_net), .I1(n1379), 
            .I2(VCC_net), .I3(n31214), .O(n1432)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_644_18_lut (.I0(duty[16]), .I1(n40620), .I2(n9), .I3(n30755), 
            .O(pwm_setpoint_22__N_11[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_add_937_14 (.CI(n31214), .I0(n1379), 
            .I1(VCC_net), .CO(n31215));
    SB_LUT4 encoder0_position_23__I_0_add_937_13_lut (.I0(GND_net), .I1(n1380), 
            .I2(VCC_net), .I3(n31213), .O(n1433)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_13 (.CI(n31213), .I0(n1380), 
            .I1(VCC_net), .CO(n31214));
    SB_LUT4 encoder0_position_23__I_0_add_937_12_lut (.I0(GND_net), .I1(n1381), 
            .I2(VCC_net), .I3(n31212), .O(n1434)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_12 (.CI(n31212), .I0(n1381), 
            .I1(VCC_net), .CO(n31213));
    SB_LUT4 encoder0_position_23__I_0_add_937_11_lut (.I0(GND_net), .I1(n1382), 
            .I2(VCC_net), .I3(n31211), .O(n1435)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_11 (.CI(n31211), .I0(n1382), 
            .I1(VCC_net), .CO(n31212));
    SB_LUT4 encoder0_position_23__I_0_add_937_10_lut (.I0(GND_net), .I1(n1383), 
            .I2(VCC_net), .I3(n31210), .O(n1436)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_10 (.CI(n31210), .I0(n1383), 
            .I1(VCC_net), .CO(n31211));
    SB_LUT4 encoder0_position_23__I_0_add_937_9_lut (.I0(GND_net), .I1(n1384), 
            .I2(VCC_net), .I3(n31209), .O(n1437)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_9 (.CI(n31209), .I0(n1384), 
            .I1(VCC_net), .CO(n31210));
    SB_DFFESR delay_counter_1507__i12 (.Q(delay_counter[12]), .C(CLK_c), 
            .E(n21971), .D(n153), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 encoder0_position_23__I_0_i1312_3_lut (.I0(n1924), .I1(n1977), 
            .I2(n1948), .I3(GND_net), .O(n2002));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_i1312_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_1507__i11 (.Q(delay_counter[11]), .C(CLK_c), 
            .E(n21971), .D(n154), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 encoder0_position_23__I_0_add_937_8_lut (.I0(GND_net), .I1(n1385), 
            .I2(VCC_net), .I3(n31208), .O(n1438)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_1507__i10 (.Q(delay_counter[10]), .C(CLK_c), 
            .E(n21971), .D(n155), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_CARRY encoder0_position_23__I_0_add_937_8 (.CI(n31208), .I0(n1385), 
            .I1(VCC_net), .CO(n31209));
    SB_LUT4 encoder0_position_23__I_0_add_937_7_lut (.I0(GND_net), .I1(n1386), 
            .I2(GND_net), .I3(n31207), .O(n1439)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_7 (.CI(n31207), .I0(n1386), 
            .I1(GND_net), .CO(n31208));
    SB_LUT4 encoder0_position_23__I_0_add_937_6_lut (.I0(GND_net), .I1(n1387), 
            .I2(GND_net), .I3(n31206), .O(n1440)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_1507__i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n21971), 
            .D(n156), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_CARRY encoder0_position_23__I_0_add_937_6 (.CI(n31206), .I0(n1387), 
            .I1(GND_net), .CO(n31207));
    SB_LUT4 encoder0_position_23__I_0_add_937_5_lut (.I0(GND_net), .I1(n1388), 
            .I2(VCC_net), .I3(n31205), .O(n1441)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_5 (.CI(n31205), .I0(n1388), 
            .I1(VCC_net), .CO(n31206));
    SB_LUT4 encoder0_position_23__I_0_add_937_4_lut (.I0(GND_net), .I1(n1389), 
            .I2(GND_net), .I3(n31204), .O(n1442)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_4 (.CI(n31204), .I0(n1389), 
            .I1(GND_net), .CO(n31205));
    SB_LUT4 encoder0_position_23__I_0_add_937_3_lut (.I0(GND_net), .I1(n1390), 
            .I2(VCC_net), .I3(n31203), .O(n1443)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_3 (.CI(n31203), .I0(n1390), 
            .I1(VCC_net), .CO(n31204));
    SB_LUT4 encoder0_position_23__I_0_add_937_2_lut (.I0(GND_net), .I1(n524), 
            .I2(GND_net), .I3(VCC_net), .O(n1444)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_937_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_937_2 (.CI(VCC_net), .I0(n524), 
            .I1(GND_net), .CO(n31203));
    SB_LUT4 encoder0_position_23__I_0_add_884_16_lut (.I0(GND_net), .I1(n1298), 
            .I2(VCC_net), .I3(n31202), .O(n1351)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_884_15_lut (.I0(GND_net), .I1(n1299), 
            .I2(VCC_net), .I3(n31201), .O(n1352)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_15 (.CI(n31201), .I0(n1299), 
            .I1(VCC_net), .CO(n31202));
    SB_LUT4 encoder0_position_23__I_0_add_884_14_lut (.I0(GND_net), .I1(n1300), 
            .I2(VCC_net), .I3(n31200), .O(n1353)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_14 (.CI(n31200), .I0(n1300), 
            .I1(VCC_net), .CO(n31201));
    SB_DFFESR delay_counter_1507__i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n21971), 
            .D(n157), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 encoder0_position_23__I_0_add_884_13_lut (.I0(GND_net), .I1(n1301), 
            .I2(VCC_net), .I3(n31199), .O(n1354)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_13 (.CI(n31199), .I0(n1301), 
            .I1(VCC_net), .CO(n31200));
    SB_LUT4 encoder0_position_23__I_0_add_884_12_lut (.I0(GND_net), .I1(n1302), 
            .I2(VCC_net), .I3(n31198), .O(n1355)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_644_18 (.CI(n30755), .I0(n40620), .I1(n9), .CO(n30756));
    SB_CARRY encoder0_position_23__I_0_add_884_12 (.CI(n31198), .I0(n1302), 
            .I1(VCC_net), .CO(n31199));
    SB_LUT4 add_644_17_lut (.I0(duty[15]), .I1(n40620), .I2(n10), .I3(n30754), 
            .O(pwm_setpoint_22__N_11[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_884_11_lut (.I0(GND_net), .I1(n1303), 
            .I2(VCC_net), .I3(n31197), .O(n1356)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_11 (.CI(n31197), .I0(n1303), 
            .I1(VCC_net), .CO(n31198));
    SB_LUT4 encoder0_position_23__I_0_add_884_10_lut (.I0(GND_net), .I1(n1304), 
            .I2(VCC_net), .I3(n31196), .O(n1357)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_10 (.CI(n31196), .I0(n1304), 
            .I1(VCC_net), .CO(n31197));
    SB_LUT4 encoder0_position_23__I_0_add_884_9_lut (.I0(GND_net), .I1(n1305), 
            .I2(VCC_net), .I3(n31195), .O(n1358)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1783_7_lut (.I0(GND_net), .I1(n509), .I2(GND_net), .I3(n32024), 
            .O(n5440)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1783_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1783_6_lut (.I0(n38316), .I1(n510), .I2(GND_net), .I3(n32023), 
            .O(n39289)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1783_6_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_1783_6 (.CI(n32023), .I0(n510), .I1(GND_net), .CO(n32024));
    SB_LUT4 add_1783_5_lut (.I0(GND_net), .I1(n511), .I2(VCC_net), .I3(n32022), 
            .O(n5442)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1783_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_9 (.CI(n31195), .I0(n1305), 
            .I1(VCC_net), .CO(n31196));
    SB_CARRY add_1783_5 (.CI(n32022), .I0(n511), .I1(VCC_net), .CO(n32023));
    SB_LUT4 encoder0_position_23__I_0_add_884_8_lut (.I0(GND_net), .I1(n1306), 
            .I2(VCC_net), .I3(n31194), .O(n1359)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1783_4_lut (.I0(GND_net), .I1(n425), .I2(GND_net), .I3(n32021), 
            .O(n5443)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1783_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_644_17 (.CI(n30754), .I0(n40620), .I1(n10), .CO(n30755));
    SB_CARRY add_1783_4 (.CI(n32021), .I0(n425), .I1(GND_net), .CO(n32022));
    SB_LUT4 add_1783_3_lut (.I0(GND_net), .I1(n513), .I2(VCC_net), .I3(n32020), 
            .O(n5444)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1783_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1783_3 (.CI(n32020), .I0(n513), .I1(VCC_net), .CO(n32021));
    SB_LUT4 add_1783_2_lut (.I0(GND_net), .I1(n514), .I2(GND_net), .I3(VCC_net), 
            .O(n5445)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1783_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_8 (.CI(n31194), .I0(n1306), 
            .I1(VCC_net), .CO(n31195));
    SB_CARRY add_1783_2 (.CI(VCC_net), .I0(n514), .I1(GND_net), .CO(n32020));
    SB_LUT4 encoder0_position_23__I_0_add_884_7_lut (.I0(GND_net), .I1(n1307), 
            .I2(GND_net), .I3(n31193), .O(n1360)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_7 (.CI(n31193), .I0(n1307), 
            .I1(GND_net), .CO(n31194));
    SB_LUT4 encoder0_position_23__I_0_add_884_6_lut (.I0(GND_net), .I1(n1308), 
            .I2(GND_net), .I3(n31192), .O(n1361)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_6 (.CI(n31192), .I0(n1308), 
            .I1(GND_net), .CO(n31193));
    SB_LUT4 encoder0_position_23__I_0_add_884_5_lut (.I0(GND_net), .I1(n1309), 
            .I2(VCC_net), .I3(n31191), .O(n1362)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_5 (.CI(n31191), .I0(n1309), 
            .I1(VCC_net), .CO(n31192));
    SB_LUT4 encoder0_position_23__I_0_add_884_4_lut (.I0(GND_net), .I1(n1310), 
            .I2(GND_net), .I3(n31190), .O(n1363)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_4 (.CI(n31190), .I0(n1310), 
            .I1(GND_net), .CO(n31191));
    SB_LUT4 encoder0_position_23__I_0_add_884_3_lut (.I0(GND_net), .I1(n1311), 
            .I2(VCC_net), .I3(n31189), .O(n1364)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_3 (.CI(n31189), .I0(n1311), 
            .I1(VCC_net), .CO(n31190));
    SB_LUT4 add_644_16_lut (.I0(duty[14]), .I1(n40620), .I2(n11), .I3(n30753), 
            .O(pwm_setpoint_22__N_11[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_644_16 (.CI(n30753), .I0(n40620), .I1(n11), .CO(n30754));
    SB_LUT4 encoder0_position_23__I_0_add_884_2_lut (.I0(GND_net), .I1(n523), 
            .I2(GND_net), .I3(VCC_net), .O(n1365)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_884_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_884_2 (.CI(VCC_net), .I0(n523), 
            .I1(GND_net), .CO(n31189));
    SB_LUT4 encoder0_position_23__I_0_add_831_15_lut (.I0(GND_net), .I1(n1220), 
            .I2(VCC_net), .I3(n31188), .O(n1273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4996));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13937_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n21865), .I3(GND_net), .O(n22340));   // verilog/coms.v(127[12] 300[6])
    defparam i13937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14019_3_lut (.I0(\data_in_frame[14] [4]), .I1(rx_data[4]), 
            .I2(n35562), .I3(GND_net), .O(n22422));   // verilog/coms.v(127[12] 300[6])
    defparam i14019_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13938_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n21865), .I3(GND_net), .O(n22341));   // verilog/coms.v(127[12] 300[6])
    defparam i13938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13939_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n21865), .I3(GND_net), .O(n22342));   // verilog/coms.v(127[12] 300[6])
    defparam i13939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13940_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n21865), .I3(GND_net), .O(n22343));   // verilog/coms.v(127[12] 300[6])
    defparam i13940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13941_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n21865), .I3(GND_net), .O(n22344));   // verilog/coms.v(127[12] 300[6])
    defparam i13941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30459_2_lut_3_lut (.I0(n3_adj_4904), .I1(n4_adj_5000), .I2(encoder0_position[23]), 
            .I3(GND_net), .O(n619));
    defparam i30459_2_lut_3_lut.LUT_INIT = 16'h7f7f;
    SB_LUT4 i26324_3_lut_4_lut (.I0(n3_adj_4904), .I1(n4_adj_5000), .I2(n5442), 
            .I3(n4_adj_4903), .O(n36334));
    defparam i26324_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i26356_3_lut_4_lut (.I0(n3_adj_4904), .I1(n4_adj_5000), .I2(n5444), 
            .I3(n6_adj_4899), .O(n36368));
    defparam i26356_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 encoder0_position_23__I_0_add_831_14_lut (.I0(GND_net), .I1(n1221), 
            .I2(VCC_net), .I3(n31187), .O(n1274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_14 (.CI(n31187), .I0(n1221), 
            .I1(VCC_net), .CO(n31188));
    SB_LUT4 encoder0_position_23__I_0_add_831_13_lut (.I0(GND_net), .I1(n1222), 
            .I2(VCC_net), .I3(n31186), .O(n1275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_13 (.CI(n31186), .I0(n1222), 
            .I1(VCC_net), .CO(n31187));
    SB_DFFESR delay_counter_1507__i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n21971), 
            .D(n158), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 encoder0_position_23__I_0_add_831_12_lut (.I0(GND_net), .I1(n1223), 
            .I2(VCC_net), .I3(n31185), .O(n1276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_12 (.CI(n31185), .I0(n1223), 
            .I1(VCC_net), .CO(n31186));
    SB_LUT4 encoder0_position_23__I_0_add_831_11_lut (.I0(GND_net), .I1(n1224), 
            .I2(VCC_net), .I3(n31184), .O(n1277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_11 (.CI(n31184), .I0(n1224), 
            .I1(VCC_net), .CO(n31185));
    SB_LUT4 encoder0_position_23__I_0_add_831_10_lut (.I0(GND_net), .I1(n1225), 
            .I2(VCC_net), .I3(n31183), .O(n1278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_10 (.CI(n31183), .I0(n1225), 
            .I1(VCC_net), .CO(n31184));
    SB_LUT4 encoder0_position_23__I_0_add_831_9_lut (.I0(GND_net), .I1(n1226), 
            .I2(VCC_net), .I3(n31182), .O(n1279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_9 (.CI(n31182), .I0(n1226), 
            .I1(VCC_net), .CO(n31183));
    SB_LUT4 add_644_15_lut (.I0(duty[13]), .I1(n40620), .I2(n12), .I3(n30752), 
            .O(pwm_setpoint_22__N_11[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_15_lut.LUT_INIT = 16'h8BB8;
    SB_DFFESR delay_counter_1507__i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n21971), 
            .D(n159), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 encoder0_position_23__I_0_add_831_8_lut (.I0(GND_net), .I1(n1227), 
            .I2(VCC_net), .I3(n31181), .O(n1280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_8 (.CI(n31181), .I0(n1227), 
            .I1(VCC_net), .CO(n31182));
    SB_LUT4 encoder0_position_23__I_0_add_831_7_lut (.I0(GND_net), .I1(n1228), 
            .I2(GND_net), .I3(n31180), .O(n1281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_7 (.CI(n31180), .I0(n1228), 
            .I1(GND_net), .CO(n31181));
    SB_LUT4 encoder0_position_23__I_0_add_831_6_lut (.I0(GND_net), .I1(n1229), 
            .I2(GND_net), .I3(n31179), .O(n1282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_6 (.CI(n31179), .I0(n1229), 
            .I1(GND_net), .CO(n31180));
    SB_LUT4 encoder0_position_23__I_0_add_831_5_lut (.I0(GND_net), .I1(n1230), 
            .I2(VCC_net), .I3(n31178), .O(n1283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_5 (.CI(n31178), .I0(n1230), 
            .I1(VCC_net), .CO(n31179));
    SB_LUT4 encoder0_position_23__I_0_add_831_4_lut (.I0(GND_net), .I1(n1231), 
            .I2(GND_net), .I3(n31177), .O(n1284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_4 (.CI(n31177), .I0(n1231), 
            .I1(GND_net), .CO(n31178));
    SB_LUT4 i26320_3_lut_4_lut (.I0(n3_adj_4904), .I1(n4_adj_5000), .I2(n5443), 
            .I3(n5_adj_4900), .O(n36330));
    defparam i26320_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 encoder0_position_23__I_0_add_831_3_lut (.I0(GND_net), .I1(n1232), 
            .I2(VCC_net), .I3(n31176), .O(n1285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_3 (.CI(n31176), .I0(n1232), 
            .I1(VCC_net), .CO(n31177));
    SB_LUT4 i26322_3_lut_4_lut (.I0(n3_adj_4904), .I1(n4_adj_5000), .I2(n5445), 
            .I3(n7_adj_4898), .O(n36332));
    defparam i26322_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 encoder0_position_23__I_0_i409_3_lut_4_lut (.I0(n2), .I1(encoder0_position[23]), 
            .I2(n619), .I3(n5440), .O(n674));
    defparam encoder0_position_23__I_0_i409_3_lut_4_lut.LUT_INIT = 16'h8f80;
    SB_LUT4 encoder0_position_23__I_0_add_831_2_lut (.I0(GND_net), .I1(n522), 
            .I2(GND_net), .I3(VCC_net), .O(n1286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_831_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_831_2 (.CI(VCC_net), .I0(n522), 
            .I1(GND_net), .CO(n31176));
    SB_LUT4 encoder0_position_23__I_0_add_778_14_lut (.I0(GND_net), .I1(n1142), 
            .I2(VCC_net), .I3(n31175), .O(n1195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_778_13_lut (.I0(GND_net), .I1(n1143), 
            .I2(VCC_net), .I3(n31174), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_13 (.CI(n31174), .I0(n1143), 
            .I1(VCC_net), .CO(n31175));
    SB_LUT4 encoder0_position_23__I_0_add_778_12_lut (.I0(GND_net), .I1(n1144), 
            .I2(VCC_net), .I3(n31173), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_12 (.CI(n31173), .I0(n1144), 
            .I1(VCC_net), .CO(n31174));
    SB_LUT4 encoder0_position_23__I_0_add_778_11_lut (.I0(GND_net), .I1(n1145), 
            .I2(VCC_net), .I3(n31172), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_11 (.CI(n31172), .I0(n1145), 
            .I1(VCC_net), .CO(n31173));
    SB_LUT4 encoder0_position_23__I_0_add_778_10_lut (.I0(GND_net), .I1(n1146), 
            .I2(VCC_net), .I3(n31171), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_10 (.CI(n31171), .I0(n1146), 
            .I1(VCC_net), .CO(n31172));
    SB_LUT4 encoder0_position_23__I_0_add_778_9_lut (.I0(GND_net), .I1(n1147), 
            .I2(VCC_net), .I3(n31170), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_9 (.CI(n31170), .I0(n1147), 
            .I1(VCC_net), .CO(n31171));
    SB_LUT4 encoder0_position_23__I_0_add_778_8_lut (.I0(GND_net), .I1(n1148), 
            .I2(VCC_net), .I3(n31169), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_8 (.CI(n31169), .I0(n1148), 
            .I1(VCC_net), .CO(n31170));
    SB_LUT4 encoder0_position_23__I_0_add_778_7_lut (.I0(GND_net), .I1(n1149), 
            .I2(GND_net), .I3(n31168), .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_7 (.CI(n31168), .I0(n1149), 
            .I1(GND_net), .CO(n31169));
    SB_LUT4 encoder0_position_23__I_0_add_778_6_lut (.I0(GND_net), .I1(n1150), 
            .I2(GND_net), .I3(n31167), .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_6 (.CI(n31167), .I0(n1150), 
            .I1(GND_net), .CO(n31168));
    SB_LUT4 encoder0_position_23__I_0_add_778_5_lut (.I0(GND_net), .I1(n1151), 
            .I2(VCC_net), .I3(n31166), .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_5 (.CI(n31166), .I0(n1151), 
            .I1(VCC_net), .CO(n31167));
    SB_LUT4 encoder0_position_23__I_0_add_778_4_lut (.I0(GND_net), .I1(n1152), 
            .I2(GND_net), .I3(n31165), .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_4 (.CI(n31165), .I0(n1152), 
            .I1(GND_net), .CO(n31166));
    SB_LUT4 encoder0_position_23__I_0_add_778_3_lut (.I0(GND_net), .I1(n1153), 
            .I2(VCC_net), .I3(n31164), .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_3 (.CI(n31164), .I0(n1153), 
            .I1(VCC_net), .CO(n31165));
    SB_LUT4 encoder0_position_23__I_0_add_778_2_lut (.I0(GND_net), .I1(n521), 
            .I2(GND_net), .I3(VCC_net), .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_778_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_778_2 (.CI(VCC_net), .I0(n521), 
            .I1(GND_net), .CO(n31164));
    SB_LUT4 encoder0_position_23__I_0_add_725_13_lut (.I0(GND_net), .I1(n1064), 
            .I2(VCC_net), .I3(n31163), .O(n1117)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_725_12_lut (.I0(GND_net), .I1(n1065), 
            .I2(VCC_net), .I3(n31162), .O(n1118)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_12 (.CI(n31162), .I0(n1065), 
            .I1(VCC_net), .CO(n31163));
    SB_LUT4 encoder0_position_23__I_0_add_725_11_lut (.I0(GND_net), .I1(n1066), 
            .I2(VCC_net), .I3(n31161), .O(n1119)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_11 (.CI(n31161), .I0(n1066), 
            .I1(VCC_net), .CO(n31162));
    SB_LUT4 encoder0_position_23__I_0_add_725_10_lut (.I0(GND_net), .I1(n1067), 
            .I2(VCC_net), .I3(n31160), .O(n1120)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_10 (.CI(n31160), .I0(n1067), 
            .I1(VCC_net), .CO(n31161));
    SB_LUT4 encoder0_position_23__I_0_add_725_9_lut (.I0(GND_net), .I1(n1068), 
            .I2(VCC_net), .I3(n31159), .O(n1121)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_9 (.CI(n31159), .I0(n1068), 
            .I1(VCC_net), .CO(n31160));
    SB_LUT4 encoder0_position_23__I_0_add_725_8_lut (.I0(GND_net), .I1(n1069), 
            .I2(VCC_net), .I3(n31158), .O(n1122)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_8 (.CI(n31158), .I0(n1069), 
            .I1(VCC_net), .CO(n31159));
    SB_LUT4 encoder0_position_23__I_0_add_725_7_lut (.I0(GND_net), .I1(n1070), 
            .I2(GND_net), .I3(n31157), .O(n1123)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_7 (.CI(n31157), .I0(n1070), 
            .I1(GND_net), .CO(n31158));
    SB_DFF ID_i0_i7 (.Q(ID[7]), .C(CLK_c), .D(n22856));   // verilog/TinyFPGA_B.v(233[10] 247[6])
    SB_DFF ID_i0_i6 (.Q(ID[6]), .C(CLK_c), .D(n22855));   // verilog/TinyFPGA_B.v(233[10] 247[6])
    SB_DFF ID_i0_i5 (.Q(ID[5]), .C(CLK_c), .D(n22854));   // verilog/TinyFPGA_B.v(233[10] 247[6])
    SB_DFF ID_i0_i4 (.Q(ID[4]), .C(CLK_c), .D(n22853));   // verilog/TinyFPGA_B.v(233[10] 247[6])
    SB_DFF ID_i0_i3 (.Q(ID[3]), .C(CLK_c), .D(n22852));   // verilog/TinyFPGA_B.v(233[10] 247[6])
    SB_DFF ID_i0_i2 (.Q(ID[2]), .C(CLK_c), .D(n22851));   // verilog/TinyFPGA_B.v(233[10] 247[6])
    SB_DFF ID_i0_i1 (.Q(ID[1]), .C(CLK_c), .D(n22850));   // verilog/TinyFPGA_B.v(233[10] 247[6])
    SB_LUT4 encoder0_position_23__I_0_add_725_6_lut (.I0(GND_net), .I1(n1071), 
            .I2(GND_net), .I3(n31156), .O(n1124)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_6 (.CI(n31156), .I0(n1071), 
            .I1(GND_net), .CO(n31157));
    SB_LUT4 encoder0_position_23__I_0_add_725_5_lut (.I0(GND_net), .I1(n1072), 
            .I2(VCC_net), .I3(n31155), .O(n1125)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_644_15 (.CI(n30752), .I0(n40620), .I1(n12), .CO(n30753));
    SB_LUT4 i13942_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n21865), .I3(GND_net), .O(n22345));   // verilog/coms.v(127[12] 300[6])
    defparam i13942_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_725_5 (.CI(n31155), .I0(n1072), 
            .I1(VCC_net), .CO(n31156));
    SB_LUT4 encoder0_position_23__I_0_add_725_4_lut (.I0(GND_net), .I1(n1073), 
            .I2(GND_net), .I3(n31154), .O(n1126)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_4 (.CI(n31154), .I0(n1073), 
            .I1(GND_net), .CO(n31155));
    SB_LUT4 encoder0_position_23__I_0_add_725_3_lut (.I0(GND_net), .I1(n1074), 
            .I2(VCC_net), .I3(n31153), .O(n1127)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_644_14_lut (.I0(duty[12]), .I1(n40620), .I2(n13), .I3(n30751), 
            .O(pwm_setpoint_22__N_11[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_add_725_3 (.CI(n31153), .I0(n1074), 
            .I1(VCC_net), .CO(n31154));
    SB_LUT4 encoder0_position_23__I_0_add_725_2_lut (.I0(GND_net), .I1(n520), 
            .I2(GND_net), .I3(VCC_net), .O(n1128)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_725_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_725_2 (.CI(VCC_net), .I0(n520), 
            .I1(GND_net), .CO(n31153));
    SB_LUT4 encoder0_position_23__I_0_add_672_12_lut (.I0(n40392), .I1(n986), 
            .I2(VCC_net), .I3(n31152), .O(n1064)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_23__I_0_add_672_11_lut (.I0(GND_net), .I1(n987), 
            .I2(VCC_net), .I3(n31151), .O(n1040)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_11 (.CI(n31151), .I0(n987), 
            .I1(VCC_net), .CO(n31152));
    SB_CARRY add_644_14 (.CI(n30751), .I0(n40620), .I1(n13), .CO(n30752));
    SB_LUT4 encoder0_position_23__I_0_add_672_10_lut (.I0(GND_net), .I1(n988), 
            .I2(VCC_net), .I3(n31150), .O(n1041)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_10 (.CI(n31150), .I0(n988), 
            .I1(VCC_net), .CO(n31151));
    SB_LUT4 encoder0_position_23__I_0_add_672_9_lut (.I0(GND_net), .I1(n989), 
            .I2(VCC_net), .I3(n31149), .O(n1042)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_9 (.CI(n31149), .I0(n989), 
            .I1(VCC_net), .CO(n31150));
    SB_LUT4 encoder0_position_23__I_0_add_672_8_lut (.I0(GND_net), .I1(n990), 
            .I2(VCC_net), .I3(n31148), .O(n1043)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_8 (.CI(n31148), .I0(n990), 
            .I1(VCC_net), .CO(n31149));
    SB_LUT4 encoder0_position_23__I_0_add_672_7_lut (.I0(GND_net), .I1(n991), 
            .I2(GND_net), .I3(n31147), .O(n1044)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_7 (.CI(n31147), .I0(n991), 
            .I1(GND_net), .CO(n31148));
    SB_LUT4 encoder0_position_23__I_0_add_672_6_lut (.I0(GND_net), .I1(n992), 
            .I2(GND_net), .I3(n31146), .O(n1045)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_6 (.CI(n31146), .I0(n992), 
            .I1(GND_net), .CO(n31147));
    SB_LUT4 encoder0_position_23__I_0_add_672_5_lut (.I0(GND_net), .I1(n993), 
            .I2(VCC_net), .I3(n31145), .O(n1046)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_5 (.CI(n31145), .I0(n993), 
            .I1(VCC_net), .CO(n31146));
    SB_LUT4 add_644_13_lut (.I0(duty[11]), .I1(n40620), .I2(n14_adj_4855), 
            .I3(n30750), .O(pwm_setpoint_22__N_11[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_13_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_add_672_4_lut (.I0(GND_net), .I1(n994), 
            .I2(GND_net), .I3(n31144), .O(n1047)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_4 (.CI(n31144), .I0(n994), 
            .I1(GND_net), .CO(n31145));
    SB_LUT4 encoder0_position_23__I_0_add_672_3_lut (.I0(GND_net), .I1(n995), 
            .I2(VCC_net), .I3(n31143), .O(n1048)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_644_13 (.CI(n30750), .I0(n40620), .I1(n14_adj_4855), 
            .CO(n30751));
    SB_CARRY encoder0_position_23__I_0_add_672_3 (.CI(n31143), .I0(n995), 
            .I1(VCC_net), .CO(n31144));
    SB_LUT4 encoder0_position_23__I_0_add_672_2_lut (.I0(GND_net), .I1(n519), 
            .I2(GND_net), .I3(VCC_net), .O(n1049)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_672_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_672_2 (.CI(VCC_net), .I0(n519), 
            .I1(GND_net), .CO(n31143));
    SB_LUT4 i1_2_lut_adj_1729 (.I0(n20602), .I1(pwm_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(n20604));
    defparam i1_2_lut_adj_1729.LUT_INIT = 16'heeee;
    SB_LUT4 i29299_4_lut (.I0(n27), .I1(n15_adj_4964), .I2(n13_adj_4963), 
            .I3(n11_adj_4961), .O(n39327));
    defparam i29299_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29591_4_lut (.I0(n9_adj_4959), .I1(n7_adj_4957), .I2(pwm_counter[2]), 
            .I3(pwm_setpoint[2]), .O(n39620));
    defparam i29591_4_lut.LUT_INIT = 16'heffe;
    SB_LUT4 encoder0_position_23__I_0_add_619_11_lut (.I0(GND_net), .I1(n908), 
            .I2(VCC_net), .I3(n31134), .O(n961)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_619_10_lut (.I0(GND_net), .I1(n909), 
            .I2(VCC_net), .I3(n31133), .O(n962)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_10 (.CI(n31133), .I0(n909), 
            .I1(VCC_net), .CO(n31134));
    SB_LUT4 encoder0_position_23__I_0_add_619_9_lut (.I0(GND_net), .I1(n910), 
            .I2(VCC_net), .I3(n31132), .O(n963)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_9 (.CI(n31132), .I0(n910), 
            .I1(VCC_net), .CO(n31133));
    SB_LUT4 i29764_4_lut (.I0(n15_adj_4964), .I1(n13_adj_4963), .I2(n11_adj_4961), 
            .I3(n39620), .O(n39793));
    defparam i29764_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i29762_4_lut (.I0(n21_adj_4967), .I1(n19_adj_4966), .I2(n17_adj_4965), 
            .I3(n39793), .O(n39791));
    defparam i29762_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 encoder0_position_23__I_0_add_619_8_lut (.I0(GND_net), .I1(n911), 
            .I2(VCC_net), .I3(n31131), .O(n964)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29301_4_lut (.I0(n27), .I1(n25_adj_4969), .I2(n23_adj_4968), 
            .I3(n39791), .O(n39329));
    defparam i29301_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY encoder0_position_23__I_0_add_619_8 (.CI(n31131), .I0(n911), 
            .I1(VCC_net), .CO(n31132));
    SB_LUT4 encoder0_position_23__I_0_add_619_7_lut (.I0(GND_net), .I1(n912), 
            .I2(GND_net), .I3(n31130), .O(n965)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_716_i4_4_lut (.I0(pwm_setpoint[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_counter[0]), .O(n4_adj_4955));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i29913_3_lut (.I0(n4_adj_4955), .I1(pwm_setpoint[13]), .I2(n27), 
            .I3(GND_net), .O(n39942));   // verilog/pwm.v(21[8:24])
    defparam i29913_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_619_7 (.CI(n31130), .I0(n912), 
            .I1(GND_net), .CO(n31131));
    SB_LUT4 encoder0_position_23__I_0_add_619_6_lut (.I0(GND_net), .I1(n913), 
            .I2(GND_net), .I3(n31129), .O(n966)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_6 (.CI(n31129), .I0(n913), 
            .I1(GND_net), .CO(n31130));
    SB_LUT4 encoder0_position_23__I_0_add_619_5_lut (.I0(GND_net), .I1(n914), 
            .I2(VCC_net), .I3(n31128), .O(n967)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_5 (.CI(n31128), .I0(n914), 
            .I1(VCC_net), .CO(n31129));
    SB_LUT4 LessThan_716_i30_3_lut (.I0(n12_adj_4962), .I1(pwm_setpoint[17]), 
            .I2(n35), .I3(GND_net), .O(n30_adj_4970));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_619_4_lut (.I0(GND_net), .I1(n915), 
            .I2(GND_net), .I3(n31127), .O(n968)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29914_3_lut (.I0(n39942), .I1(pwm_setpoint[14]), .I2(n29), 
            .I3(GND_net), .O(n39943));   // verilog/pwm.v(21[8:24])
    defparam i29914_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29295_4_lut (.I0(n33_adj_4972), .I1(n31_adj_4971), .I2(n29), 
            .I3(n39327), .O(n39323));
    defparam i29295_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY encoder0_position_23__I_0_add_619_4 (.CI(n31127), .I0(n915), 
            .I1(GND_net), .CO(n31128));
    SB_LUT4 encoder0_position_23__I_0_add_619_3_lut (.I0(GND_net), .I1(n916), 
            .I2(VCC_net), .I3(n31126), .O(n969)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30025_4_lut (.I0(n30_adj_4970), .I1(n10_adj_4960), .I2(n35), 
            .I3(n39321), .O(n40054));   // verilog/pwm.v(21[8:24])
    defparam i30025_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29897_3_lut (.I0(n39943), .I1(pwm_setpoint[15]), .I2(n31_adj_4971), 
            .I3(GND_net), .O(n39926));   // verilog/pwm.v(21[8:24])
    defparam i29897_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_619_3 (.CI(n31126), .I0(n916), 
            .I1(VCC_net), .CO(n31127));
    SB_LUT4 encoder0_position_23__I_0_add_619_2_lut (.I0(GND_net), .I1(n518), 
            .I2(GND_net), .I3(VCC_net), .O(n970)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_619_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_619_2 (.CI(VCC_net), .I0(n518), 
            .I1(GND_net), .CO(n31126));
    SB_LUT4 i29915_3_lut (.I0(n6_adj_4956), .I1(pwm_setpoint[10]), .I2(n21_adj_4967), 
            .I3(GND_net), .O(n39944));   // verilog/pwm.v(21[8:24])
    defparam i29915_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_566_10_lut (.I0(GND_net), .I1(n830), 
            .I2(VCC_net), .I3(n31125), .O(n883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_add_566_9_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n31124), .O(n884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29916_3_lut (.I0(n39944), .I1(pwm_setpoint[11]), .I2(n23_adj_4968), 
            .I3(GND_net), .O(n39945));   // verilog/pwm.v(21[8:24])
    defparam i29916_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29581_4_lut (.I0(n23_adj_4968), .I1(n21_adj_4967), .I2(n19_adj_4966), 
            .I3(n39335), .O(n39610));
    defparam i29581_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i29832_3_lut (.I0(n8_adj_4958), .I1(pwm_setpoint[9]), .I2(n19_adj_4966), 
            .I3(GND_net), .O(n39861));   // verilog/pwm.v(21[8:24])
    defparam i29832_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_23__I_0_add_566_9 (.CI(n31124), .I0(n831), 
            .I1(VCC_net), .CO(n31125));
    SB_LUT4 i29895_3_lut (.I0(n39945), .I1(pwm_setpoint[12]), .I2(n25_adj_4969), 
            .I3(GND_net), .O(n39924));   // verilog/pwm.v(21[8:24])
    defparam i29895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29846_4_lut (.I0(n33_adj_4972), .I1(n31_adj_4971), .I2(n29), 
            .I3(n39329), .O(n39875));
    defparam i29846_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_23__I_0_add_566_8_lut (.I0(GND_net), .I1(n832), 
            .I2(VCC_net), .I3(n31123), .O(n885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30076_4_lut (.I0(n39926), .I1(n40054), .I2(n35), .I3(n39323), 
            .O(n40105));   // verilog/pwm.v(21[8:24])
    defparam i30076_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_23__I_0_add_566_8 (.CI(n31123), .I0(n832), 
            .I1(VCC_net), .CO(n31124));
    SB_LUT4 i29909_4_lut (.I0(n39924), .I1(n39861), .I2(n25_adj_4969), 
            .I3(n39610), .O(n39938));   // verilog/pwm.v(21[8:24])
    defparam i29909_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i30080_4_lut (.I0(n39938), .I1(n40105), .I2(n35), .I3(n39875), 
            .O(n40109));   // verilog/pwm.v(21[8:24])
    defparam i30080_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_23__I_0_add_566_7_lut (.I0(GND_net), .I1(n833), 
            .I2(GND_net), .I3(n31122), .O(n886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_7 (.CI(n31122), .I0(n833), 
            .I1(GND_net), .CO(n31123));
    SB_LUT4 encoder0_position_23__I_0_add_566_6_lut (.I0(GND_net), .I1(n834), 
            .I2(GND_net), .I3(n31121), .O(n887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30081_3_lut (.I0(n40109), .I1(pwm_setpoint[18]), .I2(pwm_counter[18]), 
            .I3(GND_net), .O(n40110));   // verilog/pwm.v(21[8:24])
    defparam i30081_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_23__I_0_add_566_6 (.CI(n31121), .I0(n834), 
            .I1(GND_net), .CO(n31122));
    SB_LUT4 encoder0_position_23__I_0_add_566_5_lut (.I0(GND_net), .I1(n835), 
            .I2(VCC_net), .I3(n31120), .O(n888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_5 (.CI(n31120), .I0(n835), 
            .I1(VCC_net), .CO(n31121));
    SB_LUT4 encoder0_position_23__I_0_add_566_4_lut (.I0(GND_net), .I1(n836), 
            .I2(GND_net), .I3(n31119), .O(n889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_4 (.CI(n31119), .I0(n836), 
            .I1(GND_net), .CO(n31120));
    SB_LUT4 encoder0_position_23__I_0_add_566_3_lut (.I0(GND_net), .I1(n837), 
            .I2(VCC_net), .I3(n31118), .O(n890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_3 (.CI(n31118), .I0(n837), 
            .I1(VCC_net), .CO(n31119));
    SB_LUT4 encoder0_position_23__I_0_add_566_2_lut (.I0(GND_net), .I1(n517), 
            .I2(GND_net), .I3(VCC_net), .O(n891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_566_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_566_2 (.CI(VCC_net), .I0(n517), 
            .I1(GND_net), .CO(n31118));
    SB_LUT4 i30079_3_lut (.I0(n40110), .I1(pwm_setpoint[19]), .I2(pwm_counter[19]), 
            .I3(GND_net), .O(n40108));   // verilog/pwm.v(21[8:24])
    defparam i30079_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_23__I_0_add_513_9_lut (.I0(n40353), .I1(n752), 
            .I2(VCC_net), .I3(n31117), .O(n830)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_23__I_0_add_513_8_lut (.I0(GND_net), .I1(n753), 
            .I2(VCC_net), .I3(n31116), .O(n806)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_513_8 (.CI(n31116), .I0(n753), 
            .I1(VCC_net), .CO(n31117));
    SB_LUT4 encoder0_position_23__I_0_add_513_7_lut (.I0(GND_net), .I1(n754), 
            .I2(GND_net), .I3(n31115), .O(n807)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_513_7 (.CI(n31115), .I0(n754), 
            .I1(GND_net), .CO(n31116));
    SB_LUT4 encoder0_position_23__I_0_add_513_6_lut (.I0(GND_net), .I1(n755), 
            .I2(GND_net), .I3(n31114), .O(n808)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30005_3_lut (.I0(n40108), .I1(pwm_setpoint[20]), .I2(pwm_counter[20]), 
            .I3(GND_net), .O(n40034));   // verilog/pwm.v(21[8:24])
    defparam i30005_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_23__I_0_add_513_6 (.CI(n31114), .I0(n755), 
            .I1(GND_net), .CO(n31115));
    SB_LUT4 encoder0_position_23__I_0_add_513_5_lut (.I0(GND_net), .I1(n756), 
            .I2(VCC_net), .I3(n31113), .O(n809)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_513_5 (.CI(n31113), .I0(n756), 
            .I1(VCC_net), .CO(n31114));
    SB_LUT4 encoder0_position_23__I_0_add_513_4_lut (.I0(GND_net), .I1(n757), 
            .I2(GND_net), .I3(n31112), .O(n810)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_513_4 (.CI(n31112), .I0(n757), 
            .I1(GND_net), .CO(n31113));
    SB_LUT4 encoder0_position_23__I_0_add_513_3_lut (.I0(GND_net), .I1(n758), 
            .I2(VCC_net), .I3(n31111), .O(n811)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_513_3 (.CI(n31111), .I0(n758), 
            .I1(VCC_net), .CO(n31112));
    SB_LUT4 encoder0_position_23__I_0_add_513_2_lut (.I0(GND_net), .I1(n516), 
            .I2(GND_net), .I3(VCC_net), .O(n812)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_513_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_513_2 (.CI(VCC_net), .I0(n516), 
            .I1(GND_net), .CO(n31111));
    SB_LUT4 encoder0_position_23__I_0_add_460_8_lut (.I0(n40291), .I1(n674), 
            .I2(VCC_net), .I3(n31110), .O(n752)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_23__I_0_add_460_7_lut (.I0(GND_net), .I1(n675), 
            .I2(GND_net), .I3(n31109), .O(n728)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_460_7 (.CI(n31109), .I0(n675), 
            .I1(GND_net), .CO(n31110));
    SB_LUT4 encoder0_position_23__I_0_add_460_6_lut (.I0(GND_net), .I1(n676), 
            .I2(GND_net), .I3(n31108), .O(n729)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_460_6 (.CI(n31108), .I0(n676), 
            .I1(GND_net), .CO(n31109));
    SB_LUT4 encoder0_position_23__I_0_add_460_5_lut (.I0(GND_net), .I1(n677), 
            .I2(VCC_net), .I3(n31107), .O(n730)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_644_12_lut (.I0(duty[10]), .I1(n40620), .I2(n15_adj_4856), 
            .I3(n30749), .O(pwm_setpoint_22__N_11[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_23__I_0_add_460_5 (.CI(n31107), .I0(n677), 
            .I1(VCC_net), .CO(n31108));
    SB_LUT4 encoder0_position_23__I_0_add_460_4_lut (.I0(GND_net), .I1(n678), 
            .I2(GND_net), .I3(n31106), .O(n731)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_add_460_4 (.CI(n31106), .I0(n678), 
            .I1(GND_net), .CO(n31107));
    SB_LUT4 encoder0_position_23__I_0_add_460_3_lut (.I0(GND_net), .I1(n679), 
            .I2(VCC_net), .I3(n31105), .O(n732)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13943_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n21865), .I3(GND_net), .O(n22346));   // verilog/coms.v(127[12] 300[6])
    defparam i13943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13944_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n21865), .I3(GND_net), .O(n22347));   // verilog/coms.v(127[12] 300[6])
    defparam i13944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13945_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n21865), .I3(GND_net), .O(n22348));   // verilog/coms.v(127[12] 300[6])
    defparam i13945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13946_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n21865), .I3(GND_net), .O(n22349));   // verilog/coms.v(127[12] 300[6])
    defparam i13946_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_1507__i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n21971), 
            .D(n160), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_CARRY encoder0_position_23__I_0_add_460_3 (.CI(n31105), .I0(n679), 
            .I1(VCC_net), .CO(n31106));
    SB_LUT4 i13947_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n21865), .I3(GND_net), .O(n22350));   // verilog/coms.v(127[12] 300[6])
    defparam i13947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13948_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n21865), .I3(GND_net), .O(n22351));   // verilog/coms.v(127[12] 300[6])
    defparam i13948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13949_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n21865), .I3(GND_net), .O(n22352));   // verilog/coms.v(127[12] 300[6])
    defparam i13949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13950_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n21865), .I3(GND_net), .O(n22353));   // verilog/coms.v(127[12] 300[6])
    defparam i13950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13951_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n21865), .I3(GND_net), .O(n22354));   // verilog/coms.v(127[12] 300[6])
    defparam i13951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13952_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n21865), .I3(GND_net), .O(n22355));   // verilog/coms.v(127[12] 300[6])
    defparam i13952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13953_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n21865), .I3(GND_net), .O(n22356));   // verilog/coms.v(127[12] 300[6])
    defparam i13953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13954_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n21865), .I3(GND_net), .O(n22357));   // verilog/coms.v(127[12] 300[6])
    defparam i13954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13955_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n21865), .I3(GND_net), .O(n22358));   // verilog/coms.v(127[12] 300[6])
    defparam i13955_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_1507__i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n21971), 
            .D(n161), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 i13956_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n21865), .I3(GND_net), .O(n22359));   // verilog/coms.v(127[12] 300[6])
    defparam i13956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13957_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n21865), .I3(GND_net), .O(n22360));   // verilog/coms.v(127[12] 300[6])
    defparam i13957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13958_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n21865), .I3(GND_net), .O(n22361));   // verilog/coms.v(127[12] 300[6])
    defparam i13958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_23__I_0_add_460_2_lut (.I0(GND_net), .I1(n515), 
            .I2(GND_net), .I3(VCC_net), .O(n733)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_add_460_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_1507__i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n21971), 
            .D(n162), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_CARRY encoder0_position_23__I_0_add_460_2 (.CI(VCC_net), .I0(n515), 
            .I1(GND_net), .CO(n31105));
    SB_DFFESR delay_counter_1507__i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n21971), 
            .D(n163), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 i13959_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n21865), .I3(GND_net), .O(n22362));   // verilog/coms.v(127[12] 300[6])
    defparam i13959_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_1507__i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n21971), 
            .D(n164), .R(n22157));   // verilog/TinyFPGA_B.v(236[24:41])
    SB_LUT4 i13960_3_lut (.I0(\data_in_frame[21] [7]), .I1(rx_data[7]), 
            .I2(n35575), .I3(GND_net), .O(n22363));   // verilog/coms.v(127[12] 300[6])
    defparam i13960_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13961_3_lut (.I0(\data_in_frame[21] [6]), .I1(rx_data[6]), 
            .I2(n35575), .I3(GND_net), .O(n22364));   // verilog/coms.v(127[12] 300[6])
    defparam i13961_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13962_3_lut (.I0(\data_in_frame[21] [5]), .I1(rx_data[5]), 
            .I2(n35575), .I3(GND_net), .O(n22365));   // verilog/coms.v(127[12] 300[6])
    defparam i13962_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13963_3_lut (.I0(\data_in_frame[21] [4]), .I1(rx_data[4]), 
            .I2(n35575), .I3(GND_net), .O(n22366));   // verilog/coms.v(127[12] 300[6])
    defparam i13963_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13964_3_lut (.I0(\data_in_frame[21] [3]), .I1(rx_data[3]), 
            .I2(n35575), .I3(GND_net), .O(n22367));   // verilog/coms.v(127[12] 300[6])
    defparam i13964_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13965_3_lut (.I0(\data_in_frame[21] [2]), .I1(rx_data[2]), 
            .I2(n35575), .I3(GND_net), .O(n22368));   // verilog/coms.v(127[12] 300[6])
    defparam i13965_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13966_3_lut (.I0(\data_in_frame[21] [1]), .I1(rx_data[1]), 
            .I2(n35575), .I3(GND_net), .O(n22369));   // verilog/coms.v(127[12] 300[6])
    defparam i13966_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i30006_3_lut (.I0(n40034), .I1(pwm_setpoint[21]), .I2(pwm_counter[21]), 
            .I3(GND_net), .O(n40035));   // verilog/pwm.v(21[8:24])
    defparam i30006_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_644_12 (.CI(n30749), .I0(n40620), .I1(n15_adj_4856), 
            .CO(n30750));
    SB_LUT4 i13967_3_lut (.I0(\data_in_frame[21] [0]), .I1(rx_data[0]), 
            .I2(n35575), .I3(GND_net), .O(n22370));   // verilog/coms.v(127[12] 300[6])
    defparam i13967_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_644_11_lut (.I0(duty[9]), .I1(n40620), .I2(n16), .I3(n30748), 
            .O(pwm_setpoint_22__N_11[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_644_11 (.CI(n30748), .I0(n40620), .I1(n16), .CO(n30749));
    SB_LUT4 add_644_10_lut (.I0(duty[8]), .I1(n40620), .I2(n17), .I3(n30747), 
            .O(pwm_setpoint_22__N_11[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_10_lut.LUT_INIT = 16'h8BB8;
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(clk32MHz), 
           .D(encoder0_position_scaled_23__N_34[0]));   // verilog/TinyFPGA_B.v(200[10] 203[6])
    SB_DFF read_51 (.Q(read), .C(CLK_c), .D(n37894));   // verilog/TinyFPGA_B.v(233[10] 247[6])
    SB_DFF ID_i0_i0 (.Q(ID[0]), .C(CLK_c), .D(n22322));   // verilog/TinyFPGA_B.v(233[10] 247[6])
    SB_LUT4 LessThan_716_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4959));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i9_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_644_10 (.CI(n30747), .I0(n40620), .I1(n17), .CO(n30748));
    SB_LUT4 LessThan_716_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4961));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_716_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4965));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_716_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_716_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4964));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_644_9_lut (.I0(duty[7]), .I1(n40620), .I2(n18), .I3(n30746), 
            .O(pwm_setpoint_22__N_11[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 LessThan_716_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4963));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_716_i7_2_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4957));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_716_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4967));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_716_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4968));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_716_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4966));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_716_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i29_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_644_9 (.CI(n30746), .I0(n40620), .I1(n18), .CO(n30747));
    SB_LUT4 LessThan_716_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4971));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_716_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4972));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_4_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_716_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4969));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_716_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam LessThan_716_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_644_8_lut (.I0(duty[6]), .I1(n40620), .I2(n19), .I3(n30745), 
            .O(pwm_setpoint_22__N_11[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_644_8 (.CI(n30745), .I0(n40620), .I1(n19), .CO(n30746));
    SB_LUT4 add_644_7_lut (.I0(duty[5]), .I1(n40620), .I2(n20), .I3(n30744), 
            .O(pwm_setpoint_22__N_11[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 mux_3255_i20_3_lut (.I0(encoder0_position[19]), .I1(n6_adj_4899), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n513));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3255_i21_3_lut (.I0(encoder0_position[20]), .I1(n5_adj_4900), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n425));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_3255_i22_3_lut (.I0(encoder0_position[21]), .I1(n4_adj_4903), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n511));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28289_1_lut (.I0(n4_adj_5000), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n38316));
    defparam i28289_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_3255_i23_3_lut (.I0(encoder0_position[22]), .I1(n3_adj_4904), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n510));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam mux_3255_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_644_7 (.CI(n30744), .I0(n40620), .I1(n20), .CO(n30745));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4994));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_644_6_lut (.I0(duty[4]), .I1(n40620), .I2(n21), .I3(n30743), 
            .O(pwm_setpoint_22__N_11[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4993));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    GND i1 (.Y(GND_net));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4992));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4991));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13888_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n37680), .I3(GND_net), .O(n22291));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13888_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4990));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    motorControl control (.GND_net(GND_net), .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), 
            .\Ki[11] (Ki[11]), .\Kp[14] (Kp[14]), .PWMLimit({PWMLimit}), 
            .\Kp[15] (Kp[15]), .\Ki[12] (Ki[12]), .\Kp[9] (Kp[9]), .\Kp[10] (Kp[10]), 
            .\Ki[2] (Ki[2]), .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), 
            .\Kp[7] (Kp[7]), .\Ki[1] (Ki[1]), .\Ki[0] (Ki[0]), .\Kp[11] (Kp[11]), 
            .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), 
            .\Ki[7] (Ki[7]), .\Ki[8] (Ki[8]), .\Kp[1] (Kp[1]), .\Kp[0] (Kp[0]), 
            .\Kp[2] (Kp[2]), .\Kp[12] (Kp[12]), .\Kp[3] (Kp[3]), .\Kp[13] (Kp[13]), 
            .\Kp[8] (Kp[8]), .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), .IntegralLimit({IntegralLimit}), 
            .\Kp[6] (Kp[6]), .duty({duty}), .clk32MHz(clk32MHz), .VCC_net(VCC_net), 
            .setpoint({setpoint}), .motor_state({motor_state}), .n40620(n40620)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(170[16] 182[4])
    SB_LUT4 i14021_3_lut (.I0(\data_in_frame[14] [2]), .I1(rx_data[2]), 
            .I2(n35562), .I3(GND_net), .O(n22424));   // verilog/coms.v(127[12] 300[6])
    defparam i14021_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_644_6 (.CI(n30743), .I0(n40620), .I1(n21), .CO(n30744));
    SB_LUT4 add_644_5_lut (.I0(duty[3]), .I1(n40620), .I2(n22), .I3(n30742), 
            .O(pwm_setpoint_22__N_11[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_644_5_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_4976), .I3(n31816), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_4977), .I3(n31815), .O(n3_adj_4904)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4989));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_25 (.CI(n31815), 
            .I0(GND_net), .I1(n3_adj_4977), .CO(n31816));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4988));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_4978), .I3(n31814), .O(n4_adj_4903)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_24 (.CI(n31814), 
            .I0(GND_net), .I1(n4_adj_4978), .CO(n31815));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_4979), .I3(n31813), .O(n5_adj_4900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_23 (.CI(n31813), 
            .I0(GND_net), .I1(n5_adj_4979), .CO(n31814));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_4980), .I3(n31812), .O(n6_adj_4899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_22 (.CI(n31812), 
            .I0(GND_net), .I1(n6_adj_4980), .CO(n31813));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_4981), .I3(n31811), .O(n7_adj_4898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_21 (.CI(n31811), 
            .I0(GND_net), .I1(n7_adj_4981), .CO(n31812));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_4982), .I3(n31810), .O(n8_adj_4897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_20 (.CI(n31810), 
            .I0(GND_net), .I1(n8_adj_4982), .CO(n31811));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_4983), .I3(n31809), .O(n9_adj_4896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_19 (.CI(n31809), 
            .I0(GND_net), .I1(n9_adj_4983), .CO(n31810));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_4984), .I3(n31808), .O(n10_adj_4895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14022_3_lut (.I0(\data_in_frame[14] [1]), .I1(rx_data[1]), 
            .I2(n35562), .I3(GND_net), .O(n22425));   // verilog/coms.v(127[12] 300[6])
    defparam i14022_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4987));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4986));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_18 (.CI(n31808), 
            .I0(GND_net), .I1(n10_adj_4984), .CO(n31809));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_4985), .I3(n31807), .O(n11_adj_4894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_17 (.CI(n31807), 
            .I0(GND_net), .I1(n11_adj_4985), .CO(n31808));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_4986), .I3(n31806), .O(n12_adj_4893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_16 (.CI(n31806), 
            .I0(GND_net), .I1(n12_adj_4986), .CO(n31807));
    SB_CARRY add_644_5 (.CI(n30742), .I0(n40620), .I1(n22), .CO(n30743));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_4987), .I3(n31805), .O(n13_adj_4892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4985));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_15 (.CI(n31805), 
            .I0(GND_net), .I1(n13_adj_4987), .CO(n31806));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_4988), .I3(n31804), .O(n14_adj_4891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_14 (.CI(n31804), 
            .I0(GND_net), .I1(n14_adj_4988), .CO(n31805));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_4989), .I3(n31803), .O(n15_adj_4890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_13 (.CI(n31803), 
            .I0(GND_net), .I1(n15_adj_4989), .CO(n31804));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_4990), .I3(n31802), .O(n16_adj_4889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4984));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_12 (.CI(n31802), 
            .I0(GND_net), .I1(n16_adj_4990), .CO(n31803));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_4991), .I3(n31801), .O(n17_adj_4888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_11 (.CI(n31801), 
            .I0(GND_net), .I1(n17_adj_4991), .CO(n31802));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_4992), .I3(n31800), .O(n18_adj_4887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_10 (.CI(n31800), 
            .I0(GND_net), .I1(n18_adj_4992), .CO(n31801));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_4993), .I3(n31799), .O(n19_adj_4886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_9 (.CI(n31799), 
            .I0(GND_net), .I1(n19_adj_4993), .CO(n31800));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_4994), .I3(n31798), .O(n20_adj_4885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_23__I_0_unary_minus_2_add_3_8 (.CI(n31798), 
            .I0(GND_net), .I1(n20_adj_4994), .CO(n31799));
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_4995), .I3(n31797), .O(n21_adj_4884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_23__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4983));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4982));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4981));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4980));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14023_3_lut (.I0(\data_in_frame[14] [0]), .I1(rx_data[0]), 
            .I2(n35562), .I3(GND_net), .O(n22426));   // verilog/coms.v(127[12] 300[6])
    defparam i14023_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14024_3_lut (.I0(\data_in_frame[13] [7]), .I1(rx_data[7]), 
            .I2(n35568), .I3(GND_net), .O(n22427));   // verilog/coms.v(127[12] 300[6])
    defparam i14024_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4979));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14025_3_lut (.I0(\data_in_frame[13] [6]), .I1(rx_data[6]), 
            .I2(n35568), .I3(GND_net), .O(n22428));   // verilog/coms.v(127[12] 300[6])
    defparam i14025_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4978));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_23__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4977));   // verilog/TinyFPGA_B.v(201[33:55])
    defparam encoder0_position_23__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14026_3_lut (.I0(\data_in_frame[13] [5]), .I1(rx_data[5]), 
            .I2(n35568), .I3(GND_net), .O(n22429));   // verilog/coms.v(127[12] 300[6])
    defparam i14026_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14027_3_lut (.I0(\data_in_frame[13] [4]), .I1(rx_data[4]), 
            .I2(n35568), .I3(GND_net), .O(n22430));   // verilog/coms.v(127[12] 300[6])
    defparam i14027_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14028_3_lut (.I0(\data_in_frame[13] [3]), .I1(rx_data[3]), 
            .I2(n35568), .I3(GND_net), .O(n22431));   // verilog/coms.v(127[12] 300[6])
    defparam i14028_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14029_3_lut (.I0(\data_in_frame[13] [2]), .I1(rx_data[2]), 
            .I2(n35568), .I3(GND_net), .O(n22432));   // verilog/coms.v(127[12] 300[6])
    defparam i14029_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14030_3_lut (.I0(\data_in_frame[13] [1]), .I1(rx_data[1]), 
            .I2(n35568), .I3(GND_net), .O(n22433));   // verilog/coms.v(127[12] 300[6])
    defparam i14030_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14031_3_lut (.I0(\data_in_frame[13] [0]), .I1(rx_data[0]), 
            .I2(n35568), .I3(GND_net), .O(n22434));   // verilog/coms.v(127[12] 300[6])
    defparam i14031_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16_4_lut_4_lut (.I0(state_adj_5111[0]), .I1(n39285), .I2(n4760), 
            .I3(n10_adj_4908), .O(n8_adj_4879));   // verilog/i2c_controller.v(89[8] 155[6])
    defparam i16_4_lut_4_lut.LUT_INIT = 16'h3a7a;
    SB_LUT4 i29903_3_lut (.I0(n40035), .I1(pwm_setpoint[22]), .I2(pwm_counter[22]), 
            .I3(GND_net), .O(n39932));   // verilog/pwm.v(21[8:24])
    defparam i29903_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_4_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14072_3_lut (.I0(\data_in_frame[7] [7]), .I1(rx_data[7]), .I2(n35586), 
            .I3(GND_net), .O(n22475));   // verilog/coms.v(127[12] 300[6])
    defparam i14072_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14073_3_lut (.I0(\data_in_frame[7] [6]), .I1(rx_data[6]), .I2(n35586), 
            .I3(GND_net), .O(n22476));   // verilog/coms.v(127[12] 300[6])
    defparam i14073_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14074_3_lut (.I0(\data_in_frame[7] [5]), .I1(rx_data[5]), .I2(n35586), 
            .I3(GND_net), .O(n22477));   // verilog/coms.v(127[12] 300[6])
    defparam i14074_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14075_3_lut (.I0(\data_in_frame[7] [4]), .I1(rx_data[4]), .I2(n35586), 
            .I3(GND_net), .O(n22478));   // verilog/coms.v(127[12] 300[6])
    defparam i14075_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14076_3_lut (.I0(\data_in_frame[7] [3]), .I1(rx_data[3]), .I2(n35586), 
            .I3(GND_net), .O(n22479));   // verilog/coms.v(127[12] 300[6])
    defparam i14076_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14077_3_lut (.I0(\data_in_frame[7] [2]), .I1(rx_data[2]), .I2(n35586), 
            .I3(GND_net), .O(n22480));   // verilog/coms.v(127[12] 300[6])
    defparam i14077_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14078_3_lut (.I0(\data_in_frame[7] [1]), .I1(rx_data[1]), .I2(n35586), 
            .I3(GND_net), .O(n22481));   // verilog/coms.v(127[12] 300[6])
    defparam i14078_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut (.I0(control_mode[0]), .I1(control_mode[6]), 
            .I2(n10_adj_4859), .I3(control_mode[2]), .O(n20608));   // verilog/TinyFPGA_B.v(165[5:22])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14079_3_lut (.I0(\data_in_frame[7] [0]), .I1(rx_data[0]), .I2(n35586), 
            .I3(GND_net), .O(n22482));   // verilog/coms.v(127[12] 300[6])
    defparam i14079_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14080_3_lut (.I0(\data_in_frame[6] [7]), .I1(rx_data[7]), .I2(n35579), 
            .I3(GND_net), .O(n22483));   // verilog/coms.v(127[12] 300[6])
    defparam i14080_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14081_3_lut (.I0(\data_in_frame[6] [6]), .I1(rx_data[6]), .I2(n35579), 
            .I3(GND_net), .O(n22484));   // verilog/coms.v(127[12] 300[6])
    defparam i14081_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14082_3_lut (.I0(\data_in_frame[6] [5]), .I1(rx_data[5]), .I2(n35579), 
            .I3(GND_net), .O(n22485));   // verilog/coms.v(127[12] 300[6])
    defparam i14082_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i3_4_lut_4_lut (.I0(r_SM_Main_adj_5088[1]), .I1(r_SM_Main_adj_5088[0]), 
            .I2(r_SM_Main_adj_5088[2]), .I3(r_SM_Main_2__N_3454[1]), .O(n41168));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i14083_3_lut (.I0(\data_in_frame[6] [4]), .I1(rx_data[4]), .I2(n35579), 
            .I3(GND_net), .O(n22486));   // verilog/coms.v(127[12] 300[6])
    defparam i14083_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14084_3_lut (.I0(\data_in_frame[6] [3]), .I1(rx_data[3]), .I2(n35579), 
            .I3(GND_net), .O(n22487));   // verilog/coms.v(127[12] 300[6])
    defparam i14084_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14085_3_lut (.I0(\data_in_frame[6] [2]), .I1(rx_data[2]), .I2(n35579), 
            .I3(GND_net), .O(n22488));   // verilog/coms.v(127[12] 300[6])
    defparam i14085_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14086_3_lut (.I0(\data_in_frame[6] [1]), .I1(rx_data[1]), .I2(n35579), 
            .I3(GND_net), .O(n22489));   // verilog/coms.v(127[12] 300[6])
    defparam i14086_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14087_3_lut (.I0(\data_in_frame[6] [0]), .I1(rx_data[0]), .I2(n35579), 
            .I3(GND_net), .O(n22490));   // verilog/coms.v(127[12] 300[6])
    defparam i14087_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14088_3_lut (.I0(\data_in_frame[5] [7]), .I1(rx_data[7]), .I2(n35585), 
            .I3(GND_net), .O(n22491));   // verilog/coms.v(127[12] 300[6])
    defparam i14088_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14089_3_lut (.I0(\data_in_frame[5] [6]), .I1(rx_data[6]), .I2(n35585), 
            .I3(GND_net), .O(n22492));   // verilog/coms.v(127[12] 300[6])
    defparam i14089_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14090_3_lut (.I0(\data_in_frame[5] [5]), .I1(rx_data[5]), .I2(n35585), 
            .I3(GND_net), .O(n22493));   // verilog/coms.v(127[12] 300[6])
    defparam i14090_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14091_3_lut (.I0(\data_in_frame[5] [4]), .I1(rx_data[4]), .I2(n35585), 
            .I3(GND_net), .O(n22494));   // verilog/coms.v(127[12] 300[6])
    defparam i14091_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14092_3_lut (.I0(\data_in_frame[5] [3]), .I1(rx_data[3]), .I2(n35585), 
            .I3(GND_net), .O(n22495));   // verilog/coms.v(127[12] 300[6])
    defparam i14092_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14093_3_lut (.I0(\data_in_frame[5] [2]), .I1(rx_data[2]), .I2(n35585), 
            .I3(GND_net), .O(n22496));   // verilog/coms.v(127[12] 300[6])
    defparam i14093_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14094_3_lut (.I0(\data_in_frame[5] [1]), .I1(rx_data[1]), .I2(n35585), 
            .I3(GND_net), .O(n22497));   // verilog/coms.v(127[12] 300[6])
    defparam i14094_3_lut.LUT_INIT = 16'hacac;
    EEPROM eeprom (.GND_net(GND_net), .CLK_c(CLK_c), .n3460({n3461}), 
           .\state[1] (state_adj_5082[1]), .\state[1]_adj_12 (state_adj_5111[1]), 
           .\state[2] (state_adj_5111[2]), .n7(n7_adj_5015), .read(read), 
           .\state[0] (state_adj_5082[0]), .n15(n15_adj_4901), .\state[3] (state_adj_5111[3]), 
           .n6(n6_adj_5025), .n35272(n35272), .n36440(n36440), .n35591(n35591), 
           .n27098(n27098), .n35254(n35254), .VCC_net(VCC_net), .n22318(n22318), 
           .rw(rw), .n35362(n35362), .data_ready(data_ready), .n4760(n4760), 
           .\saved_addr[0] (saved_addr[0]), .\state[0]_adj_13 (state_adj_5111[0]), 
           .n3957(n3957), .n27086(n27086), .n4(n4_adj_4945), .n4_adj_14(n4_adj_4877), 
           .n10(n10_adj_4908), .n10_adj_15(n10_adj_4902), .\state_7__N_3881[3] (state_7__N_3881[3]), 
           .n10_adj_16(n10_adj_5010), .scl_enable_N_3958(scl_enable_N_3958), 
           .scl_enable(scl_enable), .sda_enable(sda_enable), .\state_7__N_3865[0] (state_7__N_3865[0]), 
           .n5180(n5180), .n15_adj_17(n15_adj_4922), .n8(n8_adj_4879), 
           .n987({scl}), .n20731(n20731), .n20726(n20726), .n39285(n39285), 
           .n22330(n22330), .\data[0] (data[0]), .n22321(n22321), .n22300(n22300), 
           .\data[1] (data[1]), .n22299(n22299), .\data[2] (data[2]), 
           .n22298(n22298), .\data[3] (data[3]), .n22297(n22297), .\data[4] (data[4]), 
           .n22296(n22296), .\data[5] (data[5]), .n22295(n22295), .\data[6] (data[6]), 
           .n22294(n22294), .\data[7] (data[7])) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(249[10] 259[6])
    SB_LUT4 i14095_3_lut (.I0(\data_in_frame[5] [0]), .I1(rx_data[0]), .I2(n35585), 
            .I3(GND_net), .O(n22498));   // verilog/coms.v(127[12] 300[6])
    defparam i14095_3_lut.LUT_INIT = 16'hacac;
    coms neopxl_color_23__I_0 (.GND_net(GND_net), .n22423(n22423), .\data_in_frame[14] ({\data_in_frame[14] }), 
         .clk32MHz(clk32MHz), .n22422(n22422), .\data_in_frame[10] ({\data_in_frame[10] }), 
         .n22421(n22421), .\data_in_frame[5] ({\data_in_frame[5] }), .n22420(n22420), 
         .n22419(n22419), .n22418(n22418), .\data_in_frame[15] ({\data_in_frame[15] }), 
         .n22417(n22417), .n22416(n22416), .n22415(n22415), .n22414(n22414), 
         .n36883(n36883), .\data_in_frame[1] ({\data_in_frame[1] }), .n22413(n22413), 
         .ID({ID}), .\data_in_frame[11] ({\data_in_frame[11] }), .\data_in_frame[12] ({\data_in_frame[12] }), 
         .\data_in_frame[8] ({\data_in_frame[8] }), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .\data_in_frame[9] ({\data_in_frame[9] }), .rx_data({rx_data}), 
         .n22412(n22412), .\data_in_frame[2] ({\data_in_frame[2] }), .rx_data_ready(rx_data_ready), 
         .\data_in_frame[21] ({\data_in_frame[21] }), .n22411(n22411), .setpoint({setpoint}), 
         .\data_in_frame[7] ({\data_in_frame[7] }), .\data_in_frame[3] ({\data_in_frame[3] }), 
         .\data_in_frame[6] ({\data_in_frame[6] }), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .\data_out_frame[25] ({\data_out_frame[25] }), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .\data_out_frame[23] ({\data_out_frame[23] }), .\data_out_frame[24] ({\data_out_frame[24] }), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .\data_out_frame[20] ({\data_out_frame[20] }), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .n18082(n18082), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .\data_out_frame[12] ({\data_out_frame[12] }), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .\data_out_frame[9] ({\data_out_frame[9] }), .\data_out_frame[11] ({\data_out_frame[11] }), 
         .\data_out_frame[10] ({\data_out_frame[10] }), .\data_out_frame[4] ({\data_out_frame[4] }), 
         .\data_out_frame[6] ({\data_out_frame[6] }), .\data_in[2] ({\data_in[2] }), 
         .\data_in[1] ({\data_in[1] }), .\data_in[3] ({\data_in[3] }), .\data_in[0] ({\data_in[0] }), 
         .tx_active(tx_active), .n35579(n35579), .n35562(n35562), .\state[0] (state_adj_5111[0]), 
         .\state[1] (state_adj_5111[1]), .\state[2] (state_adj_5111[2]), 
         .\state[3] (state_adj_5111[3]), .n15(n15_adj_4901), .n35561(n35561), 
         .n35586(n35586), .n10(n10_adj_4902), .n22370(n22370), .n22369(n22369), 
         .n22368(n22368), .n22367(n22367), .n22366(n22366), .n22365(n22365), 
         .n22364(n22364), .n22363(n22363), .n22362(n22362), .control_mode({control_mode}), 
         .n22361(n22361), .n22360(n22360), .n22359(n22359), .n22358(n22358), 
         .n22357(n22357), .n22356(n22356), .n22355(n22355), .PWMLimit({PWMLimit}), 
         .n22354(n22354), .n22353(n22353), .n22352(n22352), .n22351(n22351), 
         .n22350(n22350), .n22349(n22349), .n22348(n22348), .n22347(n22347), 
         .n22346(n22346), .n22345(n22345), .DE_c(DE_c), .n22344(n22344), 
         .n22343(n22343), .n22342(n22342), .n22341(n22341), .n22340(n22340), 
         .LED_c(LED_c), .n35575(n35575), .n35585(n35585), .n35568(n35568), 
         .n22840(n22840), .IntegralLimit({IntegralLimit}), .n22839(n22839), 
         .n22838(n22838), .n22837(n22837), .n22836(n22836), .n22835(n22835), 
         .n22834(n22834), .n22833(n22833), .n22832(n22832), .n22831(n22831), 
         .n22830(n22830), .n22829(n22829), .n22828(n22828), .n22827(n22827), 
         .n22826(n22826), .n22825(n22825), .n22824(n22824), .n22823(n22823), 
         .n22822(n22822), .n22821(n22821), .n22820(n22820), .n22819(n22819), 
         .n22818(n22818), .n22783(n22783), .n22782(n22782), .n22781(n22781), 
         .n22780(n22780), .n22779(n22779), .n22778(n22778), .n22777(n22777), 
         .n22776(n22776), .n22775(n22775), .n22774(n22774), .n22773(n22773), 
         .n22772(n22772), .n22771(n22771), .n22770(n22770), .n22769(n22769), 
         .n22768(n22768), .n22767(n22767), .n22766(n22766), .n22765(n22765), 
         .n22764(n22764), .n22763(n22763), .n22762(n22762), .n22761(n22761), 
         .n22760(n22760), .n22759(n22759), .n22758(n22758), .n22757(n22757), 
         .n22756(n22756), .n22755(n22755), .n22754(n22754), .n22753(n22753), 
         .n22752(n22752), .\Kp[1] (Kp[1]), .n22751(n22751), .\Kp[2] (Kp[2]), 
         .n22750(n22750), .\Kp[3] (Kp[3]), .n22749(n22749), .\Kp[4] (Kp[4]), 
         .n22748(n22748), .\Kp[5] (Kp[5]), .n22747(n22747), .\Kp[6] (Kp[6]), 
         .n22746(n22746), .\Kp[7] (Kp[7]), .n22745(n22745), .\Kp[8] (Kp[8]), 
         .n22744(n22744), .\Kp[9] (Kp[9]), .n22743(n22743), .\Kp[10] (Kp[10]), 
         .n22742(n22742), .\Kp[11] (Kp[11]), .n22741(n22741), .\Kp[12] (Kp[12]), 
         .n22740(n22740), .\Kp[13] (Kp[13]), .n22739(n22739), .\Kp[14] (Kp[14]), 
         .n22738(n22738), .\Kp[15] (Kp[15]), .n22737(n22737), .\Ki[1] (Ki[1]), 
         .n22736(n22736), .\Ki[2] (Ki[2]), .n22735(n22735), .\Ki[3] (Ki[3]), 
         .n22734(n22734), .\Ki[4] (Ki[4]), .n22733(n22733), .\Ki[5] (Ki[5]), 
         .n22732(n22732), .\Ki[6] (Ki[6]), .n22731(n22731), .\Ki[7] (Ki[7]), 
         .n22730(n22730), .\Ki[8] (Ki[8]), .n22729(n22729), .\Ki[9] (Ki[9]), 
         .n22728(n22728), .\Ki[10] (Ki[10]), .n22727(n22727), .\Ki[11] (Ki[11]), 
         .n22726(n22726), .\Ki[12] (Ki[12]), .n22725(n22725), .\Ki[13] (Ki[13]), 
         .n22724(n22724), .\Ki[14] (Ki[14]), .n22721(n22721), .\Ki[15] (Ki[15]), 
         .n22720(n22720), .n22719(n22719), .n22718(n22718), .n22717(n22717), 
         .n22716(n22716), .n22715(n22715), .n22714(n22714), .n22713(n22713), 
         .n22712(n22712), .n22711(n22711), .n22710(n22710), .n22709(n22709), 
         .n22708(n22708), .n22707(n22707), .n22706(n22706), .n22705(n22705), 
         .n22704(n22704), .n22703(n22703), .n22702(n22702), .n22701(n22701), 
         .n22700(n22700), .n22699(n22699), .n22698(n22698), .n22697(n22697), 
         .n22696(n22696), .n22695(n22695), .n22694(n22694), .n22693(n22693), 
         .n22692(n22692), .n22691(n22691), .n22690(n22690), .n22689(n22689), 
         .n22688(n22688), .n22687(n22687), .n22686(n22686), .n22685(n22685), 
         .n22684(n22684), .n22683(n22683), .n22682(n22682), .n22681(n22681), 
         .n22680(n22680), .n22679(n22679), .n22678(n22678), .n22677(n22677), 
         .n22676(n22676), .n22675(n22675), .n22674(n22674), .n22673(n22673), 
         .n22672(n22672), .n22671(n22671), .n22670(n22670), .n22669(n22669), 
         .n22668(n22668), .n22667(n22667), .n22666(n22666), .n22665(n22665), 
         .n22664(n22664), .n22663(n22663), .n22662(n22662), .n22661(n22661), 
         .n22660(n22660), .n22659(n22659), .n22658(n22658), .n22657(n22657), 
         .n22656(n22656), .n21865(n21865), .n22339(n22339), .n22338(n22338), 
         .n22337(n22337), .n22336(n22336), .n22335(n22335), .n22334(n22334), 
         .n22333(n22333), .n22315(n22315), .n22314(n22314), .n22312(n22312), 
         .neopxl_color({neopxl_color}), .n22311(n22311), .\Ki[0] (Ki[0]), 
         .n22310(n22310), .\Kp[0] (Kp[0]), .n22309(n22309), .n22655(n22655), 
         .n22654(n22654), .n22653(n22653), .n22652(n22652), .n22651(n22651), 
         .n22650(n22650), .n22649(n22649), .n22648(n22648), .n22647(n22647), 
         .n22646(n22646), .n22645(n22645), .n22644(n22644), .n22643(n22643), 
         .n22642(n22642), .n22641(n22641), .n22640(n22640), .n22639(n22639), 
         .n22638(n22638), .n22637(n22637), .n22636(n22636), .n22635(n22635), 
         .n22634(n22634), .n22633(n22633), .n22632(n22632), .n22631(n22631), 
         .n22630(n22630), .n22629(n22629), .n22628(n22628), .n22627(n22627), 
         .n22626(n22626), .n22625(n22625), .n22624(n22624), .n22623(n22623), 
         .n22622(n22622), .n22621(n22621), .n22620(n22620), .n22619(n22619), 
         .n22618(n22618), .n22617(n22617), .n22616(n22616), .n22615(n22615), 
         .n22614(n22614), .n22613(n22613), .n22612(n22612), .n22611(n22611), 
         .n22610(n22610), .n22609(n22609), .n22608(n22608), .n22607(n22607), 
         .n22606(n22606), .n22605(n22605), .n22604(n22604), .n22603(n22603), 
         .n22602(n22602), .n22601(n22601), .n22600(n22600), .n22599(n22599), 
         .n22598(n22598), .n22597(n22597), .n22596(n22596), .n22595(n22595), 
         .n22594(n22594), .n22593(n22593), .n22592(n22592), .n22591(n22591), 
         .n22590(n22590), .n22589(n22589), .n22588(n22588), .n22587(n22587), 
         .n22586(n22586), .n22585(n22585), .n22584(n22584), .n22583(n22583), 
         .n22582(n22582), .n22581(n22581), .n22580(n22580), .n22579(n22579), 
         .n22578(n22578), .n22577(n22577), .n22576(n22576), .n22575(n22575), 
         .n22574(n22574), .n22573(n22573), .n22572(n22572), .n22571(n22571), 
         .n22570(n22570), .n22569(n22569), .n22568(n22568), .n22567(n22567), 
         .n22566(n22566), .n22565(n22565), .n22564(n22564), .n22563(n22563), 
         .n22292(n22292), .n22562(n22562), .n3957(n3957), .n15_adj_3(n15_adj_4922), 
         .scl_enable_N_3958(scl_enable_N_3958), .n22561(n22561), .n22560(n22560), 
         .n22559(n22559), .n22558(n22558), .n22557(n22557), .n22556(n22556), 
         .n22555(n22555), .n22554(n22554), .n22553(n22553), .n22552(n22552), 
         .n22551(n22551), .n22550(n22550), .n22549(n22549), .n22548(n22548), 
         .n22547(n22547), .n22546(n22546), .n22545(n22545), .n22544(n22544), 
         .n22543(n22543), .n22542(n22542), .n22541(n22541), .n22540(n22540), 
         .n22539(n22539), .n22538(n22538), .n22498(n22498), .n22497(n22497), 
         .n22496(n22496), .n22495(n22495), .n22494(n22494), .n22493(n22493), 
         .n22492(n22492), .n22491(n22491), .n22490(n22490), .n22489(n22489), 
         .n22488(n22488), .n22487(n22487), .n22486(n22486), .n22485(n22485), 
         .n22484(n22484), .n22483(n22483), .n22482(n22482), .n22481(n22481), 
         .n22480(n22480), .n22479(n22479), .n22478(n22478), .n22477(n22477), 
         .n22476(n22476), .n22475(n22475), .n5180(n5180), .n22434(n22434), 
         .n22433(n22433), .n22432(n22432), .n22431(n22431), .n22430(n22430), 
         .n22429(n22429), .n22428(n22428), .n22427(n22427), .n22426(n22426), 
         .n22425(n22425), .n22424(n22424), .n21920(n21920), .n22195(n22195), 
         .r_SM_Main({r_SM_Main_adj_5088}), .\r_SM_Main_2__N_3454[1] (r_SM_Main_2__N_3454[1]), 
         .tx_o(tx_o), .n13920(n13920), .VCC_net(VCC_net), .\r_Bit_Index[0] (r_Bit_Index_adj_5090[0]), 
         .n4(n4_adj_4868), .n22817(n22817), .n22319(n22319), .n41168(n41168), 
         .tx_enable(tx_enable), .n22012(n22012), .n22193(n22193), .n26980(n26980), 
         .n4_adj_4(n4_adj_4921), .n4_adj_5(n4_adj_4920), .\r_Bit_Index[0]_adj_6 (r_Bit_Index[0]), 
         .n20781(n20781), .r_Rx_Data(r_Rx_Data), .RX_N_10(RX_N_10), .n20776(n20776), 
         .n4_adj_7(n4_adj_4914), .n22843(n22843), .n22847(n22847), .n22308(n22308), 
         .n22307(n22307), .n22306(n22306), .n22305(n22305), .n22304(n22304), 
         .n22303(n22303), .n22302(n22302)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(137[8] 160[4])
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.encoder1_position({encoder1_position}), 
            .GND_net(GND_net), .clk32MHz(clk32MHz), .data_o({quadA_debounced_adj_4905, 
            quadB_debounced_adj_4906}), .n37217(n37217), .reg_B({reg_B_adj_5099}), 
            .VCC_net(VCC_net), .ENCODER1_A_c_1(ENCODER1_A_c_1), .ENCODER1_B_c_0(ENCODER1_B_c_0), 
            .n22849(n22849), .n22320(n22320)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(193[15] 198[4])
    pwm PWM (.n39932(n39932), .VCC_net(VCC_net), .INHA_c(INHA_c), .clk32MHz(clk32MHz), 
        .n20604(n20604), .GND_net(GND_net), .n20602(n20602), .\pwm_counter[6] (pwm_counter[6]), 
        .\pwm_counter[8] (pwm_counter[8]), .\pwm_counter[7] (pwm_counter[7]), 
        .\pwm_counter[13] (pwm_counter[13]), .\pwm_counter[10] (pwm_counter[10]), 
        .\pwm_counter[9] (pwm_counter[9]), .\pwm_counter[17] (pwm_counter[17]), 
        .\pwm_counter[22] (pwm_counter[22]), .\pwm_counter[14] (pwm_counter[14]), 
        .\pwm_counter[18] (pwm_counter[18]), .\pwm_counter[21] (pwm_counter[21]), 
        .\pwm_counter[16] (pwm_counter[16]), .\pwm_counter[12] (pwm_counter[12]), 
        .\pwm_counter[15] (pwm_counter[15]), .\pwm_counter[19] (pwm_counter[19]), 
        .\pwm_counter[11] (pwm_counter[11]), .\pwm_counter[20] (pwm_counter[20]), 
        .\pwm_counter[31] (pwm_counter[31]), .\pwm_counter[0] (pwm_counter[0]), 
        .\pwm_counter[5] (pwm_counter[5]), .\pwm_counter[4] (pwm_counter[4]), 
        .\pwm_counter[3] (pwm_counter[3]), .\pwm_counter[2] (pwm_counter[2]), 
        .\pwm_counter[1] (pwm_counter[1])) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(89[6] 94[3])
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (encoder0_position, GND_net, clk32MHz, 
            data_o, n38219, reg_B, VCC_net, ENCODER0_B_c_0, n22848, 
            n22316, ENCODER0_A_c_1) /* synthesis syn_module_defined=1 */ ;
    output [23:0]encoder0_position;
    input GND_net;
    input clk32MHz;
    output [1:0]data_o;
    output n38219;
    output [1:0]reg_B;
    input VCC_net;
    input ENCODER0_B_c_0;
    input n22848;
    input n22316;
    input ENCODER0_A_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n30838, n3038, n30839;
    wire [23:0]n3042;
    
    wire n30837, n30836, n30835, n30834, count_enable, B_delayed, 
        A_delayed, n30833, n30832, n30831, n30830, n30829, n30828, 
        n30827, n30826, n30825, n30824, n30823, n30822, n30821, 
        n30820, n30819, n30818, count_direction, n30817, n30840;
    
    SB_CARRY add_713_23 (.CI(n30838), .I0(encoder0_position[21]), .I1(n3038), 
            .CO(n30839));
    SB_LUT4 add_713_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n3038), 
            .I3(n30837), .O(n3042[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_22 (.CI(n30837), .I0(encoder0_position[20]), .I1(n3038), 
            .CO(n30838));
    SB_LUT4 add_713_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n3038), 
            .I3(n30836), .O(n3042[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_21 (.CI(n30836), .I0(encoder0_position[19]), .I1(n3038), 
            .CO(n30837));
    SB_LUT4 add_713_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n3038), 
            .I3(n30835), .O(n3042[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_20 (.CI(n30835), .I0(encoder0_position[18]), .I1(n3038), 
            .CO(n30836));
    SB_LUT4 add_713_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n3038), 
            .I3(n30834), .O(n3042[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_19 (.CI(n30834), .I0(encoder0_position[17]), .I1(n3038), 
            .CO(n30835));
    SB_DFFE count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[0]));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 add_713_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n3038), 
            .I3(n30833), .O(n3042[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_18 (.CI(n30833), .I0(encoder0_position[16]), .I1(n3038), 
            .CO(n30834));
    SB_LUT4 add_713_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n3038), 
            .I3(n30832), .O(n3042[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_17 (.CI(n30832), .I0(encoder0_position[15]), .I1(n3038), 
            .CO(n30833));
    SB_LUT4 add_713_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n3038), 
            .I3(n30831), .O(n3042[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_16 (.CI(n30831), .I0(encoder0_position[14]), .I1(n3038), 
            .CO(n30832));
    SB_LUT4 add_713_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n3038), 
            .I3(n30830), .O(n3042[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_15 (.CI(n30830), .I0(encoder0_position[13]), .I1(n3038), 
            .CO(n30831));
    SB_LUT4 add_713_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n3038), 
            .I3(n30829), .O(n3042[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_14 (.CI(n30829), .I0(encoder0_position[12]), .I1(n3038), 
            .CO(n30830));
    SB_LUT4 add_713_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n3038), 
            .I3(n30828), .O(n3042[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_13 (.CI(n30828), .I0(encoder0_position[11]), .I1(n3038), 
            .CO(n30829));
    SB_LUT4 add_713_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n3038), 
            .I3(n30827), .O(n3042[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_12 (.CI(n30827), .I0(encoder0_position[10]), .I1(n3038), 
            .CO(n30828));
    SB_LUT4 add_713_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n3038), 
            .I3(n30826), .O(n3042[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_11 (.CI(n30826), .I0(encoder0_position[9]), .I1(n3038), 
            .CO(n30827));
    SB_LUT4 add_713_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n3038), 
            .I3(n30825), .O(n3042[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_10 (.CI(n30825), .I0(encoder0_position[8]), .I1(n3038), 
            .CO(n30826));
    SB_LUT4 add_713_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n3038), 
            .I3(n30824), .O(n3042[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_9 (.CI(n30824), .I0(encoder0_position[7]), .I1(n3038), 
            .CO(n30825));
    SB_LUT4 add_713_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n3038), 
            .I3(n30823), .O(n3042[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_8 (.CI(n30823), .I0(encoder0_position[6]), .I1(n3038), 
            .CO(n30824));
    SB_LUT4 add_713_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n3038), 
            .I3(n30822), .O(n3042[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFE count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[23]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[22]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[21]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[20]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[19]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[18]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[17]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[16]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[15]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[14]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[13]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[12]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[11]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[10]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[9]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[8]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[7]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[6]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[5]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[4]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[3]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[2]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .E(count_enable), 
            .D(n3042[1]));   // quad.v(35[10] 41[6])
    SB_CARRY add_713_7 (.CI(n30822), .I0(encoder0_position[5]), .I1(n3038), 
            .CO(n30823));
    SB_LUT4 add_713_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n3038), 
            .I3(n30821), .O(n3042[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_6 (.CI(n30821), .I0(encoder0_position[4]), .I1(n3038), 
            .CO(n30822));
    SB_LUT4 add_713_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n3038), 
            .I3(n30820), .O(n3042[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_5 (.CI(n30820), .I0(encoder0_position[3]), .I1(n3038), 
            .CO(n30821));
    SB_LUT4 add_713_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n3038), 
            .I3(n30819), .O(n3042[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_4 (.CI(n30819), .I0(encoder0_position[2]), .I1(n3038), 
            .CO(n30820));
    SB_LUT4 add_713_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n3038), 
            .I3(n30818), .O(n3042[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_3 (.CI(n30818), .I0(encoder0_position[1]), .I1(n3038), 
            .CO(n30819));
    SB_LUT4 add_713_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n30817), .O(n3042[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_2 (.CI(n30817), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n30818));
    SB_CARRY add_713_1 (.CI(GND_net), .I0(n3038), .I1(n3038), .CO(n30817));
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1133_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n3038));   // quad.v(37[5] 40[8])
    defparam i1133_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_713_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n3038), 
            .I3(n30840), .O(n3042[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_713_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n3038), 
            .I3(n30839), .O(n3042[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_713_24 (.CI(n30839), .I0(encoder0_position[22]), .I1(n3038), 
            .CO(n30840));
    SB_LUT4 add_713_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n3038), 
            .I3(n30838), .O(n3042[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_713_23_lut.LUT_INIT = 16'hC33C;
    \grp_debouncer(2,100)_U0  debounce (.n38219(n38219), .reg_B({reg_B}), 
            .GND_net(GND_net), .clk32MHz(clk32MHz), .VCC_net(VCC_net), 
            .ENCODER0_B_c_0(ENCODER0_B_c_0), .n22848(n22848), .data_o({data_o}), 
            .n22316(n22316), .ENCODER0_A_c_1(ENCODER0_A_c_1));   // quad.v(15[37] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,100)_U0 
//

module \grp_debouncer(2,100)_U0  (n38219, reg_B, GND_net, clk32MHz, 
            VCC_net, ENCODER0_B_c_0, n22848, data_o, n22316, ENCODER0_A_c_1);
    output n38219;
    output [1:0]reg_B;
    input GND_net;
    input clk32MHz;
    input VCC_net;
    input ENCODER0_B_c_0;
    input n22848;
    output [1:0]data_o;
    input n22316;
    input ENCODER0_A_c_1;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [6:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n12;
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_6__N_3697;
    wire [6:0]n33;
    
    wire n31688, n31687, n31686, n31685, n31684, n31683;
    
    SB_LUT4 i5_4_lut (.I0(cnt_reg[1]), .I1(cnt_reg[4]), .I2(cnt_reg[3]), 
            .I3(cnt_reg[6]), .O(n12));
    defparam i5_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut (.I0(cnt_reg[5]), .I1(n12), .I2(cnt_reg[0]), .I3(cnt_reg[2]), 
            .O(n38219));
    defparam i6_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n38219), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_6__N_3697));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 cnt_reg_1514_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n31688), .O(n33[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1514_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_1514_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n31687), .O(n33[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1514_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1514_add_4_7 (.CI(n31687), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n31688));
    SB_LUT4 cnt_reg_1514_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n31686), .O(n33[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1514_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1514_add_4_6 (.CI(n31686), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n31687));
    SB_LUT4 cnt_reg_1514_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n31685), .O(n33[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1514_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1514_add_4_5 (.CI(n31685), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n31686));
    SB_LUT4 cnt_reg_1514_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n31684), .O(n33[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1514_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1514_add_4_4 (.CI(n31684), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n31685));
    SB_LUT4 cnt_reg_1514_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n31683), .O(n33[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1514_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_CARRY cnt_reg_1514_add_4_3 (.CI(n31683), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n31684));
    SB_LUT4 cnt_reg_1514_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n33[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1514_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1514_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n31683));
    SB_DFFSR cnt_reg_1514__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n33[0]), 
            .R(cnt_next_6__N_3697));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(ENCODER0_B_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n22848));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n22316));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1514__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n33[1]), 
            .R(cnt_next_6__N_3697));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1514__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n33[2]), 
            .R(cnt_next_6__N_3697));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1514__i3 (.Q(cnt_reg[3]), .C(clk32MHz), .D(n33[3]), 
            .R(cnt_next_6__N_3697));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1514__i4 (.Q(cnt_reg[4]), .C(clk32MHz), .D(n33[4]), 
            .R(cnt_next_6__N_3697));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1514__i5 (.Q(cnt_reg[5]), .C(clk32MHz), .D(n33[5]), 
            .R(cnt_next_6__N_3697));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1514__i6 (.Q(cnt_reg[6]), .C(clk32MHz), .D(n33[6]), 
            .R(cnt_next_6__N_3697));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(ENCODER0_A_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    
endmodule
//
// Verilog Description of module neopixel
//

module neopixel (GND_net, VCC_net, clk32MHz, \neo_pixel_transmitter.done , 
            \neo_pixel_transmitter.t0 , start, \state[1] , LED_c, \state_3__N_369[1] , 
            n14, n36364, n21969, timer, n37680, neopxl_color, n22814, 
            n22813, n22812, n22811, n22810, n22809, n22808, n22807, 
            n22806, n22805, n22804, n22803, n22802, n22801, n22800, 
            n22799, n22798, n22797, n22796, n22795, n22794, n22793, 
            n22792, n22791, n22790, n22789, n22788, n22787, n22786, 
            n22785, n22784, n22326, \neo_pixel_transmitter.done_N_583 , 
            NEOPXL_c, n34460, n22291, n39196) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input VCC_net;
    input clk32MHz;
    output \neo_pixel_transmitter.done ;
    output [31:0]\neo_pixel_transmitter.t0 ;
    output start;
    output \state[1] ;
    input LED_c;
    output \state_3__N_369[1] ;
    output n14;
    output n36364;
    output n21969;
    output [31:0]timer;
    output n37680;
    input [23:0]neopxl_color;
    input n22814;
    input n22813;
    input n22812;
    input n22811;
    input n22810;
    input n22809;
    input n22808;
    input n22807;
    input n22806;
    input n22805;
    input n22804;
    input n22803;
    input n22802;
    input n22801;
    input n22800;
    input n22799;
    input n22798;
    input n22797;
    input n22796;
    input n22795;
    input n22794;
    input n22793;
    input n22792;
    input n22791;
    input n22790;
    input n22789;
    input n22788;
    input n22787;
    input n22786;
    input n22785;
    input n22784;
    input n22326;
    input \neo_pixel_transmitter.done_N_583 ;
    output NEOPXL_c;
    input n34460;
    input n22291;
    output n39196;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [31:0]n971;
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    wire [31:0]n255;
    
    wire n21935, n22215, n30970, \neo_pixel_transmitter.done_N_577 , 
        n40929;
    wire [31:0]n1;
    
    wire n2819, n40624, n31588, n3001, n3017, n31589, n2302, n2292, 
        n22, n2299, n2309, n30, n2294, n2306, n2297, n34, n2301, 
        n2307, n2291, n2305, n32, n2298, n2295, n2304, n2300, 
        n33, n2308, n2296, n2303, n2293, n31, n2324, n2225, 
        n40637, n21, n23, n22_adj_4705, n24, n36, n2193, n2194, 
        n2206, n2204, n28, n2203, n2209, n32_adj_4706, n2208, 
        n2201, n2192, n2196, n30_adj_4707, n2195, n2207, n2205, 
        n2199, n31_adj_4708, n2202, n2197, n2198, n2200, n29, 
        n2126, n40636, n2918, n40625, n30650, n2093, n2103, n2097, 
        n26, n2104, n2096, n2094, n2098, n29_adj_4709, n2099, 
        n2109, n20, n2101, n2105, n2095, n2108, n28_adj_4710, 
        n2102, n2100, n32_adj_4711, n2106, n2107, n19, n2693, 
        n2704, n28_adj_4712, n2699, n2706, n2694, n2691, n38, 
        n2709, n27886, n2701, n2696, n2697, n36_adj_4713, n2700, 
        n2705, n42, n2702, n2690, n2689, n2708, n40, n2687, 
        n2703, n2695, n41, n2688, n2698, n2692, n2707, n39, 
        n2720, n2798, n2804, n2791, n2795, n40_adj_4714, n2796, 
        n2793, n2788, n2808, n38_adj_4715, n2789, n2800, n2803, 
        n2805, n39_adj_4716, n2792, n2787, n2801, n2799, n37, 
        n2786, n2797, n34_adj_4717, n1037, n40622, n2794, n2806, 
        n2807, n2790, n42_adj_4718, n46, n2621, n40619, n2802, 
        n2809, n33_adj_4719, n2, n1007, n40623, n1006, n3102, 
        n3090, n3103, n3085, n42_adj_4720, n3089, n3094, n3101, 
        n3098, n46_adj_4721, n3099, n3091, n3106, n3100, n44, 
        n3097, n3088, n3104, n3092, n45, n3105, n3083, n3093, 
        n3096, n43, n3108, n3109, n40_adj_4722, n3107, n3087, 
        n3086, n48, n52, n3095, n3084, n39_adj_4723, n3116, n3002, 
        n31587, n906, n1005, n608, n708, n8234, n7764, n36524, 
        n19304, n807, n36370, n9244, n838, n36488, n905, n38308, 
        n22070, n19296, n1009, n1008, n38343, n6_adj_4724, n4, 
        n40618, n25, n27, n26_adj_4725, n28_adj_4726, n37_adj_4727, 
        n20592, n36428, n32422, n36426;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    
    wire n39580, n28022, n36512, n39581, n36536, n1334, n40635, 
        n2588, n31792, n2589, n31791, n3003, n31586, n2590, n31790, 
        n29_adj_4729, n30_adj_4730, n20697, n3004, n31585, n32530;
    wire [31:0]one_wire_N_520;
    
    wire n2591, n31789, n3005, n31584, n2592, n31788, n14_adj_4731, 
        n9_adj_4732, n1158, n28010, n3006, n31583, n2593, n31787, 
        n3007, n31582, n1308, n1304, n1305, n14_adj_4733, n1302, 
        n1307, n12_adj_4734, n3008, n31581, n2594, n31786, n1303, 
        n1309, n16, n1301, n1306, n2027, n40633, n3209, n27896, 
        n35, n11_adj_4735, n29_adj_4736, n51, n48_adj_4737, n37_adj_4738, 
        n23_adj_4739, n53, n39_adj_4740, n46_adj_4741, n27_adj_4742, 
        n57, n63, n43_adj_4743, n47, n25_adj_4744, n33_adj_4745, 
        n47_adj_4746, n61, n45_adj_4747, n59, n17, n15_adj_4748, 
        n55, n44_adj_4749, n31_adj_4750, n41_adj_4751, n49, n43_adj_4752, 
        n54, n45_adj_4753, n13_adj_4754, n19_adj_4755, n21_adj_4756, 
        n49_adj_4757, n32566, n1172, n39203, n20719, n36326, n41597;
    wire [4:0]color_bit_N_563;
    
    wire n40723, n40729, n39243, n40657;
    wire [3:0]state_3__N_369;
    
    wire n3009, n31580, n2595, n31785, n30658, n40621, n1103, 
        n30778, n2596, n31784, n1104, n30777, n31579, n31578, 
        n2597, n31783, n31577, n31576, n30651, n30659, n31575, 
        n2598, n31782, n2599, n31781, n4983, n1105, n30776, n2600, 
        n31780, n2601, n31779, n1235, n40634, n2602, n31778, n31574, 
        n1205, n1206, n1204, n1207, n14_adj_4760, n31573, n2603, 
        n31777, n31572, n1203, n1209, n9_adj_4761, n2604, n31776, 
        n2605, n31775, n31571, n1202, n1208, n1106, n30775, n2606, 
        n31774, n2607, n31773, n1107, n30774, n2608, n31772, n31570, 
        n2609, n31771, n1108, n30773, n31569, n1109, n31568, n31567, 
        n31770, n31566, n31769, n31565, n31768, n31564, n31563, 
        n31767, n31562, n31766, n31561, n31765, n31560, n31559, 
        n31764, n31558, n31557, n27850, n31556, n31763, n31555, 
        n31554, n31762, n31761, n31553, n30876, n30875, n30657, 
        n30874, n31760, n31759, n31758, n30873, n31757, n30649, 
        n31756, n31755, n31754, n39270, n30678, n31753, n30677, 
        n31752, n31751, n31750, n31749, n31748, n30872, n2885, 
        n31747, n2886, n31746, n2887, n31745, n2888, n31744, n30676, 
        n2889, n31743, n2890, n31742, n2891, n31741, n2892, n31740;
    wire [31:0]n133;
    
    wire n36470, n27516, n38147, n36538, n2893, n31739, n30656, 
        n2894, n31738, n2895, n31737, n30675, n2896, n31736, n30871, 
        n36_adj_4764, n25_adj_4765, n34_adj_4766, n40_adj_4767, n38_adj_4768, 
        n2897, n31735, n30870, n30655, n30869, n39_adj_4769, n37_adj_4770, 
        n30674, n2898, n31734, n31636, n30673, n30648, n31635, 
        n30868, n2899, n31733, n2900, n31732, n31634, n31633, 
        n2901, n31731, n30672, n30654, n31632, n2902, n31730, 
        n30671, n31631, n30867, n31630, n2903, n31729, n2904, 
        n31728, n30670, n31629, n2905, n31727, n31628, n31627, 
        n30866, n31626, n31625, n2906, n31726, n31624, n30865, 
        n30864, n31623, n2907, n31725, n2908, n31724, n30863, 
        n2909, n31622, n30862, n40840, n38446, n40834, n38449, 
        n40822, n38455, n2989, n2990, n40_adj_4772, n2984, n2988, 
        n2986, n44_adj_4773, n2994, n42_adj_4774, n2999, n3000, 
        n2992, n2997, n43_adj_4775, n30861, n30860, n30669, n2996, 
        n2985, n2995, n2987, n41_adj_4777, n2993, n38_adj_4778, 
        n2998, n2991, n46_adj_4779, n50, n37_adj_4780, n2003, n2008, 
        n18_adj_4782, n1996, n1998, n2006, n2007, n28_adj_4783, 
        n1997, n1999, n2005, n2000, n26_adj_4784, n1994, n2001, 
        n2004, n1995, n27_adj_4785, n2002, n2009, n25_adj_4786, 
        n1928, n40632, n1895, n1902, n1899, n1897, n26_adj_4787, 
        n30859, n1907, n1909, n19_adj_4789, n1908, n1900, n16_adj_4790, 
        n30858, n1904, n1901, n1906, n1898, n24_adj_4792, n1905, 
        n1903, n28_adj_4793, n1896, n1829, n40631, n31723, n30857, 
        n31621, n31722, n30856, n31721, n31720, n31719, n31620, 
        n31619, n31718, n31618, n31617, n1806, n1803, n1798, n1805, 
        n24_adj_4796, n1808, n1804, n1802, n1807, n22_adj_4797, 
        n1800, n1799, n1797, n1801, n23_adj_4798, n1796, n1809, 
        n21_adj_4799, n31717, n1730, n40630, n31616, n30855, n31716, 
        n31615, n1499, n1400, n1433, n32019, n1500, n1401, n32018, 
        n30854, n1501, n1402, n32017, n1502, n1403, n32016, n1503, 
        n1404, n32015, n1504, n1405, n32014, n1505, n1406, n32013, 
        n31614, n1506, n1407, n32012, n1507, n1408, n32011, n1508, 
        n1409, n40626, n32010, n1704, n1709, n16_adj_4803, n1509, 
        n30853, n1136, n32009, n32008, n32007, n31715, n31613, 
        n32006, n1707, n1697, n1702, n1699, n22_adj_4805, n1706, 
        n1701, n1708, n20_adj_4806, n1703, n1698, n24_adj_4807, 
        n1705, n1700, n1631, n40629, n1608, n1606, n1604, n1603, 
        n20_adj_4809, n1602, n1609, n13_adj_4810, n1598, n1600, 
        n18_adj_4811, n1605, n1599, n22_adj_4812, n1601, n1607, 
        n1532, n40628, n31714, n31612, n30653, n30668, n30852, 
        n30667, n30851, n32005, n32004, n40627, n32003, n31611, 
        n30652, n31992, n31713, n31991, n30850, n31990, n30666, 
        n31989, n31988, n31987, n31986, n31985, n31984, n31983, 
        n31982, n31981, n31980, n30849, n31979, n31978, n31977, 
        n31976, n31975, n31974, n31973, n31972, n31971, n31970, 
        n31969, n31968, n31967, n31966, n31965, n31964, n30848, 
        n31963, n31610, n31962, n31961, n31960, n31959, n31958, 
        n31957, n30665, n31956, n31955, n31954, n31953, n31952, 
        n31951, n31950, n31949, n31948, n31947, n31946, n31945, 
        n31944, n31943, n31942, n31941, n31940, n31939, n31938, 
        n31937, n31936, n31935, n31934, n31933, n31932, n31931, 
        n31930, n35558, n18_adj_4816, n20_adj_4817, n15_adj_4818, 
        n31929, n31928, n31927, n31926, n31925, n31924, n31923, 
        n31922, n31921, n31920, n31919, n31918, n30847, n111, 
        n40726, n31712, n31609, n30846, n4_adj_4819, n31608, n31711, 
        n31607, n31606, n31917, n31710, n31142, n31141, n31140, 
        n31139, n31709, n31138, n31137, n31136, n31135, n31916, 
        n116, n31708, n31915, n31707, n31605, n31604, n30664, 
        n30663, n38337, n40720, n31914, n31913, n31912, n20_adj_4820, 
        n31706, n31603, n31602, n31097, n31096, n31705, n31095, 
        n31094, n31601, n31093, n31092, n31091, n31090, n31089, 
        n36830, n31704, n31600, n27860, n12_adj_4821, n31911, n31910, 
        n31703, n31599, n31909, n31598, n31702, n31908, n31907, 
        n31597, n31701, n31596, n31906, n31700, n30662, n31699, 
        n27902, n16_adj_4822, n31905, n31595, n17_adj_4823, n30661, 
        n30660, n30974, n31904, n31903, n31902, n31901, n31900, 
        n31594, n31899, n31898, n31897, n31896, n31895, n31593, 
        n31592, n31894, n31893, n31892, n31891, n31890, n31889, 
        n31888, n31887, n31886, n31885, n31884, n31883, n31882, 
        n31881, n31880, n31879, n31878, n31877, n2390, n31876, 
        n2391, n31875, n2392, n31874, n2393, n31873, n2394, n31872, 
        n2395, n31871, n2396, n31870, n2397, n31869, n2398, n31868, 
        n2399, n31867, n2400, n31866, n2401, n31865, n2402, n31864, 
        n2403, n31863, n2404, n31862, n2405, n31861, n2406, n31860, 
        n2407, n31859, n2408, n40638, n31858, n2409, n2489, n2423, 
        n31857, n2490, n31856, n2491, n31855, n2492, n31854, n2493, 
        n31853, n2494, n31852, n2495, n31851, n2496, n31850, n2497, 
        n31849, n2498, n31848, n2499, n31847, n2500, n31846, n2501, 
        n31845, n2502, n31844, n2503, n31843, n2504, n31842, n2505, 
        n31841, n2506, n31840, n2507, n31839, n2508, n40639, n31838, 
        n2509, n2522, n31837, n31836, n31835, n31834, n31833, 
        n31832, n31831, n31830, n30973, n31829, n31828, n31827, 
        n31826, n31591, n31825, n31824, n31823, n31822, n31821, 
        n31820, n31819, n30972, n31818, n40640, n31817, n31590, 
        n30971, n7_adj_4824, n40702, n39869, n30_adj_4825, n48_adj_4826, 
        n46_adj_4827, n24_adj_4828, n34_adj_4829, n22_adj_4830, n47_adj_4831, 
        n38_adj_4832, n36_adj_4833, n37_adj_4834, n35_adj_4835, n45_adj_4836, 
        n44_adj_4837, n40_adj_4838, n27_adj_4839, n38_adj_4840, n43_adj_4841, 
        n42_adj_4842, n41_adj_4843, n43_adj_4844, n45_adj_4845, n47_adj_4846, 
        n54_adj_4847, n49_adj_4848, n40654, n27_adj_4849, n33_adj_4850, 
        n32_adj_4851, n31_adj_4852, n35_adj_4853, n37_adj_4854;
    
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(clk32MHz), .E(n21935), 
            .D(n255[19]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n30970));
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk32MHz), .E(n40929), .D(\neo_pixel_transmitter.done_N_577 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30597_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40624));
    defparam i30597_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2076_11 (.CI(n31588), .I0(n3001), .I1(n3017), .CO(n31589));
    SB_DFFESR bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(clk32MHz), .E(n21935), 
            .D(n255[18]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_2_lut (.I0(n2302), .I1(n2292), .I2(GND_net), .I3(GND_net), 
            .O(n22));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i11_4_lut (.I0(bit_ctr[12]), .I1(n22), .I2(n2299), .I3(n2309), 
            .O(n30));
    defparam i11_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 i15_4_lut (.I0(n2294), .I1(n30), .I2(n2306), .I3(n2297), 
            .O(n34));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(n2301), .I1(n2307), .I2(n2291), .I3(n2305), 
            .O(n32));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n2298), .I1(n2295), .I2(n2304), .I3(n2300), 
            .O(n33));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n2308), .I1(n2296), .I2(n2303), .I3(n2293), 
            .O(n31));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(n31), .I1(n33), .I2(n32), .I3(n34), .O(n2324));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30610_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40637));
    defparam i30610_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(clk32MHz), .E(n21935), 
            .D(n255[17]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(clk32MHz), .E(n21935), 
            .D(n255[16]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(clk32MHz), .E(n21935), 
            .D(n255[15]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(clk32MHz), .E(n21935), 
            .D(n255[14]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(clk32MHz), .E(n21935), 
            .D(n255[13]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(clk32MHz), .E(n21935), 
            .D(n255[12]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(clk32MHz), .E(n21935), 
            .D(n255[11]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(clk32MHz), .E(n21935), 
            .D(n255[10]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(clk32MHz), .E(n21935), 
            .D(n255[9]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(clk32MHz), .E(n21935), 
            .D(n255[8]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(clk32MHz), .E(n21935), 
            .D(n255[7]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(clk32MHz), .E(n21935), 
            .D(n255[6]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(clk32MHz), .E(n21935), 
            .D(n255[5]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(clk32MHz), .E(n21935), 
            .D(n255[4]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(clk32MHz), .E(n21935), 
            .D(n255[3]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(clk32MHz), .E(n21935), 
            .D(n255[2]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(clk32MHz), .E(n21935), 
            .D(n255[1]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i16_4_lut (.I0(n21), .I1(n23), .I2(n22_adj_4705), .I3(n24), 
            .O(n36));   // verilog/neopixel.v(104[14:39])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(n2193), .I1(n2194), .I2(n2206), .I3(n2204), 
            .O(n28));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1527 (.I0(n2203), .I1(n28), .I2(bit_ctr[13]), 
            .I3(n2209), .O(n32_adj_4706));
    defparam i14_4_lut_adj_1527.LUT_INIT = 16'hfeee;
    SB_LUT4 i12_4_lut_adj_1528 (.I0(n2208), .I1(n2201), .I2(n2192), .I3(n2196), 
            .O(n30_adj_4707));
    defparam i12_4_lut_adj_1528.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1529 (.I0(n2195), .I1(n2207), .I2(n2205), .I3(n2199), 
            .O(n31_adj_4708));
    defparam i13_4_lut_adj_1529.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1530 (.I0(n2202), .I1(n2197), .I2(n2198), .I3(n2200), 
            .O(n29));
    defparam i11_4_lut_adj_1530.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n29), .I1(n31_adj_4708), .I2(n30_adj_4707), 
            .I3(n32_adj_4706), .O(n2225));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30609_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40636));
    defparam i30609_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30598_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40625));
    defparam i30598_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_5_lut (.I0(GND_net), .I1(bit_ctr[3]), .I2(GND_net), 
            .I3(n30650), .O(n255[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9_3_lut (.I0(n2093), .I1(n2103), .I2(n2097), .I3(GND_net), 
            .O(n26));
    defparam i9_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12_4_lut_adj_1531 (.I0(n2104), .I1(n2096), .I2(n2094), .I3(n2098), 
            .O(n29_adj_4709));
    defparam i12_4_lut_adj_1531.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut (.I0(bit_ctr[14]), .I1(n2099), .I2(n2109), .I3(GND_net), 
            .O(n20));
    defparam i3_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i11_4_lut_adj_1532 (.I0(n2101), .I1(n2105), .I2(n2095), .I3(n2108), 
            .O(n28_adj_4710));
    defparam i11_4_lut_adj_1532.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1533 (.I0(n29_adj_4709), .I1(n2102), .I2(n26), 
            .I3(n2100), .O(n32_adj_4711));
    defparam i15_4_lut_adj_1533.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(n2106), .I1(n2107), .I2(GND_net), .I3(GND_net), 
            .O(n19));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i16_4_lut_adj_1534 (.I0(n19), .I1(n32_adj_4711), .I2(n28_adj_4710), 
            .I3(n20), .O(n2126));
    defparam i16_4_lut_adj_1534.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut (.I0(n2693), .I1(n2704), .I2(GND_net), .I3(GND_net), 
            .O(n28_adj_4712));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1535 (.I0(n2699), .I1(n2706), .I2(n2694), .I3(n2691), 
            .O(n38));
    defparam i15_4_lut_adj_1535.LUT_INIT = 16'hfffe;
    SB_LUT4 i19480_2_lut (.I0(bit_ctr[8]), .I1(n2709), .I2(GND_net), .I3(GND_net), 
            .O(n27886));
    defparam i19480_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1536 (.I0(n2701), .I1(n2696), .I2(n2697), .I3(n27886), 
            .O(n36_adj_4713));
    defparam i13_4_lut_adj_1536.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n2700), .I1(n38), .I2(n28_adj_4712), .I3(n2705), 
            .O(n42));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1537 (.I0(n2702), .I1(n2690), .I2(n2689), .I3(n2708), 
            .O(n40));
    defparam i17_4_lut_adj_1537.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1538 (.I0(n2687), .I1(n36_adj_4713), .I2(n2703), 
            .I3(n2695), .O(n41));
    defparam i18_4_lut_adj_1538.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1539 (.I0(n2688), .I1(n2698), .I2(n2692), .I3(n2707), 
            .O(n39));
    defparam i16_4_lut_adj_1539.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n39), .I1(n41), .I2(n40), .I3(n42), .O(n2720));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1540 (.I0(n2798), .I1(n2804), .I2(n2791), .I3(n2795), 
            .O(n40_adj_4714));
    defparam i16_4_lut_adj_1540.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1541 (.I0(n2796), .I1(n2793), .I2(n2788), .I3(n2808), 
            .O(n38_adj_4715));
    defparam i14_4_lut_adj_1541.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1542 (.I0(n2789), .I1(n2800), .I2(n2803), .I3(n2805), 
            .O(n39_adj_4716));
    defparam i15_4_lut_adj_1542.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1543 (.I0(n2792), .I1(n2787), .I2(n2801), .I3(n2799), 
            .O(n37));
    defparam i13_4_lut_adj_1543.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_2_lut (.I0(n2786), .I1(n2797), .I2(GND_net), .I3(GND_net), 
            .O(n34_adj_4717));
    defparam i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i30595_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40622));
    defparam i30595_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i18_4_lut_adj_1544 (.I0(n2794), .I1(n2806), .I2(n2807), .I3(n2790), 
            .O(n42_adj_4718));
    defparam i18_4_lut_adj_1544.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1545 (.I0(n37), .I1(n39_adj_4716), .I2(n38_adj_4715), 
            .I3(n40_adj_4714), .O(n46));
    defparam i22_4_lut_adj_1545.LUT_INIT = 16'hfffe;
    SB_LUT4 i30592_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40619));
    defparam i30592_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i9_3_lut_adj_1546 (.I0(bit_ctr[7]), .I1(n2802), .I2(n2809), 
            .I3(GND_net), .O(n33_adj_4719));
    defparam i9_3_lut_adj_1546.LUT_INIT = 16'hecec;
    SB_LUT4 i30156_2_lut (.I0(n2), .I1(n971[28]), .I2(GND_net), .I3(GND_net), 
            .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i30156_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i23_4_lut (.I0(n33_adj_4719), .I1(n46), .I2(n42_adj_4718), 
            .I3(n34_adj_4717), .O(n2819));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30596_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40623));
    defparam i30596_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30154_2_lut (.I0(n2), .I1(n971[29]), .I2(GND_net), .I3(GND_net), 
            .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam i30154_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i15_4_lut_adj_1547 (.I0(n3102), .I1(n3090), .I2(n3103), .I3(n3085), 
            .O(n42_adj_4720));
    defparam i15_4_lut_adj_1547.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1548 (.I0(n3089), .I1(n3094), .I2(n3101), .I3(n3098), 
            .O(n46_adj_4721));
    defparam i19_4_lut_adj_1548.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1549 (.I0(n3099), .I1(n3091), .I2(n3106), .I3(n3100), 
            .O(n44));
    defparam i17_4_lut_adj_1549.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1550 (.I0(n3097), .I1(n3088), .I2(n3104), .I3(n3092), 
            .O(n45));
    defparam i18_4_lut_adj_1550.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1551 (.I0(n3105), .I1(n3083), .I2(n3093), .I3(n3096), 
            .O(n43));
    defparam i16_4_lut_adj_1551.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(bit_ctr[4]), .I1(n3108), .I2(n3109), .I3(GND_net), 
            .O(n40_adj_4722));
    defparam i13_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i21_4_lut (.I0(n3107), .I1(n42_adj_4720), .I2(n3087), .I3(n3086), 
            .O(n48));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n43), .I1(n45), .I2(n44), .I3(n46_adj_4721), 
            .O(n52));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut (.I0(n3095), .I1(n3084), .I2(GND_net), .I3(GND_net), 
            .O(n39_adj_4723));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i26_4_lut (.I0(n39_adj_4723), .I1(n52), .I2(n48), .I3(n40_adj_4722), 
            .O(n3116));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n31587), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_i672_3_lut (.I0(n906), .I1(n971[30]), .I2(n2), .I3(GND_net), 
            .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19387_2_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(GND_net), .O(n608));   // verilog/neopixel.v(22[26:36])
    defparam i19387_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_4_lut (.I0(n708), .I1(n8234), .I2(n7764), .I3(n608), 
            .O(n36524));
    defparam i2_4_lut.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_2_lut (.I0(bit_ctr[28]), .I1(n36524), .I2(GND_net), .I3(GND_net), 
            .O(n19304));
    defparam i1_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i28254_3_lut (.I0(n36524), .I1(n708), .I2(n7764), .I3(GND_net), 
            .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam i28254_3_lut.LUT_INIT = 16'h8282;
    SB_LUT4 mod_5_i606_3_lut (.I0(n36370), .I1(n9244), .I2(n838), .I3(GND_net), 
            .O(n36488));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i606_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 i28281_3_lut (.I0(n906), .I1(n905), .I2(n36488), .I3(GND_net), 
            .O(n38308));
    defparam i28281_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(n22070), .I1(n38308), .I2(bit_ctr[26]), .I3(n19296), 
            .O(n2));   // verilog/neopixel.v(22[26:36])
    defparam i4_4_lut.LUT_INIT = 16'h0111;
    SB_LUT4 i1_2_lut_adj_1552 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n19296));
    defparam i1_2_lut_adj_1552.LUT_INIT = 16'h9999;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n2), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i675_3_lut (.I0(n19296), .I1(n971[27]), .I2(n2), .I3(GND_net), 
            .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i28315_3_lut (.I0(n971[28]), .I1(n971[31]), .I2(n971[29]), 
            .I3(GND_net), .O(n38343));
    defparam i28315_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), .I3(GND_net), 
            .O(n6_adj_4724));
    defparam i2_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i3_4_lut (.I0(n2), .I1(n6_adj_4724), .I2(n1005), .I3(n38343), 
            .O(n1037));
    defparam i3_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i30207_2_lut (.I0(n2), .I1(n971[31]), .I2(GND_net), .I3(GND_net), 
            .O(n4));   // verilog/neopixel.v(22[26:36])
    defparam i30207_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i30591_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40618));
    defparam i30591_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17_4_lut_adj_1553 (.I0(n25), .I1(n27), .I2(n26_adj_4725), 
            .I3(n28_adj_4726), .O(n37_adj_4727));   // verilog/neopixel.v(104[14:39])
    defparam i17_4_lut_adj_1553.LUT_INIT = 16'hfffe;
    SB_LUT4 i26414_2_lut (.I0(start), .I1(n20592), .I2(GND_net), .I3(GND_net), 
            .O(n36428));
    defparam i26414_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i29743_4_lut (.I0(n32422), .I1(n36426), .I2(\neo_pixel_transmitter.done ), 
            .I3(state[0]), .O(n39580));
    defparam i29743_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i53_4_lut (.I0(n36428), .I1(n28022), .I2(\state[1] ), .I3(n36426), 
            .O(n36512));
    defparam i53_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i52_4_lut (.I0(n36512), .I1(n39581), .I2(state[0]), .I3(\neo_pixel_transmitter.done ), 
            .O(n36536));
    defparam i52_4_lut.LUT_INIT = 16'h3335;
    SB_LUT4 i30608_1_lut (.I0(n1334), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40635));
    defparam i30608_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2076_10 (.CI(n31587), .I0(n3002), .I1(n3017), .CO(n31588));
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n31792), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(clk32MHz), .E(n21935), 
            .D(n255[22]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n31791), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(clk32MHz), .E(n21935), 
            .D(n255[29]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1808_23 (.CI(n31791), .I0(n2589), .I1(n2621), .CO(n31792));
    SB_DFFESR bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(clk32MHz), .E(n21935), 
            .D(n255[28]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n31586), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n31790), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i19_4_lut_adj_1554 (.I0(n37_adj_4727), .I1(n29_adj_4729), .I2(n36), 
            .I3(n30_adj_4730), .O(n20697));   // verilog/neopixel.v(104[14:39])
    defparam i19_4_lut_adj_1554.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(clk32MHz), .E(n21935), 
            .D(n255[21]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_2076_9 (.CI(n31586), .I0(n3003), .I1(n3017), .CO(n31587));
    SB_CARRY mod_5_add_1808_22 (.CI(n31790), .I0(n2590), .I1(n2621), .CO(n31791));
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n31585), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_8 (.CI(n31585), .I0(n3004), .I1(n3017), .CO(n31586));
    SB_LUT4 i1_3_lut (.I0(n32530), .I1(one_wire_N_520[4]), .I2(one_wire_N_520[3]), 
            .I3(GND_net), .O(n36426));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n31789), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n31584), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_21 (.CI(n31789), .I0(n2591), .I1(n2621), .CO(n31790));
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n31788), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6_4_lut (.I0(one_wire_N_520[5]), .I1(one_wire_N_520[11]), .I2(one_wire_N_520[7]), 
            .I3(n20697), .O(n14_adj_4731));   // verilog/neopixel.v(104[14:39])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(n9_adj_4732), .I1(n14_adj_4731), .I2(one_wire_N_520[10]), 
            .I3(one_wire_N_520[8]), .O(n20592));   // verilog/neopixel.v(104[14:39])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i261_2_lut (.I0(LED_c), .I1(\state_3__N_369[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n1158));   // verilog/neopixel.v(40[18] 45[12])
    defparam i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_adj_1555 (.I0(n20592), .I1(n36426), .I2(GND_net), 
            .I3(GND_net), .O(n28010));
    defparam i2_2_lut_adj_1555.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_1808_20 (.CI(n31788), .I0(n2592), .I1(n2621), .CO(n31789));
    SB_CARRY mod_5_add_2076_7 (.CI(n31584), .I0(n3005), .I1(n3017), .CO(n31585));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n31583), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n31787), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_6 (.CI(n31583), .I0(n3006), .I1(n3017), .CO(n31584));
    SB_CARRY mod_5_add_1808_19 (.CI(n31787), .I0(n2593), .I1(n2621), .CO(n31788));
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n31582), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_5 (.CI(n31582), .I0(n3007), .I1(n3017), .CO(n31583));
    SB_DFFESR bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(clk32MHz), .E(n21935), 
            .D(n255[20]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i5_3_lut (.I0(n1308), .I1(n1304), .I2(n1305), .I3(GND_net), 
            .O(n14_adj_4733));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_2_lut_adj_1556 (.I0(n1302), .I1(n1307), .I2(GND_net), .I3(GND_net), 
            .O(n12_adj_4734));
    defparam i3_2_lut_adj_1556.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n31581), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_4 (.CI(n31581), .I0(n3008), .I1(n3017), .CO(n31582));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n31786), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7_4_lut_adj_1557 (.I0(bit_ctr[22]), .I1(n14_adj_4733), .I2(n1303), 
            .I3(n1309), .O(n16));
    defparam i7_4_lut_adj_1557.LUT_INIT = 16'hfefc;
    SB_LUT4 i8_4_lut (.I0(n1301), .I1(n16), .I2(n12_adj_4734), .I3(n1306), 
            .O(n1334));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30606_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40633));
    defparam i30606_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19614_4_lut (.I0(one_wire_N_520[9]), .I1(n20697), .I2(one_wire_N_520[11]), 
            .I3(one_wire_N_520[10]), .O(n28022));
    defparam i19614_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i19490_2_lut (.I0(bit_ctr[3]), .I1(n3209), .I2(GND_net), .I3(GND_net), 
            .O(n27896));
    defparam i19490_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20_4_lut (.I0(n35), .I1(n11_adj_4735), .I2(n29_adj_4736), 
            .I3(n51), .O(n48_adj_4737));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1558 (.I0(n37_adj_4738), .I1(n23_adj_4739), .I2(n53), 
            .I3(n39_adj_4740), .O(n46_adj_4741));
    defparam i18_4_lut_adj_1558.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1559 (.I0(n27_adj_4742), .I1(n57), .I2(n63), 
            .I3(n43_adj_4743), .O(n47));
    defparam i19_4_lut_adj_1559.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1560 (.I0(n25_adj_4744), .I1(n33_adj_4745), .I2(n47_adj_4746), 
            .I3(n61), .O(n45_adj_4747));
    defparam i17_4_lut_adj_1560.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1561 (.I0(n59), .I1(n17), .I2(n15_adj_4748), 
            .I3(n55), .O(n44_adj_4749));
    defparam i16_4_lut_adj_1561.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1562 (.I0(n31_adj_4750), .I1(n41_adj_4751), .I2(n49), 
            .I3(n27896), .O(n43_adj_4752));
    defparam i15_4_lut_adj_1562.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1563 (.I0(n45_adj_4747), .I1(n47), .I2(n46_adj_4741), 
            .I3(n48_adj_4737), .O(n54));
    defparam i26_4_lut_adj_1563.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1564 (.I0(n45_adj_4753), .I1(n13_adj_4754), .I2(n19_adj_4755), 
            .I3(n21_adj_4756), .O(n49_adj_4757));
    defparam i21_4_lut_adj_1564.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n49_adj_4757), .I1(n54), .I2(n43_adj_4752), 
            .I3(n44_adj_4749), .O(n32566));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i275_2_lut (.I0(n28022), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n1172));   // verilog/neopixel.v(103[9] 111[12])
    defparam i275_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i15_4_lut_adj_1565 (.I0(n14), .I1(n39203), .I2(\state[1] ), 
            .I3(n20719), .O(n36364));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15_4_lut_adj_1565.LUT_INIT = 16'h303a;
    SB_LUT4 i1_4_lut (.I0(state[0]), .I1(n36326), .I2(n1172), .I3(\state[1] ), 
            .O(n21969));
    defparam i1_4_lut.LUT_INIT = 16'hafcc;
    SB_LUT4 i1_rep_319_2_lut (.I0(bit_ctr[3]), .I1(n32566), .I2(GND_net), 
            .I3(GND_net), .O(n41597));
    defparam i1_rep_319_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29633_3_lut (.I0(n3209), .I1(bit_ctr[3]), .I2(n32566), .I3(GND_net), 
            .O(color_bit_N_563[4]));
    defparam i29633_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i29739_4_lut (.I0(n40723), .I1(n41597), .I2(n40729), .I3(bit_ctr[2]), 
            .O(n39243));
    defparam i29739_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i18673_4_lut (.I0(n40657), .I1(\state_3__N_369[1] ), .I2(n39243), 
            .I3(color_bit_N_563[4]), .O(state_3__N_369[0]));   // verilog/neopixel.v(40[18] 45[12])
    defparam i18673_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY mod_5_add_1808_18 (.CI(n31786), .I0(n2594), .I1(n2621), .CO(n31787));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n3009), .I1(n3009), .I2(n40618), 
            .I3(n31580), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n31785), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_17 (.CI(n31785), .I0(n2595), .I1(n2621), .CO(n31786));
    SB_LUT4 add_21_13_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(n30658), .O(n255[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_3 (.CI(n31580), .I0(n3009), .I1(n40618), .CO(n31581));
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i30594_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40621));
    defparam i30594_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_736_8_lut (.I0(n4), .I1(n4), .I2(n1037), .I3(n30778), 
            .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n31784), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n40618), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_736_7_lut (.I0(n1005), .I1(n1005), .I2(n1037), .I3(n30777), 
            .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_16 (.CI(n31784), .I0(n2596), .I1(n2621), .CO(n31785));
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n40618), 
            .CO(n31580));
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n31579), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n31578), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n31783), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_28 (.CI(n31578), .I0(n3084), .I1(n3116), .CO(n31579));
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n31577), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_27 (.CI(n31577), .I0(n3085), .I1(n3116), .CO(n31578));
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n31576), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_5 (.CI(n30650), .I0(bit_ctr[3]), .I1(GND_net), .CO(n30651));
    SB_CARRY add_21_13 (.CI(n30658), .I0(bit_ctr[11]), .I1(GND_net), .CO(n30659));
    SB_CARRY mod_5_add_2143_26 (.CI(n31576), .I0(n3086), .I1(n3116), .CO(n31577));
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n31575), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_15 (.CI(n31783), .I0(n2597), .I1(n2621), .CO(n31784));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n31782), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_25 (.CI(n31575), .I0(n3087), .I1(n3116), .CO(n31576));
    SB_CARRY mod_5_add_1808_14 (.CI(n31782), .I0(n2598), .I1(n2621), .CO(n31783));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n31781), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_7 (.CI(n30777), .I0(n1005), .I1(n1037), .CO(n30778));
    SB_LUT4 i3322_4_lut (.I0(n28010), .I1(n1158), .I2(\state[1] ), .I3(n20719), 
            .O(n4983));
    defparam i3322_4_lut.LUT_INIT = 16'h3f35;
    SB_LUT4 mod_5_add_736_6_lut (.I0(n1006), .I1(n1006), .I2(n1037), .I3(n30776), 
            .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_13 (.CI(n31781), .I0(n2599), .I1(n2621), .CO(n31782));
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n31780), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_12 (.CI(n31780), .I0(n2600), .I1(n2621), .CO(n31781));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n31779), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_11 (.CI(n31779), .I0(n2601), .I1(n2621), .CO(n31780));
    SB_LUT4 i30607_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40634));
    defparam i30607_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n31778), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_10 (.CI(n31778), .I0(n2602), .I1(n2621), .CO(n31779));
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n31574), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i6_4_lut_adj_1566 (.I0(n1205), .I1(n1206), .I2(n1204), .I3(n1207), 
            .O(n14_adj_4760));
    defparam i6_4_lut_adj_1566.LUT_INIT = 16'hfffe;
    SB_DFFESR bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(clk32MHz), .E(n21935), 
            .D(n255[0]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_2143_24 (.CI(n31574), .I0(n3088), .I1(n3116), .CO(n31575));
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n31573), .O(n51)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_6 (.CI(n30776), .I0(n1006), .I1(n1037), .CO(n30777));
    SB_CARRY mod_5_add_2143_23 (.CI(n31573), .I0(n3089), .I1(n3116), .CO(n31574));
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n31777), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n31572), .O(n49)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_22 (.CI(n31572), .I0(n3090), .I1(n3116), .CO(n31573));
    SB_LUT4 i1_3_lut_adj_1567 (.I0(bit_ctr[23]), .I1(n1203), .I2(n1209), 
            .I3(GND_net), .O(n9_adj_4761));
    defparam i1_3_lut_adj_1567.LUT_INIT = 16'hecec;
    SB_CARRY mod_5_add_1808_9 (.CI(n31777), .I0(n2603), .I1(n2621), .CO(n31778));
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n31776), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_8 (.CI(n31776), .I0(n2604), .I1(n2621), .CO(n31777));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n31775), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n31571), .O(n47_adj_4746)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7_4_lut_adj_1568 (.I0(n9_adj_4761), .I1(n14_adj_4760), .I2(n1202), 
            .I3(n1208), .O(n1235));
    defparam i7_4_lut_adj_1568.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_736_5_lut (.I0(n1007), .I1(n1007), .I2(n1037), .I3(n30775), 
            .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_7 (.CI(n31775), .I0(n2605), .I1(n2621), .CO(n31776));
    SB_CARRY mod_5_add_736_5 (.CI(n30775), .I0(n1007), .I1(n1037), .CO(n30776));
    SB_CARRY mod_5_add_2143_21 (.CI(n31571), .I0(n3091), .I1(n3116), .CO(n31572));
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n31774), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_6 (.CI(n31774), .I0(n2606), .I1(n2621), .CO(n31775));
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n31773), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_5 (.CI(n31773), .I0(n2607), .I1(n2621), .CO(n31774));
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n30774), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n31772), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n31570), .O(n45_adj_4753)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_4 (.CI(n31772), .I0(n2608), .I1(n2621), .CO(n31773));
    SB_CARRY mod_5_add_2143_20 (.CI(n31570), .I0(n3092), .I1(n3116), .CO(n31571));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n40619), 
            .I3(n31771), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_3 (.CI(n31771), .I0(n2609), .I1(n40619), .CO(n31772));
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n40619), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_4 (.CI(n30774), .I0(n1008), .I1(n1037), .CO(n30775));
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n40622), 
            .I3(n30773), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n31569), .O(n43_adj_4743)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_3 (.CI(n30773), .I0(n1009), .I1(n40622), .CO(n30774));
    SB_CARRY mod_5_add_2143_19 (.CI(n31569), .I0(n3093), .I1(n3116), .CO(n31570));
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n40622), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n31568), .O(n41_adj_4751)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_18 (.CI(n31568), .I0(n3094), .I1(n3116), .CO(n31569));
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n40622), 
            .CO(n30773));
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n31567), .O(n39_adj_4740)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n40619), 
            .CO(n31771));
    SB_CARRY mod_5_add_2143_17 (.CI(n31567), .I0(n3095), .I1(n3116), .CO(n31568));
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n31770), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n31566), .O(n37_adj_4738)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_16 (.CI(n31566), .I0(n3096), .I1(n3116), .CO(n31567));
    SB_LUT4 mod_5_add_1875_24_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n31769), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_24 (.CI(n31769), .I0(n2688), .I1(n2720), .CO(n31770));
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n31565), .O(n35)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_23_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n31768), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_15 (.CI(n31565), .I0(n3097), .I1(n3116), .CO(n31566));
    SB_CARRY mod_5_add_1875_23 (.CI(n31768), .I0(n2689), .I1(n2720), .CO(n31769));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n31564), .O(n33_adj_4745)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_14 (.CI(n31564), .I0(n3098), .I1(n3116), .CO(n31565));
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n31563), .O(n31_adj_4750)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_13 (.CI(n31563), .I0(n3099), .I1(n3116), .CO(n31564));
    SB_LUT4 mod_5_add_1875_22_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n31767), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n31562), .O(n29_adj_4736)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_12 (.CI(n31562), .I0(n3100), .I1(n3116), .CO(n31563));
    SB_CARRY mod_5_add_1875_22 (.CI(n31767), .I0(n2690), .I1(n2720), .CO(n31768));
    SB_LUT4 mod_5_add_1875_21_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n31766), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_21 (.CI(n31766), .I0(n2691), .I1(n2720), .CO(n31767));
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n31561), .O(n27_adj_4742)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_11 (.CI(n31561), .I0(n3101), .I1(n3116), .CO(n31562));
    SB_LUT4 mod_5_add_1875_20_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n31765), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n31560), .O(n25_adj_4744)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_10 (.CI(n31560), .I0(n3102), .I1(n3116), .CO(n31561));
    SB_LUT4 i3_4_lut_4_lut (.I0(n36370), .I1(n19304), .I2(n807), .I3(bit_ctr[27]), 
            .O(n838));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n31559), .O(n23_adj_4739)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_9 (.CI(n31559), .I0(n3103), .I1(n3116), .CO(n31560));
    SB_CARRY mod_5_add_1875_20 (.CI(n31765), .I0(n2692), .I1(n2720), .CO(n31766));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n31764), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n31558), .O(n21_adj_4756)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_8 (.CI(n31558), .I0(n3104), .I1(n3116), .CO(n31559));
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n31557), .O(n19_adj_4755)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3814_2_lut_3_lut (.I0(bit_ctr[29]), .I1(n27850), .I2(bit_ctr[28]), 
            .I3(GND_net), .O(n7764));
    defparam i3814_2_lut_3_lut.LUT_INIT = 16'h6060;
    SB_CARRY mod_5_add_2143_7 (.CI(n31557), .I0(n3105), .I1(n3116), .CO(n31558));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n31556), .O(n17)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_19 (.CI(n31764), .I0(n2693), .I1(n2720), .CO(n31765));
    SB_LUT4 mod_5_add_1875_18_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n31763), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_6 (.CI(n31556), .I0(n3106), .I1(n3116), .CO(n31557));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n31555), .O(n15_adj_4748)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_5 (.CI(n31555), .I0(n3107), .I1(n3116), .CO(n31556));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n31554), .O(n13_adj_4754)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i29405_3_lut_4_lut (.I0(bit_ctr[29]), .I1(n27850), .I2(n36524), 
            .I3(bit_ctr[28]), .O(n36370));
    defparam i29405_3_lut_4_lut.LUT_INIT = 16'h9666;
    SB_CARRY mod_5_add_2143_4 (.CI(n31554), .I0(n3108), .I1(n3116), .CO(n31555));
    SB_CARRY mod_5_add_1875_18 (.CI(n31763), .I0(n2694), .I1(n2720), .CO(n31764));
    SB_LUT4 mod_5_add_1875_17_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n31762), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_17 (.CI(n31762), .I0(n2695), .I1(n2720), .CO(n31763));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n31761), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n40621), 
            .I3(n31553), .O(n11_adj_4735)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_add_2_33_lut (.I0(one_wire_N_520[16]), .I1(timer[31]), 
            .I2(n1[31]), .I3(n30876), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2143_3 (.CI(n31553), .I0(n3109), .I1(n40621), .CO(n31554));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n40621), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_16 (.CI(n31761), .I0(n2696), .I1(n2720), .CO(n31762));
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n40621), 
            .CO(n31553));
    SB_LUT4 sub_14_add_2_32_lut (.I0(one_wire_N_520[24]), .I1(timer[30]), 
            .I2(n1[30]), .I3(n30875), .O(n22_adj_4705)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_32 (.CI(n30875), .I0(timer[30]), .I1(n1[30]), 
            .CO(n30876));
    SB_LUT4 add_21_12_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(n30657), .O(n255[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_31_lut (.I0(one_wire_N_520[22]), .I1(timer[29]), 
            .I2(n1[29]), .I3(n30874), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1875_15_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n31760), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_31 (.CI(n30874), .I0(timer[29]), .I1(n1[29]), 
            .CO(n30875));
    SB_CARRY mod_5_add_1875_15 (.CI(n31760), .I0(n2697), .I1(n2720), .CO(n31761));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n31759), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_14 (.CI(n31759), .I0(n2698), .I1(n2720), .CO(n31760));
    SB_LUT4 mod_5_add_1875_13_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n31758), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_30_lut (.I0(one_wire_N_520[18]), .I1(timer[28]), 
            .I2(n1[28]), .I3(n30873), .O(n28_adj_4726)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1875_13 (.CI(n31758), .I0(n2699), .I1(n2720), .CO(n31759));
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1875_12_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n31757), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_12 (.CI(n31757), .I0(n2700), .I1(n2720), .CO(n31758));
    SB_LUT4 i4175_2_lut_3_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(bit_ctr[29]), 
            .I3(GND_net), .O(n8234));   // verilog/neopixel.v(22[26:36])
    defparam i4175_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 add_21_4_lut (.I0(GND_net), .I1(bit_ctr[2]), .I2(GND_net), 
            .I3(n30649), .O(n255[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1875_11_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n31756), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_11 (.CI(n31756), .I0(n2701), .I1(n2720), .CO(n31757));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n31755), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_12 (.CI(n30657), .I0(bit_ctr[10]), .I1(GND_net), .CO(n30658));
    SB_CARRY mod_5_add_1875_10 (.CI(n31755), .I0(n2702), .I1(n2720), .CO(n31756));
    SB_LUT4 mod_5_add_1875_9_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n31754), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_9 (.CI(n31754), .I0(n2703), .I1(n2720), .CO(n31755));
    SB_LUT4 mod_5_i471_3_lut_3_lut_4_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), 
            .I2(n27850), .I3(bit_ctr[29]), .O(n708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i471_3_lut_3_lut_4_lut.LUT_INIT = 16'hd222;
    SB_LUT4 i30096_4_lut (.I0(\state[1] ), .I1(n39270), .I2(n4983), .I3(state[0]), 
            .O(n21935));
    defparam i30096_4_lut.LUT_INIT = 16'h0f11;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i604_4_lut_4_lut (.I0(n36370), .I1(n9244), .I2(n838), 
            .I3(n807), .O(n905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i604_4_lut_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 add_21_33_lut (.I0(GND_net), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(n30678), .O(n255[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1875_8_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n31753), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_32_lut (.I0(GND_net), .I1(bit_ctr[30]), .I2(GND_net), 
            .I3(n30677), .O(n255[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_8 (.CI(n31753), .I0(n2704), .I1(n2720), .CO(n31754));
    SB_LUT4 mod_5_add_1875_7_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n31752), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_7 (.CI(n31752), .I0(n2705), .I1(n2720), .CO(n31753));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n31751), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_6 (.CI(n31751), .I0(n2706), .I1(n2720), .CO(n31752));
    SB_LUT4 mod_5_add_1875_5_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n31750), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_32 (.CI(n30677), .I0(bit_ctr[30]), .I1(GND_net), .CO(n30678));
    SB_CARRY mod_5_add_1875_5 (.CI(n31750), .I0(n2707), .I1(n2720), .CO(n31751));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n31749), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_4 (.CI(n31749), .I0(n2708), .I1(n2720), .CO(n31750));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(n2709), .I1(n2709), .I2(n40623), 
            .I3(n31748), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_3 (.CI(n31748), .I0(n2709), .I1(n40623), .CO(n31749));
    SB_LUT4 mod_5_add_1875_2_lut (.I0(bit_ctr[8]), .I1(bit_ctr[8]), .I2(n40623), 
            .I3(VCC_net), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(n40623), 
            .CO(n31748));
    SB_CARRY sub_14_add_2_30 (.CI(n30873), .I0(timer[28]), .I1(n1[28]), 
            .CO(n30874));
    SB_LUT4 sub_14_add_2_29_lut (.I0(one_wire_N_520[25]), .I1(timer[27]), 
            .I2(n1[27]), .I3(n30872), .O(n26_adj_4725)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n31747), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n31746), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_25 (.CI(n31746), .I0(n2787), .I1(n2819), .CO(n31747));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n31745), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_24 (.CI(n31745), .I0(n2788), .I1(n2819), .CO(n31746));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n31744), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_31_lut (.I0(GND_net), .I1(bit_ctr[29]), .I2(GND_net), 
            .I3(n30676), .O(n255[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_23 (.CI(n31744), .I0(n2789), .I1(n2819), .CO(n31745));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n31743), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_22 (.CI(n31743), .I0(n2790), .I1(n2819), .CO(n31744));
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n31742), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_21 (.CI(n31742), .I0(n2791), .I1(n2819), .CO(n31743));
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n31741), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_20 (.CI(n31741), .I0(n2792), .I1(n2819), .CO(n31742));
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n31740), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_i605_3_lut_4_lut (.I0(n36370), .I1(n9244), .I2(n838), 
            .I3(n807), .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_3_lut_4_lut.LUT_INIT = 16'hfe01;
    SB_DFF timer_1508__i0 (.Q(timer[0]), .C(clk32MHz), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY add_21_31 (.CI(n30676), .I0(bit_ctr[29]), .I1(GND_net), .CO(n30677));
    SB_LUT4 i26492_4_lut (.I0(n20592), .I1(n32422), .I2(n36426), .I3(state[0]), 
            .O(n14));
    defparam i26492_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i23_3_lut (.I0(n36426), .I1(n32422), .I2(state[0]), .I3(GND_net), 
            .O(n36470));
    defparam i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1569 (.I0(n27516), .I1(\state[1] ), .I2(n20592), 
            .I3(n36470), .O(n38147));
    defparam i3_4_lut_adj_1569.LUT_INIT = 16'heeef;
    SB_LUT4 i2_4_lut_adj_1570 (.I0(\state[1] ), .I1(n38147), .I2(start), 
            .I3(n36538), .O(n37680));
    defparam i2_4_lut_adj_1570.LUT_INIT = 16'h8c00;
    SB_CARRY mod_5_add_1942_19 (.CI(n31740), .I0(n2793), .I1(n2819), .CO(n31741));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n31739), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_11_lut (.I0(GND_net), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(n30656), .O(n255[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_18 (.CI(n31739), .I0(n2794), .I1(n2819), .CO(n31740));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n31738), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_11 (.CI(n30656), .I0(bit_ctr[9]), .I1(GND_net), .CO(n30657));
    SB_CARRY mod_5_add_1942_17 (.CI(n31738), .I0(n2795), .I1(n2819), .CO(n31739));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n31737), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_16 (.CI(n31737), .I0(n2796), .I1(n2819), .CO(n31738));
    SB_CARRY sub_14_add_2_29 (.CI(n30872), .I0(timer[27]), .I1(n1[27]), 
            .CO(n30873));
    SB_LUT4 add_21_30_lut (.I0(GND_net), .I1(bit_ctr[28]), .I2(GND_net), 
            .I3(n30675), .O(n255[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_30 (.CI(n30675), .I0(bit_ctr[28]), .I1(GND_net), .CO(n30676));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n31736), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_15 (.CI(n31736), .I0(n2797), .I1(n2819), .CO(n31737));
    SB_LUT4 sub_14_add_2_28_lut (.I0(one_wire_N_520[17]), .I1(timer[26]), 
            .I2(n1[26]), .I3(n30871), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i14_4_lut_adj_1571 (.I0(n2591), .I1(n2608), .I2(n2601), .I3(n2605), 
            .O(n36_adj_4764));
    defparam i14_4_lut_adj_1571.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_3_lut_adj_1572 (.I0(n2606), .I1(bit_ctr[9]), .I2(n2609), 
            .I3(GND_net), .O(n25_adj_4765));
    defparam i3_3_lut_adj_1572.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1573 (.I0(n2593), .I1(n2596), .I2(n2600), .I3(n2590), 
            .O(n34_adj_4766));
    defparam i12_4_lut_adj_1573.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1574 (.I0(n25_adj_4765), .I1(n36_adj_4764), .I2(n2594), 
            .I3(n2589), .O(n40_adj_4767));
    defparam i18_4_lut_adj_1574.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1575 (.I0(n2602), .I1(n2588), .I2(n2604), .I3(n2607), 
            .O(n38_adj_4768));
    defparam i16_4_lut_adj_1575.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n31735), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_28 (.CI(n30871), .I0(timer[26]), .I1(n1[26]), 
            .CO(n30872));
    SB_LUT4 sub_14_add_2_27_lut (.I0(GND_net), .I1(timer[25]), .I2(n1[25]), 
            .I3(n30870), .O(one_wire_N_520[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_10_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(n30655), .O(n255[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_14 (.CI(n31735), .I0(n2798), .I1(n2819), .CO(n31736));
    SB_CARRY sub_14_add_2_27 (.CI(n30870), .I0(timer[25]), .I1(n1[25]), 
            .CO(n30871));
    SB_LUT4 sub_14_add_2_26_lut (.I0(GND_net), .I1(timer[24]), .I2(n1[24]), 
            .I3(n30869), .O(one_wire_N_520[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_4 (.CI(n30649), .I0(bit_ctr[2]), .I1(GND_net), .CO(n30650));
    SB_LUT4 i17_3_lut (.I0(n2598), .I1(n34_adj_4766), .I2(n2603), .I3(GND_net), 
            .O(n39_adj_4769));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1576 (.I0(n2592), .I1(n2597), .I2(n2595), .I3(n2599), 
            .O(n37_adj_4770));
    defparam i15_4_lut_adj_1576.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1577 (.I0(n37_adj_4770), .I1(n39_adj_4769), .I2(n38_adj_4768), 
            .I3(n40_adj_4767), .O(n2621));
    defparam i21_4_lut_adj_1577.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_29_lut (.I0(GND_net), .I1(bit_ctr[27]), .I2(GND_net), 
            .I3(n30674), .O(n255[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_29 (.CI(n30674), .I0(bit_ctr[27]), .I1(GND_net), .CO(n30675));
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n31734), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_13 (.CI(n31734), .I0(n2799), .I1(n2819), .CO(n31735));
    SB_LUT4 timer_1508_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n31636), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_26 (.CI(n30869), .I0(timer[24]), .I1(n1[24]), 
            .CO(n30870));
    SB_LUT4 add_21_28_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(n30673), .O(n255[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_3_lut (.I0(GND_net), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(n30648), .O(n255[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1508_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n31635), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_25_lut (.I0(one_wire_N_520[14]), .I1(timer[23]), 
            .I2(n1[23]), .I3(n30868), .O(n29_adj_4729)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n31733), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_10 (.CI(n30655), .I0(bit_ctr[8]), .I1(GND_net), .CO(n30656));
    SB_CARRY mod_5_add_1942_12 (.CI(n31733), .I0(n2800), .I1(n2819), .CO(n31734));
    SB_CARRY timer_1508_add_4_32 (.CI(n31635), .I0(GND_net), .I1(timer[30]), 
            .CO(n31636));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n31732), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1508_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n31634), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1508_add_4_31 (.CI(n31634), .I0(GND_net), .I1(timer[29]), 
            .CO(n31635));
    SB_CARRY sub_14_add_2_25 (.CI(n30868), .I0(timer[23]), .I1(n1[23]), 
            .CO(n30869));
    SB_LUT4 timer_1508_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n31633), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_28 (.CI(n30673), .I0(bit_ctr[26]), .I1(GND_net), .CO(n30674));
    SB_CARRY mod_5_add_1942_11 (.CI(n31732), .I0(n2801), .I1(n2819), .CO(n31733));
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n31731), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1508_add_4_30 (.CI(n31633), .I0(GND_net), .I1(timer[28]), 
            .CO(n31634));
    SB_LUT4 add_21_27_lut (.I0(GND_net), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(n30672), .O(n255[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_10 (.CI(n31731), .I0(n2802), .I1(n2819), .CO(n31732));
    SB_LUT4 add_21_9_lut (.I0(GND_net), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(n30654), .O(n255[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_27 (.CI(n30672), .I0(bit_ctr[25]), .I1(GND_net), .CO(n30673));
    SB_LUT4 timer_1508_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n31632), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n31730), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1508_add_4_29 (.CI(n31632), .I0(GND_net), .I1(timer[27]), 
            .CO(n31633));
    SB_LUT4 add_21_26_lut (.I0(GND_net), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(n30671), .O(n255[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1508_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n31631), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_24_lut (.I0(GND_net), .I1(timer[22]), .I2(n1[22]), 
            .I3(n30867), .O(one_wire_N_520[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_26 (.CI(n30671), .I0(bit_ctr[24]), .I1(GND_net), .CO(n30672));
    SB_CARRY timer_1508_add_4_28 (.CI(n31631), .I0(GND_net), .I1(timer[26]), 
            .CO(n31632));
    SB_CARRY mod_5_add_1942_9 (.CI(n31730), .I0(n2803), .I1(n2819), .CO(n31731));
    SB_LUT4 timer_1508_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n31630), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n31729), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_8 (.CI(n31729), .I0(n2804), .I1(n2819), .CO(n31730));
    SB_CARRY sub_14_add_2_24 (.CI(n30867), .I0(timer[22]), .I1(n1[22]), 
            .CO(n30868));
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n31728), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_25_lut (.I0(GND_net), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(n30670), .O(n255[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1508_add_4_27 (.CI(n31630), .I0(GND_net), .I1(timer[25]), 
            .CO(n31631));
    SB_LUT4 timer_1508_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n31629), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_7 (.CI(n31728), .I0(n2805), .I1(n2819), .CO(n31729));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n31727), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1508_add_4_26 (.CI(n31629), .I0(GND_net), .I1(timer[24]), 
            .CO(n31630));
    SB_LUT4 timer_1508_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n31628), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1508_add_4_25 (.CI(n31628), .I0(GND_net), .I1(timer[23]), 
            .CO(n31629));
    SB_LUT4 timer_1508_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n31627), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_6 (.CI(n31727), .I0(n2806), .I1(n2819), .CO(n31728));
    SB_LUT4 sub_14_add_2_23_lut (.I0(one_wire_N_520[15]), .I1(timer[21]), 
            .I2(n1[21]), .I3(n30866), .O(n30_adj_4730)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY timer_1508_add_4_24 (.CI(n31627), .I0(GND_net), .I1(timer[22]), 
            .CO(n31628));
    SB_LUT4 timer_1508_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n31626), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_9 (.CI(n30654), .I0(bit_ctr[7]), .I1(GND_net), .CO(n30655));
    SB_CARRY timer_1508_add_4_23 (.CI(n31626), .I0(GND_net), .I1(timer[21]), 
            .CO(n31627));
    SB_LUT4 timer_1508_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n31625), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n31726), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_25 (.CI(n30670), .I0(bit_ctr[23]), .I1(GND_net), .CO(n30671));
    SB_CARRY sub_14_add_2_23 (.CI(n30866), .I0(timer[21]), .I1(n1[21]), 
            .CO(n30867));
    SB_CARRY timer_1508_add_4_22 (.CI(n31625), .I0(GND_net), .I1(timer[20]), 
            .CO(n31626));
    SB_LUT4 timer_1508_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n31624), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_5 (.CI(n31726), .I0(n2807), .I1(n2819), .CO(n31727));
    SB_LUT4 sub_14_add_2_22_lut (.I0(one_wire_N_520[12]), .I1(timer[20]), 
            .I2(n1[20]), .I3(n30865), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_22 (.CI(n30865), .I0(timer[20]), .I1(n1[20]), 
            .CO(n30866));
    SB_LUT4 sub_14_add_2_21_lut (.I0(one_wire_N_520[13]), .I1(timer[19]), 
            .I2(n1[19]), .I3(n30864), .O(n25)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_21 (.CI(n30864), .I0(timer[19]), .I1(n1[19]), 
            .CO(n30865));
    SB_CARRY timer_1508_add_4_21 (.CI(n31624), .I0(GND_net), .I1(timer[19]), 
            .CO(n31625));
    SB_LUT4 timer_1508_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n31623), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n31725), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_4 (.CI(n31725), .I0(n2808), .I1(n2819), .CO(n31726));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n40624), 
            .I3(n31724), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_add_2_20_lut (.I0(GND_net), .I1(timer[18]), .I2(n1[18]), 
            .I3(n30863), .O(one_wire_N_520[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1508_add_4_20 (.CI(n31623), .I0(GND_net), .I1(timer[18]), 
            .CO(n31624));
    SB_CARRY sub_14_add_2_20 (.CI(n30863), .I0(timer[18]), .I1(n1[18]), 
            .CO(n30864));
    SB_CARRY mod_5_add_1942_3 (.CI(n31724), .I0(n2809), .I1(n40624), .CO(n31725));
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n40624), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 timer_1508_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n31622), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1508_add_4_19 (.CI(n31622), .I0(GND_net), .I1(timer[17]), 
            .CO(n31623));
    SB_LUT4 sub_14_add_2_19_lut (.I0(GND_net), .I1(timer[17]), .I2(n1[17]), 
            .I3(n30862), .O(one_wire_N_520[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_753_Mux_0_i3_3_lut_3_lut (.I0(\neo_pixel_transmitter.done ), 
            .I1(start), .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_577 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_753_Mux_0_i3_3_lut_3_lut.LUT_INIT = 16'ha1a1;
    SB_LUT4 bit_ctr_0__bdd_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[10]), 
            .I2(neopxl_color[11]), .I3(bit_ctr[1]), .O(n40840));
    defparam bit_ctr_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n40840_bdd_4_lut (.I0(n40840), .I1(neopxl_color[9]), .I2(neopxl_color[8]), 
            .I3(bit_ctr[1]), .O(n38446));
    defparam n40840_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_30777 (.I0(bit_ctr[0]), .I1(neopxl_color[14]), 
            .I2(neopxl_color[15]), .I3(bit_ctr[1]), .O(n40834));
    defparam bit_ctr_0__bdd_4_lut_30777.LUT_INIT = 16'he4aa;
    SB_LUT4 n40834_bdd_4_lut (.I0(n40834), .I1(neopxl_color[13]), .I2(neopxl_color[12]), 
            .I3(bit_ctr[1]), .O(n38449));
    defparam n40834_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 bit_ctr_0__bdd_4_lut_30772 (.I0(bit_ctr[0]), .I1(neopxl_color[2]), 
            .I2(neopxl_color[3]), .I3(bit_ctr[1]), .O(n40822));
    defparam bit_ctr_0__bdd_4_lut_30772.LUT_INIT = 16'he4aa;
    SB_LUT4 n40822_bdd_4_lut (.I0(n40822), .I1(neopxl_color[1]), .I2(neopxl_color[0]), 
            .I3(bit_ctr[1]), .O(n38455));
    defparam n40822_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY sub_14_add_2_19 (.CI(n30862), .I0(timer[17]), .I1(n1[17]), 
            .CO(n30863));
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n40624), 
            .CO(n31724));
    SB_LUT4 i14_4_lut_adj_1578 (.I0(n3004), .I1(n2989), .I2(n2990), .I3(n3007), 
            .O(n40_adj_4772));
    defparam i14_4_lut_adj_1578.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1579 (.I0(n3006), .I1(n2984), .I2(n2988), .I3(n2986), 
            .O(n44_adj_4773));
    defparam i18_4_lut_adj_1579.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1580 (.I0(n3008), .I1(n3003), .I2(n2994), .I3(n3002), 
            .O(n42_adj_4774));
    defparam i16_4_lut_adj_1580.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1581 (.I0(n2999), .I1(n3000), .I2(n2992), .I3(n2997), 
            .O(n43_adj_4775));
    defparam i17_4_lut_adj_1581.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_18_lut (.I0(GND_net), .I1(timer[16]), .I2(n1[16]), 
            .I3(n30861), .O(one_wire_N_520[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_18 (.CI(n30861), .I0(timer[16]), .I1(n1[16]), 
            .CO(n30862));
    SB_LUT4 sub_14_add_2_17_lut (.I0(GND_net), .I1(timer[15]), .I2(n1[15]), 
            .I3(n30860), .O(one_wire_N_520[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_24_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(n30669), .O(n255[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15_4_lut_adj_1582 (.I0(n2996), .I1(n2985), .I2(n2995), .I3(n2987), 
            .O(n41_adj_4777));
    defparam i15_4_lut_adj_1582.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut_adj_1583 (.I0(n3001), .I1(n2993), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_4778));
    defparam i12_2_lut_adj_1583.LUT_INIT = 16'heeee;
    SB_LUT4 i20_3_lut (.I0(n2998), .I1(n40_adj_4772), .I2(n2991), .I3(GND_net), 
            .O(n46_adj_4779));
    defparam i20_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i24_4_lut (.I0(n41_adj_4777), .I1(n43_adj_4775), .I2(n42_adj_4774), 
            .I3(n44_adj_4773), .O(n50));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_3_lut (.I0(n3005), .I1(bit_ctr[5]), .I2(n3009), .I3(GND_net), 
            .O(n37_adj_4780));
    defparam i11_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut_adj_1584 (.I0(n2003), .I1(n2008), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4782));
    defparam i2_2_lut_adj_1584.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1585 (.I0(n1996), .I1(n1998), .I2(n2006), .I3(n2007), 
            .O(n28_adj_4783));
    defparam i12_4_lut_adj_1585.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut_adj_1586 (.I0(n37_adj_4780), .I1(n50), .I2(n46_adj_4779), 
            .I3(n38_adj_4778), .O(n3017));
    defparam i25_4_lut_adj_1586.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1587 (.I0(n1997), .I1(n1999), .I2(n2005), .I3(n2000), 
            .O(n26_adj_4784));
    defparam i10_4_lut_adj_1587.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1588 (.I0(n1994), .I1(n2001), .I2(n2004), .I3(n1995), 
            .O(n27_adj_4785));
    defparam i11_4_lut_adj_1588.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(bit_ctr[15]), .I1(n18_adj_4782), .I2(n2002), 
            .I3(n2009), .O(n25_adj_4786));
    defparam i9_4_lut.LUT_INIT = 16'hfefc;
    SB_CARRY sub_14_add_2_17 (.CI(n30860), .I0(timer[15]), .I1(n1[15]), 
            .CO(n30861));
    SB_LUT4 i15_4_lut_adj_1589 (.I0(n25_adj_4786), .I1(n27_adj_4785), .I2(n26_adj_4784), 
            .I3(n28_adj_4783), .O(n2027));
    defparam i15_4_lut_adj_1589.LUT_INIT = 16'hfffe;
    SB_LUT4 i30605_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40632));
    defparam i30605_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11_4_lut_adj_1590 (.I0(n1895), .I1(n1902), .I2(n1899), .I3(n1897), 
            .O(n26_adj_4787));
    defparam i11_4_lut_adj_1590.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_16_lut (.I0(GND_net), .I1(timer[14]), .I2(n1[14]), 
            .I3(n30859), .O(one_wire_N_520[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_3_lut (.I0(n1907), .I1(bit_ctr[16]), .I2(n1909), .I3(GND_net), 
            .O(n19_adj_4789));
    defparam i4_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut_adj_1591 (.I0(n1908), .I1(n1900), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4790));
    defparam i1_2_lut_adj_1591.LUT_INIT = 16'heeee;
    SB_CARRY add_21_24 (.CI(n30669), .I0(bit_ctr[22]), .I1(GND_net), .CO(n30670));
    SB_CARRY sub_14_add_2_16 (.CI(n30859), .I0(timer[14]), .I1(n1[14]), 
            .CO(n30860));
    SB_LUT4 sub_14_add_2_15_lut (.I0(GND_net), .I1(timer[13]), .I2(n1[13]), 
            .I3(n30858), .O(one_wire_N_520[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_15 (.CI(n30858), .I0(timer[13]), .I1(n1[13]), 
            .CO(n30859));
    SB_LUT4 i9_4_lut_adj_1592 (.I0(n1904), .I1(n1901), .I2(n1906), .I3(n1898), 
            .O(n24_adj_4792));
    defparam i9_4_lut_adj_1592.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1593 (.I0(n19_adj_4789), .I1(n26_adj_4787), .I2(n1905), 
            .I3(n1903), .O(n28_adj_4793));
    defparam i13_4_lut_adj_1593.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1594 (.I0(n1896), .I1(n28_adj_4793), .I2(n24_adj_4792), 
            .I3(n16_adj_4790), .O(n1928));
    defparam i14_4_lut_adj_1594.LUT_INIT = 16'hfffe;
    SB_LUT4 i30604_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40631));
    defparam i30604_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n31723), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_14_lut (.I0(GND_net), .I1(timer[12]), .I2(n1[12]), 
            .I3(n30857), .O(one_wire_N_520[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1508_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n31621), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_14 (.CI(n30857), .I0(timer[12]), .I1(n1[12]), 
            .CO(n30858));
    SB_LUT4 mod_5_add_2009_26_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n31722), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1508_add_4_18 (.CI(n31621), .I0(GND_net), .I1(timer[16]), 
            .CO(n31622));
    SB_CARRY mod_5_add_2009_26 (.CI(n31722), .I0(n2886), .I1(n2918), .CO(n31723));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n30856), .O(one_wire_N_520[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2009_25_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n31721), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_25 (.CI(n31721), .I0(n2887), .I1(n2918), .CO(n31722));
    SB_LUT4 mod_5_add_2009_24_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n31720), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_24 (.CI(n31720), .I0(n2888), .I1(n2918), .CO(n31721));
    SB_LUT4 mod_5_add_2009_23_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n31719), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1508_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n31620), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1508_add_4_17 (.CI(n31620), .I0(GND_net), .I1(timer[15]), 
            .CO(n31621));
    SB_CARRY mod_5_add_2009_23 (.CI(n31719), .I0(n2889), .I1(n2918), .CO(n31720));
    SB_LUT4 timer_1508_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n31619), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1508_add_4_16 (.CI(n31619), .I0(GND_net), .I1(timer[14]), 
            .CO(n31620));
    SB_LUT4 mod_5_add_2009_22_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n31718), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1508_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n31618), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_13 (.CI(n30856), .I0(timer[11]), .I1(n1[11]), 
            .CO(n30857));
    SB_CARRY mod_5_add_2009_22 (.CI(n31718), .I0(n2890), .I1(n2918), .CO(n31719));
    SB_CARRY timer_1508_add_4_15 (.CI(n31618), .I0(GND_net), .I1(timer[13]), 
            .CO(n31619));
    SB_LUT4 timer_1508_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n31617), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10_4_lut_adj_1595 (.I0(n1806), .I1(n1803), .I2(n1798), .I3(n1805), 
            .O(n24_adj_4796));
    defparam i10_4_lut_adj_1595.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1596 (.I0(n1808), .I1(n1804), .I2(n1802), .I3(n1807), 
            .O(n22_adj_4797));
    defparam i8_4_lut_adj_1596.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1597 (.I0(n1800), .I1(n1799), .I2(n1797), .I3(n1801), 
            .O(n23_adj_4798));
    defparam i9_4_lut_adj_1597.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut (.I0(n1796), .I1(bit_ctr[17]), .I2(n1809), .I3(GND_net), 
            .O(n21_adj_4799));
    defparam i7_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 mod_5_add_2009_21_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n31717), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1508_add_4_14 (.CI(n31617), .I0(GND_net), .I1(timer[12]), 
            .CO(n31618));
    SB_LUT4 i13_4_lut_adj_1598 (.I0(n21_adj_4799), .I1(n23_adj_4798), .I2(n22_adj_4797), 
            .I3(n24_adj_4796), .O(n1829));
    defparam i13_4_lut_adj_1598.LUT_INIT = 16'hfffe;
    SB_LUT4 i30603_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40630));
    defparam i30603_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(clk32MHz), .E(n21935), 
            .D(n255[27]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(clk32MHz), .E(n21935), 
            .D(n255[26]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(clk32MHz), .E(n21935), 
            .D(n255[25]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_2009_21 (.CI(n31717), .I0(n2891), .I1(n2918), .CO(n31718));
    SB_LUT4 timer_1508_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n31616), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1508_add_4_13 (.CI(n31616), .I0(GND_net), .I1(timer[11]), 
            .CO(n31617));
    SB_DFFESR bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(clk32MHz), .E(n21935), 
            .D(n255[24]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n30855), .O(one_wire_N_520[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_12 (.CI(n30855), .I0(timer[10]), .I1(n1[10]), 
            .CO(n30856));
    SB_LUT4 mod_5_add_2009_20_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n31716), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1508_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n31615), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2009_20 (.CI(n31716), .I0(n2892), .I1(n2918), .CO(n31717));
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1400), .I1(n1400), .I2(n1433), 
            .I3(n32019), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1508_add_4_12 (.CI(n31615), .I0(GND_net), .I1(timer[10]), 
            .CO(n31616));
    SB_LUT4 mod_5_add_1004_11_lut (.I0(n1401), .I1(n1401), .I2(n1433), 
            .I3(n32018), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n30854), .O(one_wire_N_520[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_11 (.CI(n32018), .I0(n1401), .I1(n1433), .CO(n32019));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(n1402), .I1(n1402), .I2(n1433), 
            .I3(n32017), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_10 (.CI(n32017), .I0(n1402), .I1(n1433), .CO(n32018));
    SB_LUT4 mod_5_add_1004_9_lut (.I0(n1403), .I1(n1403), .I2(n1433), 
            .I3(n32016), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_9 (.CI(n32016), .I0(n1403), .I1(n1433), .CO(n32017));
    SB_LUT4 mod_5_add_1004_8_lut (.I0(n1404), .I1(n1404), .I2(n1433), 
            .I3(n32015), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_8 (.CI(n32015), .I0(n1404), .I1(n1433), .CO(n32016));
    SB_LUT4 mod_5_add_1004_7_lut (.I0(n1405), .I1(n1405), .I2(n1433), 
            .I3(n32014), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_7 (.CI(n32014), .I0(n1405), .I1(n1433), .CO(n32015));
    SB_LUT4 mod_5_add_1004_6_lut (.I0(n1406), .I1(n1406), .I2(n1433), 
            .I3(n32013), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_6 (.CI(n32013), .I0(n1406), .I1(n1433), .CO(n32014));
    SB_LUT4 timer_1508_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n31614), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1004_5_lut (.I0(n1407), .I1(n1407), .I2(n1433), 
            .I3(n32012), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1508_add_4_11 (.CI(n31614), .I0(GND_net), .I1(timer[9]), 
            .CO(n31615));
    SB_CARRY mod_5_add_1004_5 (.CI(n32012), .I0(n1407), .I1(n1433), .CO(n32013));
    SB_LUT4 mod_5_add_1004_4_lut (.I0(n1408), .I1(n1408), .I2(n1433), 
            .I3(n32011), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_4 (.CI(n32011), .I0(n1408), .I1(n1433), .CO(n32012));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(n1409), .I1(n1409), .I2(n40626), 
            .I3(n32010), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i3_3_lut_adj_1599 (.I0(bit_ctr[18]), .I1(n1704), .I2(n1709), 
            .I3(GND_net), .O(n16_adj_4803));
    defparam i3_3_lut_adj_1599.LUT_INIT = 16'hecec;
    SB_CARRY mod_5_add_1004_3 (.CI(n32010), .I0(n1409), .I1(n40626), .CO(n32011));
    SB_LUT4 mod_5_add_1004_2_lut (.I0(bit_ctr[21]), .I1(bit_ctr[21]), .I2(n40626), 
            .I3(VCC_net), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY sub_14_add_2_11 (.CI(n30854), .I0(timer[9]), .I1(n1[9]), 
            .CO(n30855));
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(n40626), 
            .CO(n32010));
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n30853), .O(one_wire_N_520[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n32009), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_10 (.CI(n30853), .I0(timer[8]), .I1(n1[8]), 
            .CO(n30854));
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n32008), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_8 (.CI(n32008), .I0(n1104), .I1(n1136), .CO(n32009));
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n32007), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_7 (.CI(n32007), .I0(n1105), .I1(n1136), .CO(n32008));
    SB_LUT4 mod_5_add_2009_19_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n31715), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1508_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n31613), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n32006), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_6 (.CI(n32006), .I0(n1106), .I1(n1136), .CO(n32007));
    SB_LUT4 i9_4_lut_adj_1600 (.I0(n1707), .I1(n1697), .I2(n1702), .I3(n1699), 
            .O(n22_adj_4805));
    defparam i9_4_lut_adj_1600.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1601 (.I0(n1706), .I1(n1701), .I2(n1708), .I3(GND_net), 
            .O(n20_adj_4806));
    defparam i7_3_lut_adj_1601.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1602 (.I0(n1703), .I1(n22_adj_4805), .I2(n16_adj_4803), 
            .I3(n1698), .O(n24_adj_4807));
    defparam i11_4_lut_adj_1602.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1603 (.I0(n1705), .I1(n24_adj_4807), .I2(n20_adj_4806), 
            .I3(n1700), .O(n1730));
    defparam i12_4_lut_adj_1603.LUT_INIT = 16'hfffe;
    SB_LUT4 i30602_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40629));
    defparam i30602_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_4_lut_adj_1604 (.I0(n1608), .I1(n1606), .I2(n1604), .I3(n1603), 
            .O(n20_adj_4809));
    defparam i8_4_lut_adj_1604.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1605 (.I0(bit_ctr[19]), .I1(n1602), .I2(n1609), 
            .I3(GND_net), .O(n13_adj_4810));
    defparam i1_3_lut_adj_1605.LUT_INIT = 16'hecec;
    SB_LUT4 i6_2_lut (.I0(n1598), .I1(n1600), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4811));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1606 (.I0(n13_adj_4810), .I1(n20_adj_4809), .I2(n1605), 
            .I3(n1599), .O(n22_adj_4812));
    defparam i10_4_lut_adj_1606.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1607 (.I0(n1601), .I1(n22_adj_4812), .I2(n18_adj_4811), 
            .I3(n1607), .O(n1631));
    defparam i11_4_lut_adj_1607.LUT_INIT = 16'hfffe;
    SB_LUT4 i30601_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40628));
    defparam i30601_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2009_19 (.CI(n31715), .I0(n2893), .I1(n2918), .CO(n31716));
    SB_CARRY timer_1508_add_4_10 (.CI(n31613), .I0(GND_net), .I1(timer[8]), 
            .CO(n31614));
    SB_CARRY add_21_3 (.CI(n30648), .I0(bit_ctr[1]), .I1(GND_net), .CO(n30649));
    SB_DFFESR bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(clk32MHz), .E(n21935), 
            .D(n255[23]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2009_18_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n31714), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1508_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n31612), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1508_add_4_9 (.CI(n31612), .I0(GND_net), .I1(timer[7]), 
            .CO(n31613));
    SB_LUT4 add_21_8_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(n30653), .O(n255[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_23_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(n30668), .O(n255[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_23 (.CI(n30668), .I0(bit_ctr[21]), .I1(GND_net), .CO(n30669));
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n30852), .O(one_wire_N_520[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_9 (.CI(n30852), .I0(timer[7]), .I1(n1[7]), .CO(n30853));
    SB_LUT4 add_21_22_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(n30667), .O(n255[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_8_lut (.I0(one_wire_N_520[9]), .I1(timer[6]), .I2(n1[6]), 
            .I3(n30851), .O(n9_adj_4732)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_21_2_lut (.I0(GND_net), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n255[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_22 (.CI(n30667), .I0(bit_ctr[20]), .I1(GND_net), .CO(n30668));
    SB_LUT4 i19120_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(GND_net), .I3(GND_net), .O(n27516));
    defparam i19120_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n32005), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_5 (.CI(n32005), .I0(n1107), .I1(n1136), .CO(n32006));
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n32004), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_4 (.CI(n32004), .I0(n1108), .I1(n1136), .CO(n32005));
    SB_CARRY mod_5_add_2009_18 (.CI(n31714), .I0(n2894), .I1(n2918), .CO(n31715));
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n40627), 
            .I3(n32003), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_3 (.CI(n32003), .I0(n1109), .I1(n40627), .CO(n32004));
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n40627), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 timer_1508_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n31611), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n40627), 
            .CO(n32003));
    SB_CARRY add_21_8 (.CI(n30653), .I0(bit_ctr[6]), .I1(GND_net), .CO(n30654));
    SB_LUT4 add_21_7_lut (.I0(GND_net), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(n30652), .O(n255[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_8 (.CI(n30851), .I0(timer[6]), .I1(n1[6]), .CO(n30852));
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n31992), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_17_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n31713), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_12_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n31991), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n30850), .O(one_wire_N_520[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_12 (.CI(n31991), .I0(n1500), .I1(n1532), .CO(n31992));
    SB_LUT4 mod_5_add_1071_11_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n31990), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_21_lut (.I0(GND_net), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(n30666), .O(n255[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_11 (.CI(n31990), .I0(n1501), .I1(n1532), .CO(n31991));
    SB_CARRY sub_14_add_2_7 (.CI(n30850), .I0(timer[5]), .I1(n1[5]), .CO(n30851));
    SB_LUT4 mod_5_add_1071_10_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n31989), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_10 (.CI(n31989), .I0(n1502), .I1(n1532), .CO(n31990));
    SB_LUT4 mod_5_add_1071_9_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n31988), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_9 (.CI(n31988), .I0(n1503), .I1(n1532), .CO(n31989));
    SB_LUT4 mod_5_add_1071_8_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n31987), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_8 (.CI(n31987), .I0(n1504), .I1(n1532), .CO(n31988));
    SB_LUT4 mod_5_add_1071_7_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n31986), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_7 (.CI(n31986), .I0(n1505), .I1(n1532), .CO(n31987));
    SB_LUT4 mod_5_add_1071_6_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n31985), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_6 (.CI(n31985), .I0(n1506), .I1(n1532), .CO(n31986));
    SB_LUT4 mod_5_add_1071_5_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n31984), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_5 (.CI(n31984), .I0(n1507), .I1(n1532), .CO(n31985));
    SB_LUT4 mod_5_add_1071_4_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n31983), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_4 (.CI(n31983), .I0(n1508), .I1(n1532), .CO(n31984));
    SB_LUT4 mod_5_add_1071_3_lut (.I0(n1509), .I1(n1509), .I2(n40628), 
            .I3(n31982), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_3 (.CI(n31982), .I0(n1509), .I1(n40628), .CO(n31983));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(bit_ctr[20]), .I1(bit_ctr[20]), .I2(n40628), 
            .I3(VCC_net), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(n40628), 
            .CO(n31982));
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n31981), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n31980), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n30849), .O(one_wire_N_520[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_13 (.CI(n31980), .I0(n1599), .I1(n1631), .CO(n31981));
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n31979), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_12 (.CI(n31979), .I0(n1600), .I1(n1631), .CO(n31980));
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n31978), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_11 (.CI(n31978), .I0(n1601), .I1(n1631), .CO(n31979));
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n31977), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_10 (.CI(n31977), .I0(n1602), .I1(n1631), .CO(n31978));
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n31976), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_9 (.CI(n31976), .I0(n1603), .I1(n1631), .CO(n31977));
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n31975), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_8 (.CI(n31975), .I0(n1604), .I1(n1631), .CO(n31976));
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n31974), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_7 (.CI(n31974), .I0(n1605), .I1(n1631), .CO(n31975));
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n31973), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_6 (.CI(n31973), .I0(n1606), .I1(n1631), .CO(n31974));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n31972), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_5 (.CI(n31972), .I0(n1607), .I1(n1631), .CO(n31973));
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n31971), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_4 (.CI(n31971), .I0(n1608), .I1(n1631), .CO(n31972));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n40629), 
            .I3(n31970), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_3 (.CI(n31970), .I0(n1609), .I1(n40629), .CO(n31971));
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n40629), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n40629), 
            .CO(n31970));
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n31969), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n31968), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_14 (.CI(n31968), .I0(n1698), .I1(n1730), .CO(n31969));
    SB_CARRY sub_14_add_2_6 (.CI(n30849), .I0(timer[4]), .I1(n1[4]), .CO(n30850));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n31967), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_13 (.CI(n31967), .I0(n1699), .I1(n1730), .CO(n31968));
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n31966), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_17 (.CI(n31713), .I0(n2895), .I1(n2918), .CO(n31714));
    SB_CARRY mod_5_add_1205_12 (.CI(n31966), .I0(n1700), .I1(n1730), .CO(n31967));
    SB_CARRY timer_1508_add_4_8 (.CI(n31611), .I0(GND_net), .I1(timer[6]), 
            .CO(n31612));
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n31965), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_11 (.CI(n31965), .I0(n1701), .I1(n1730), .CO(n31966));
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n31964), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n30848), .O(one_wire_N_520[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_10 (.CI(n31964), .I0(n1702), .I1(n1730), .CO(n31965));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n31963), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_9 (.CI(n31963), .I0(n1703), .I1(n1730), .CO(n31964));
    SB_LUT4 timer_1508_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n31610), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n31962), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_8 (.CI(n31962), .I0(n1704), .I1(n1730), .CO(n31963));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n31961), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_7 (.CI(n31961), .I0(n1705), .I1(n1730), .CO(n31962));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n31960), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_21 (.CI(n30666), .I0(bit_ctr[19]), .I1(GND_net), .CO(n30667));
    SB_CARRY mod_5_add_1205_6 (.CI(n31960), .I0(n1706), .I1(n1730), .CO(n31961));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n31959), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_5 (.CI(n31959), .I0(n1707), .I1(n1730), .CO(n31960));
    SB_CARRY sub_14_add_2_5 (.CI(n30848), .I0(timer[3]), .I1(n1[3]), .CO(n30849));
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n31958), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_4 (.CI(n31958), .I0(n1708), .I1(n1730), .CO(n31959));
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n40630), 
            .I3(n31957), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_20_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(n30665), .O(n255[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1205_3 (.CI(n31957), .I0(n1709), .I1(n40630), .CO(n31958));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n40630), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n40630), 
            .CO(n31957));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n31956), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n31955), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_15 (.CI(n31955), .I0(n1797), .I1(n1829), .CO(n31956));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n31954), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_14 (.CI(n31954), .I0(n1798), .I1(n1829), .CO(n31955));
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n31953), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_13 (.CI(n31953), .I0(n1799), .I1(n1829), .CO(n31954));
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n31952), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_12 (.CI(n31952), .I0(n1800), .I1(n1829), .CO(n31953));
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n31951), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_11 (.CI(n31951), .I0(n1801), .I1(n1829), .CO(n31952));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n31950), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_10 (.CI(n31950), .I0(n1802), .I1(n1829), .CO(n31951));
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n31949), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_9 (.CI(n31949), .I0(n1803), .I1(n1829), .CO(n31950));
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n31948), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_8 (.CI(n31948), .I0(n1804), .I1(n1829), .CO(n31949));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n31947), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_7 (.CI(n31947), .I0(n1805), .I1(n1829), .CO(n31948));
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n31946), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_6 (.CI(n31946), .I0(n1806), .I1(n1829), .CO(n31947));
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n31945), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_5 (.CI(n31945), .I0(n1807), .I1(n1829), .CO(n31946));
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n31944), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_4 (.CI(n31944), .I0(n1808), .I1(n1829), .CO(n31945));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n40631), 
            .I3(n31943), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_3 (.CI(n31943), .I0(n1809), .I1(n40631), .CO(n31944));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n40631), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n40631), 
            .CO(n31943));
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n31942), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_16_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n31941), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_16 (.CI(n31941), .I0(n1896), .I1(n1928), .CO(n31942));
    SB_LUT4 mod_5_add_1339_15_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n31940), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_15 (.CI(n31940), .I0(n1897), .I1(n1928), .CO(n31941));
    SB_LUT4 mod_5_add_1339_14_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n31939), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_14 (.CI(n31939), .I0(n1898), .I1(n1928), .CO(n31940));
    SB_LUT4 mod_5_add_1339_13_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n31938), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_13 (.CI(n31938), .I0(n1899), .I1(n1928), .CO(n31939));
    SB_LUT4 mod_5_add_1339_12_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n31937), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_12 (.CI(n31937), .I0(n1900), .I1(n1928), .CO(n31938));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n31936), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_11 (.CI(n31936), .I0(n1901), .I1(n1928), .CO(n31937));
    SB_LUT4 mod_5_add_1339_10_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n31935), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_10 (.CI(n31935), .I0(n1902), .I1(n1928), .CO(n31936));
    SB_LUT4 mod_5_add_1339_9_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n31934), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_9 (.CI(n31934), .I0(n1903), .I1(n1928), .CO(n31935));
    SB_LUT4 mod_5_add_1339_8_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n31933), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_8 (.CI(n31933), .I0(n1904), .I1(n1928), .CO(n31934));
    SB_LUT4 mod_5_add_1339_7_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n31932), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_7 (.CI(n31932), .I0(n1905), .I1(n1928), .CO(n31933));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n31931), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_6 (.CI(n31931), .I0(n1906), .I1(n1928), .CO(n31932));
    SB_LUT4 mod_5_add_1339_5_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n31930), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i30083_2_lut (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n35558));
    defparam i30083_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_4_lut_adj_1608 (.I0(n1506), .I1(n1503), .I2(n1500), .I3(n1501), 
            .O(n18_adj_4816));
    defparam i7_4_lut_adj_1608.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1609 (.I0(n1504), .I1(n18_adj_4816), .I2(n1502), 
            .I3(n1499), .O(n20_adj_4817));
    defparam i9_4_lut_adj_1609.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1610 (.I0(bit_ctr[20]), .I1(n1505), .I2(n1509), 
            .I3(GND_net), .O(n15_adj_4818));
    defparam i4_3_lut_adj_1610.LUT_INIT = 16'hecec;
    SB_LUT4 i10_4_lut_adj_1611 (.I0(n15_adj_4818), .I1(n20_adj_4817), .I2(n1508), 
            .I3(n1507), .O(n1532));
    defparam i10_4_lut_adj_1611.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1339_5 (.CI(n31930), .I0(n1907), .I1(n1928), .CO(n31931));
    SB_LUT4 mod_5_add_1339_4_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n31929), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_4 (.CI(n31929), .I0(n1908), .I1(n1928), .CO(n31930));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(n1909), .I1(n1909), .I2(n40632), 
            .I3(n31928), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1339_3 (.CI(n31928), .I0(n1909), .I1(n40632), .CO(n31929));
    SB_LUT4 mod_5_add_1339_2_lut (.I0(bit_ctr[16]), .I1(bit_ctr[16]), .I2(n40632), 
            .I3(VCC_net), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(n40632), 
            .CO(n31928));
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n31927), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_17_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n31926), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_17 (.CI(n31926), .I0(n1995), .I1(n2027), .CO(n31927));
    SB_LUT4 mod_5_add_1406_16_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n31925), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_16 (.CI(n31925), .I0(n1996), .I1(n2027), .CO(n31926));
    SB_LUT4 mod_5_add_1406_15_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n31924), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_15 (.CI(n31924), .I0(n1997), .I1(n2027), .CO(n31925));
    SB_LUT4 mod_5_add_1406_14_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n31923), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_14 (.CI(n31923), .I0(n1998), .I1(n2027), .CO(n31924));
    SB_LUT4 mod_5_add_1406_13_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n31922), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_13 (.CI(n31922), .I0(n1999), .I1(n2027), .CO(n31923));
    SB_LUT4 mod_5_add_1406_12_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n31921), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_12 (.CI(n31921), .I0(n2000), .I1(n2027), .CO(n31922));
    SB_LUT4 mod_5_add_1406_11_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n31920), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_11 (.CI(n31920), .I0(n2001), .I1(n2027), .CO(n31921));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n31919), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_10 (.CI(n31919), .I0(n2002), .I1(n2027), .CO(n31920));
    SB_LUT4 mod_5_add_1406_9_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n31918), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n30847), .O(one_wire_N_520[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1612 (.I0(one_wire_N_520[4]), .I1(one_wire_N_520[3]), 
            .I2(n35558), .I3(n32530), .O(n111));
    defparam i1_4_lut_adj_1612.LUT_INIT = 16'h5155;
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk32MHz), .D(n22814));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk32MHz), .D(n22813));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk32MHz), .D(n22812));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk32MHz), .D(n22811));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk32MHz), .D(n22810));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk32MHz), .D(n22809));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk32MHz), .D(n22808));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk32MHz), .D(n22807));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 bit_ctr_0__bdd_4_lut_30762 (.I0(bit_ctr[0]), .I1(neopxl_color[22]), 
            .I2(neopxl_color[23]), .I3(bit_ctr[1]), .O(n40726));
    defparam bit_ctr_0__bdd_4_lut_30762.LUT_INIT = 16'he4aa;
    SB_LUT4 i30600_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40627));
    defparam i30600_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk32MHz), .D(n22806));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1406_9 (.CI(n31918), .I0(n2003), .I1(n2027), .CO(n31919));
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk32MHz), .D(n22805));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2009_16_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n31712), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk32MHz), .D(n22804));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY timer_1508_add_4_7 (.CI(n31610), .I0(GND_net), .I1(timer[5]), 
            .CO(n31611));
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk32MHz), .D(n22803));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk32MHz), .D(n22802));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk32MHz), .D(n22801));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk32MHz), .D(n22800));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk32MHz), .D(n22799));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY sub_14_add_2_4 (.CI(n30847), .I0(timer[2]), .I1(n1[2]), .CO(n30848));
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk32MHz), .D(n22798));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk32MHz), .D(n22797));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk32MHz), .D(n22796));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk32MHz), .D(n22795));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk32MHz), .D(n22794));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk32MHz), .D(n22793));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk32MHz), .D(n22792));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk32MHz), .D(n22791));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk32MHz), .D(n22790));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk32MHz), .D(n22789));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk32MHz), .D(n22788));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk32MHz), .D(n22787));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk32MHz), .D(n22786));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk32MHz), .D(n22785));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk32MHz), .D(n22784));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 timer_1508_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n31609), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_3_lut (.I0(n4_adj_4819), .I1(timer[1]), .I2(n1[1]), 
            .I3(n30846), .O(n32530)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_2009_16 (.CI(n31712), .I0(n2896), .I1(n2918), .CO(n31713));
    SB_CARRY timer_1508_add_4_6 (.CI(n31609), .I0(GND_net), .I1(timer[4]), 
            .CO(n31610));
    SB_CARRY sub_14_add_2_3 (.CI(n30846), .I0(timer[1]), .I1(n1[1]), .CO(n30847));
    SB_LUT4 n40726_bdd_4_lut (.I0(n40726), .I1(neopxl_color[21]), .I2(neopxl_color[20]), 
            .I3(bit_ctr[1]), .O(n40729));
    defparam n40726_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_1508_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n31608), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_2_lut (.I0(one_wire_N_520[2]), .I1(timer[0]), .I2(n1[0]), 
            .I3(VCC_net), .O(n4_adj_4819)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_2009_15_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n31711), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1508_add_4_5 (.CI(n31608), .I0(GND_net), .I1(timer[3]), 
            .CO(n31609));
    SB_LUT4 timer_1508_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n31607), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_15 (.CI(n31711), .I0(n2897), .I1(n2918), .CO(n31712));
    SB_CARRY timer_1508_add_4_4 (.CI(n31607), .I0(GND_net), .I1(timer[2]), 
            .CO(n31608));
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n30846));
    SB_LUT4 timer_1508_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n31606), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_20 (.CI(n30665), .I0(bit_ctr[18]), .I1(GND_net), .CO(n30666));
    SB_LUT4 mod_5_add_1406_8_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n31917), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_14_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n31710), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_14 (.CI(n31710), .I0(n2898), .I1(n2918), .CO(n31711));
    SB_CARRY timer_1508_add_4_3 (.CI(n31606), .I0(GND_net), .I1(timer[1]), 
            .CO(n31607));
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n31142), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n31141), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n31141), .I0(n1203), .I1(n1235), .CO(n31142));
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n31140), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_8 (.CI(n31140), .I0(n1204), .I1(n1235), .CO(n31141));
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n31139), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_8 (.CI(n31917), .I0(n2004), .I1(n2027), .CO(n31918));
    SB_LUT4 mod_5_add_2009_13_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n31709), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_7 (.CI(n31139), .I0(n1205), .I1(n1235), .CO(n31140));
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n31138), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_6 (.CI(n31138), .I0(n1206), .I1(n1235), .CO(n31139));
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n31137), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_5 (.CI(n31137), .I0(n1207), .I1(n1235), .CO(n31138));
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n31136), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_4 (.CI(n31136), .I0(n1208), .I1(n1235), .CO(n31137));
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n40634), 
            .I3(n31135), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_3 (.CI(n31135), .I0(n1209), .I1(n40634), .CO(n31136));
    SB_CARRY mod_5_add_2009_13 (.CI(n31709), .I0(n2899), .I1(n2918), .CO(n31710));
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n40634), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n40634), 
            .CO(n31135));
    SB_LUT4 timer_1508_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1508_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1406_7_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n31916), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_4_lut_adj_1613 (.I0(n111), .I1(n35558), .I2(one_wire_N_520[2]), 
            .I3(one_wire_N_520[3]), .O(n116));
    defparam i1_4_lut_adj_1613.LUT_INIT = 16'haeee;
    SB_LUT4 mod_5_add_2009_12_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n31708), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_12 (.CI(n31708), .I0(n2900), .I1(n2918), .CO(n31709));
    SB_CARRY timer_1508_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n31606));
    SB_CARRY mod_5_add_1406_7 (.CI(n31916), .I0(n2005), .I1(n2027), .CO(n31917));
    SB_LUT4 mod_5_add_1406_6_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n31915), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_11_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n31707), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n31605), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_11 (.CI(n31707), .I0(n2901), .I1(n2918), .CO(n31708));
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n31604), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_27 (.CI(n31604), .I0(n2985), .I1(n3017), .CO(n31605));
    SB_LUT4 add_21_19_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(n30664), .O(n255[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_19 (.CI(n30664), .I0(bit_ctr[17]), .I1(GND_net), .CO(n30665));
    SB_LUT4 add_21_18_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(n30663), .O(n255[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i28310_3_lut (.I0(n20697), .I1(one_wire_N_520[8]), .I2(start), 
            .I3(GND_net), .O(n38337));
    defparam i28310_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 bit_ctr_0__bdd_4_lut_30683 (.I0(bit_ctr[0]), .I1(neopxl_color[18]), 
            .I2(neopxl_color[19]), .I3(bit_ctr[1]), .O(n40720));
    defparam bit_ctr_0__bdd_4_lut_30683.LUT_INIT = 16'he4aa;
    SB_CARRY mod_5_add_1406_6 (.CI(n31915), .I0(n2006), .I1(n2027), .CO(n31916));
    SB_LUT4 mod_5_add_1406_5_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n31914), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n30648));
    SB_CARRY mod_5_add_1406_5 (.CI(n31914), .I0(n2007), .I1(n2027), .CO(n31915));
    SB_LUT4 mod_5_add_1406_4_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n31913), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESS state_i0 (.Q(state[0]), .C(clk32MHz), .E(n21969), .D(state_3__N_369[0]), 
            .S(n36364));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1406_4 (.CI(n31913), .I0(n2008), .I1(n2027), .CO(n31914));
    SB_LUT4 mod_5_add_1406_3_lut (.I0(n2009), .I1(n2009), .I2(n40633), 
            .I3(n31912), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 n40720_bdd_4_lut (.I0(n40720), .I1(neopxl_color[17]), .I2(neopxl_color[16]), 
            .I3(bit_ctr[1]), .O(n40723));
    defparam n40720_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9_4_lut_adj_1614 (.I0(n38337), .I1(one_wire_N_520[10]), .I2(n9_adj_4732), 
            .I3(n116), .O(n20_adj_4820));
    defparam i9_4_lut_adj_1614.LUT_INIT = 16'h0100;
    SB_CARRY mod_5_add_1406_3 (.CI(n31912), .I0(n2009), .I1(n40633), .CO(n31913));
    SB_LUT4 mod_5_add_2009_10_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n31706), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n31603), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_10 (.CI(n31706), .I0(n2902), .I1(n2918), .CO(n31707));
    SB_CARRY mod_5_add_2076_26 (.CI(n31603), .I0(n2986), .I1(n3017), .CO(n31604));
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n31602), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(clk32MHz), .E(n21935), 
            .D(n255[31]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1301), .I1(n1301), .I2(n1334), 
            .I3(n31097), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_10_lut (.I0(n1302), .I1(n1302), .I2(n1334), 
            .I3(n31096), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_10 (.CI(n31096), .I0(n1302), .I1(n1334), .CO(n31097));
    SB_LUT4 mod_5_add_2009_9_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n31705), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_25 (.CI(n31602), .I0(n2987), .I1(n3017), .CO(n31603));
    SB_LUT4 mod_5_add_937_9_lut (.I0(n1303), .I1(n1303), .I2(n1334), .I3(n31095), 
            .O(n1402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_9 (.CI(n31095), .I0(n1303), .I1(n1334), .CO(n31096));
    SB_LUT4 mod_5_add_937_8_lut (.I0(n1304), .I1(n1304), .I2(n1334), .I3(n31094), 
            .O(n1403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n31601), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_8 (.CI(n31094), .I0(n1304), .I1(n1334), .CO(n31095));
    SB_LUT4 mod_5_add_937_7_lut (.I0(n1305), .I1(n1305), .I2(n1334), .I3(n31093), 
            .O(n1404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_7 (.CI(n31093), .I0(n1305), .I1(n1334), .CO(n31094));
    SB_LUT4 mod_5_add_937_6_lut (.I0(n1306), .I1(n1306), .I2(n1334), .I3(n31092), 
            .O(n1405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_6 (.CI(n31092), .I0(n1306), .I1(n1334), .CO(n31093));
    SB_LUT4 mod_5_add_937_5_lut (.I0(n1307), .I1(n1307), .I2(n1334), .I3(n31091), 
            .O(n1406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk32MHz), .E(VCC_net), .D(n22326));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF timer_1508__i1 (.Q(timer[1]), .C(clk32MHz), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 i2_3_lut_4_lut (.I0(n14), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[1] ), .O(n36538));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_CARRY mod_5_add_937_5 (.CI(n31091), .I0(n1307), .I1(n1334), .CO(n31092));
    SB_CARRY mod_5_add_2076_24 (.CI(n31601), .I0(n2988), .I1(n3017), .CO(n31602));
    SB_LUT4 mod_5_add_937_4_lut (.I0(n1308), .I1(n1308), .I2(n1334), .I3(n31090), 
            .O(n1407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_4 (.CI(n31090), .I0(n1308), .I1(n1334), .CO(n31091));
    SB_LUT4 mod_5_add_937_3_lut (.I0(n1309), .I1(n1309), .I2(n40635), 
            .I3(n31089), .O(n1408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_3 (.CI(n31089), .I0(n1309), .I1(n40635), .CO(n31090));
    SB_LUT4 mod_5_add_937_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[22]), .I2(n40635), 
            .I3(VCC_net), .O(n1409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(n40635), 
            .CO(n31089));
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(clk32MHz), .E(n36536), .D(\neo_pixel_transmitter.done_N_583 ), 
            .R(n36830));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_7 (.CI(n30652), .I0(bit_ctr[5]), .I1(GND_net), .CO(n30653));
    SB_DFF timer_1508__i2 (.Q(timer[2]), .C(clk32MHz), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY mod_5_add_2009_9 (.CI(n31705), .I0(n2903), .I1(n2918), .CO(n31706));
    SB_LUT4 mod_5_add_1406_2_lut (.I0(bit_ctr[15]), .I1(bit_ctr[15]), .I2(n40633), 
            .I3(VCC_net), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(n40633), 
            .CO(n31912));
    SB_LUT4 mod_5_add_2009_8_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n31704), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n31600), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i19454_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n27860));
    defparam i19454_2_lut.LUT_INIT = 16'h8888;
    SB_DFF timer_1508__i3 (.Q(timer[3]), .C(clk32MHz), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i4 (.Q(timer[4]), .C(clk32MHz), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i5 (.Q(timer[5]), .C(clk32MHz), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i6 (.Q(timer[6]), .C(clk32MHz), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i7 (.Q(timer[7]), .C(clk32MHz), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i8 (.Q(timer[8]), .C(clk32MHz), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i9 (.Q(timer[9]), .C(clk32MHz), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i10 (.Q(timer[10]), .C(clk32MHz), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i11 (.Q(timer[11]), .C(clk32MHz), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i12 (.Q(timer[12]), .C(clk32MHz), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i13 (.Q(timer[13]), .C(clk32MHz), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i14 (.Q(timer[14]), .C(clk32MHz), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i15 (.Q(timer[15]), .C(clk32MHz), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i16 (.Q(timer[16]), .C(clk32MHz), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i17 (.Q(timer[17]), .C(clk32MHz), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i18 (.Q(timer[18]), .C(clk32MHz), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i19 (.Q(timer[19]), .C(clk32MHz), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i20 (.Q(timer[20]), .C(clk32MHz), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i21 (.Q(timer[21]), .C(clk32MHz), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i22 (.Q(timer[22]), .C(clk32MHz), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i23 (.Q(timer[23]), .C(clk32MHz), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i24 (.Q(timer[24]), .C(clk32MHz), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i25 (.Q(timer[25]), .C(clk32MHz), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i26 (.Q(timer[26]), .C(clk32MHz), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i27 (.Q(timer[27]), .C(clk32MHz), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i28 (.Q(timer[28]), .C(clk32MHz), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i29 (.Q(timer[29]), .C(clk32MHz), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i30 (.Q(timer[30]), .C(clk32MHz), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1508__i31 (.Q(timer[31]), .C(clk32MHz), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 i5_4_lut (.I0(n1105), .I1(n1103), .I2(n27860), .I3(n1108), 
            .O(n12_adj_4821));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF start_103 (.Q(start), .C(clk32MHz), .D(n34460));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n31911), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_18_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n31910), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_18 (.CI(n31910), .I0(n2094), .I1(n2126), .CO(n31911));
    SB_LUT4 i6_4_lut_adj_1615 (.I0(n1107), .I1(n12_adj_4821), .I2(n1106), 
            .I3(n1104), .O(n1136));
    defparam i6_4_lut_adj_1615.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2009_8 (.CI(n31704), .I0(n2904), .I1(n2918), .CO(n31705));
    SB_CARRY mod_5_add_2076_23 (.CI(n31600), .I0(n2989), .I1(n3017), .CO(n31601));
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2009_7_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n31703), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n31599), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i30599_1_lut (.I0(n1433), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40626));
    defparam i30599_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_18 (.CI(n30663), .I0(bit_ctr[16]), .I1(GND_net), .CO(n30664));
    SB_CARRY mod_5_add_2076_22 (.CI(n31599), .I0(n2990), .I1(n3017), .CO(n31600));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n31909), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_7 (.CI(n31703), .I0(n2905), .I1(n2918), .CO(n31704));
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n31598), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_17 (.CI(n31909), .I0(n2095), .I1(n2126), .CO(n31910));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n31702), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_21 (.CI(n31598), .I0(n2991), .I1(n3017), .CO(n31599));
    SB_CARRY mod_5_add_2009_6 (.CI(n31702), .I0(n2906), .I1(n2918), .CO(n31703));
    SB_LUT4 mod_5_add_1473_16_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n31908), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_16 (.CI(n31908), .I0(n2096), .I1(n2126), .CO(n31909));
    SB_LUT4 mod_5_add_1473_15_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n31907), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n31597), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_15 (.CI(n31907), .I0(n2097), .I1(n2126), .CO(n31908));
    SB_LUT4 mod_5_add_2009_5_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n31701), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_20 (.CI(n31597), .I0(n2992), .I1(n3017), .CO(n31598));
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n31596), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_14_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n31906), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_5 (.CI(n31701), .I0(n2907), .I1(n2918), .CO(n31702));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n31700), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_17_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(n30662), .O(n255[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_4 (.CI(n31700), .I0(n2908), .I1(n2918), .CO(n31701));
    SB_LUT4 mod_5_add_2009_3_lut (.I0(n2909), .I1(n2909), .I2(n40625), 
            .I3(n31699), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_19 (.CI(n31596), .I0(n2993), .I1(n3017), .CO(n31597));
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_17 (.CI(n30662), .I0(bit_ctr[15]), .I1(GND_net), .CO(n30663));
    SB_LUT4 i19496_2_lut (.I0(bit_ctr[21]), .I1(n1409), .I2(GND_net), 
            .I3(GND_net), .O(n27902));
    defparam i19496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_1616 (.I0(n1405), .I1(n27902), .I2(n1403), .I3(n1406), 
            .O(n16_adj_4822));
    defparam i6_4_lut_adj_1616.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1473_14 (.CI(n31906), .I0(n2098), .I1(n2126), .CO(n31907));
    SB_LUT4 mod_5_add_1473_13_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n31905), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_3 (.CI(n31699), .I0(n2909), .I1(n40625), .CO(n31700));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n31595), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7_4_lut_adj_1617 (.I0(n1402), .I1(n1404), .I2(n1400), .I3(n1407), 
            .O(n17_adj_4823));
    defparam i7_4_lut_adj_1617.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_16_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(n30661), .O(n255[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9_4_lut_adj_1618 (.I0(n17_adj_4823), .I1(n1408), .I2(n16_adj_4822), 
            .I3(n1401), .O(n1433));
    defparam i9_4_lut_adj_1618.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2009_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[6]), .I2(n40625), 
            .I3(VCC_net), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_18 (.CI(n31595), .I0(n2994), .I1(n3017), .CO(n31596));
    SB_CARRY add_21_16 (.CI(n30661), .I0(bit_ctr[14]), .I1(GND_net), .CO(n30662));
    SB_LUT4 add_21_15_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(n30660), .O(n255[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(n905), .I2(VCC_net), 
            .I3(n30974), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_13 (.CI(n31905), .I0(n2099), .I1(n2126), .CO(n31906));
    SB_LUT4 mod_5_add_1473_12_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n31904), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_12 (.CI(n31904), .I0(n2100), .I1(n2126), .CO(n31905));
    SB_LUT4 mod_5_add_1473_11_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n31903), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_11 (.CI(n31903), .I0(n2101), .I1(n2126), .CO(n31904));
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(n40625), 
            .CO(n31699));
    SB_LUT4 mod_5_add_1473_10_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n31902), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_10 (.CI(n31902), .I0(n2102), .I1(n2126), .CO(n31903));
    SB_LUT4 mod_5_add_1473_9_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n31901), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_9 (.CI(n31901), .I0(n2103), .I1(n2126), .CO(n31902));
    SB_LUT4 mod_5_add_1473_8_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n31900), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_8 (.CI(n31900), .I0(n2104), .I1(n2126), .CO(n31901));
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n31594), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_7_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n31899), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_7 (.CI(n31899), .I0(n2105), .I1(n2126), .CO(n31900));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n31898), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_6 (.CI(n31898), .I0(n2106), .I1(n2126), .CO(n31899));
    SB_LUT4 mod_5_add_1473_5_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n31897), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_5 (.CI(n31897), .I0(n2107), .I1(n2126), .CO(n31898));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n31896), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_4 (.CI(n31896), .I0(n2108), .I1(n2126), .CO(n31897));
    SB_LUT4 mod_5_add_1473_3_lut (.I0(n2109), .I1(n2109), .I2(n40636), 
            .I3(n31895), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_3 (.CI(n31895), .I0(n2109), .I1(n40636), .CO(n31896));
    SB_CARRY mod_5_add_2076_17 (.CI(n31594), .I0(n2995), .I1(n3017), .CO(n31595));
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n31593), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_16 (.CI(n31593), .I0(n2996), .I1(n3017), .CO(n31594));
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n31592), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_2_lut (.I0(bit_ctr[14]), .I1(bit_ctr[14]), .I2(n40636), 
            .I3(VCC_net), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(n40636), 
            .CO(n31895));
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n31894), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(clk32MHz), .E(n21935), 
            .D(n255[30]), .R(n22215));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1540_19_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n31893), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_15 (.CI(n30660), .I0(bit_ctr[13]), .I1(GND_net), .CO(n30661));
    SB_CARRY mod_5_add_1540_19 (.CI(n31893), .I0(n2193), .I1(n2225), .CO(n31894));
    SB_LUT4 mod_5_add_1540_18_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n31892), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_18 (.CI(n31892), .I0(n2194), .I1(n2225), .CO(n31893));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n31891), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_17 (.CI(n31891), .I0(n2195), .I1(n2225), .CO(n31892));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n31890), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_16 (.CI(n31890), .I0(n2196), .I1(n2225), .CO(n31891));
    SB_LUT4 mod_5_add_1540_15_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n31889), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_15 (.CI(n31889), .I0(n2197), .I1(n2225), .CO(n31890));
    SB_LUT4 mod_5_add_1540_14_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n31888), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_14 (.CI(n31888), .I0(n2198), .I1(n2225), .CO(n31889));
    SB_LUT4 mod_5_add_1540_13_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n31887), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_13 (.CI(n31887), .I0(n2199), .I1(n2225), .CO(n31888));
    SB_LUT4 mod_5_add_1540_12_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n31886), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_12 (.CI(n31886), .I0(n2200), .I1(n2225), .CO(n31887));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n31885), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_11 (.CI(n31885), .I0(n2201), .I1(n2225), .CO(n31886));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n31884), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_10 (.CI(n31884), .I0(n2202), .I1(n2225), .CO(n31885));
    SB_LUT4 mod_5_add_1540_9_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n31883), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1540_9 (.CI(n31883), .I0(n2203), .I1(n2225), .CO(n31884));
    SB_LUT4 mod_5_add_1540_8_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n31882), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_8 (.CI(n31882), .I0(n2204), .I1(n2225), .CO(n31883));
    SB_LUT4 mod_5_add_1540_7_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n31881), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_7 (.CI(n31881), .I0(n2205), .I1(n2225), .CO(n31882));
    SB_LUT4 mod_5_add_1540_6_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n31880), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_6 (.CI(n31880), .I0(n2206), .I1(n2225), .CO(n31881));
    SB_LUT4 mod_5_add_1540_5_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n31879), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_5 (.CI(n31879), .I0(n2207), .I1(n2225), .CO(n31880));
    SB_LUT4 mod_5_add_1540_4_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n31878), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_4 (.CI(n31878), .I0(n2208), .I1(n2225), .CO(n31879));
    SB_LUT4 mod_5_add_1540_3_lut (.I0(n2209), .I1(n2209), .I2(n40637), 
            .I3(n31877), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_3 (.CI(n31877), .I0(n2209), .I1(n40637), .CO(n31878));
    SB_LUT4 mod_5_add_1540_2_lut (.I0(bit_ctr[13]), .I1(bit_ctr[13]), .I2(n40637), 
            .I3(VCC_net), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(n40637), 
            .CO(n31877));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n31876), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n31875), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_20 (.CI(n31875), .I0(n2292), .I1(n2324), .CO(n31876));
    SB_LUT4 mod_5_add_1607_19_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n31874), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_19 (.CI(n31874), .I0(n2293), .I1(n2324), .CO(n31875));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n31873), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_15 (.CI(n31592), .I0(n2997), .I1(n3017), .CO(n31593));
    SB_CARRY mod_5_add_1607_18 (.CI(n31873), .I0(n2294), .I1(n2324), .CO(n31874));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n31872), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_17 (.CI(n31872), .I0(n2295), .I1(n2324), .CO(n31873));
    SB_LUT4 mod_5_add_1607_16_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n31871), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_16 (.CI(n31871), .I0(n2296), .I1(n2324), .CO(n31872));
    SB_LUT4 mod_5_add_1607_15_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n31870), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_15 (.CI(n31870), .I0(n2297), .I1(n2324), .CO(n31871));
    SB_LUT4 mod_5_add_1607_14_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n31869), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_14 (.CI(n31869), .I0(n2298), .I1(n2324), .CO(n31870));
    SB_LUT4 mod_5_add_1607_13_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n31868), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_13 (.CI(n31868), .I0(n2299), .I1(n2324), .CO(n31869));
    SB_LUT4 mod_5_add_1607_12_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n31867), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_12 (.CI(n31867), .I0(n2300), .I1(n2324), .CO(n31868));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n31866), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_11 (.CI(n31866), .I0(n2301), .I1(n2324), .CO(n31867));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n31865), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_10 (.CI(n31865), .I0(n2302), .I1(n2324), .CO(n31866));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n31864), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_9 (.CI(n31864), .I0(n2303), .I1(n2324), .CO(n31865));
    SB_LUT4 mod_5_add_1607_8_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n31863), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_8 (.CI(n31863), .I0(n2304), .I1(n2324), .CO(n31864));
    SB_LUT4 mod_5_add_1607_7_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n31862), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_7 (.CI(n31862), .I0(n2305), .I1(n2324), .CO(n31863));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n31861), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_6 (.CI(n31861), .I0(n2306), .I1(n2324), .CO(n31862));
    SB_LUT4 mod_5_add_1607_5_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n31860), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_5 (.CI(n31860), .I0(n2307), .I1(n2324), .CO(n31861));
    SB_LUT4 mod_5_add_1607_4_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n31859), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_4 (.CI(n31859), .I0(n2308), .I1(n2324), .CO(n31860));
    SB_LUT4 mod_5_add_1607_3_lut (.I0(n2309), .I1(n2309), .I2(n40638), 
            .I3(n31858), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_3 (.CI(n31858), .I0(n2309), .I1(n40638), .CO(n31859));
    SB_LUT4 mod_5_add_1607_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[12]), .I2(n40638), 
            .I3(VCC_net), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(n40638), 
            .CO(n31858));
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n31857), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n31856), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_21 (.CI(n31856), .I0(n2391), .I1(n2423), .CO(n31857));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n31855), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_20 (.CI(n31855), .I0(n2392), .I1(n2423), .CO(n31856));
    SB_LUT4 mod_5_add_1674_19_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n31854), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_19 (.CI(n31854), .I0(n2393), .I1(n2423), .CO(n31855));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n31853), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_18 (.CI(n31853), .I0(n2394), .I1(n2423), .CO(n31854));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n31852), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_17 (.CI(n31852), .I0(n2395), .I1(n2423), .CO(n31853));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n31851), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_16 (.CI(n31851), .I0(n2396), .I1(n2423), .CO(n31852));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n31850), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_15 (.CI(n31850), .I0(n2397), .I1(n2423), .CO(n31851));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n31849), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_14 (.CI(n31849), .I0(n2398), .I1(n2423), .CO(n31850));
    SB_LUT4 mod_5_add_1674_13_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n31848), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_13 (.CI(n31848), .I0(n2399), .I1(n2423), .CO(n31849));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n31847), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_12 (.CI(n31847), .I0(n2400), .I1(n2423), .CO(n31848));
    SB_LUT4 mod_5_add_1674_11_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n31846), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_11 (.CI(n31846), .I0(n2401), .I1(n2423), .CO(n31847));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n31845), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_10 (.CI(n31845), .I0(n2402), .I1(n2423), .CO(n31846));
    SB_LUT4 mod_5_add_1674_9_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n31844), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_9 (.CI(n31844), .I0(n2403), .I1(n2423), .CO(n31845));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n31843), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_8 (.CI(n31843), .I0(n2404), .I1(n2423), .CO(n31844));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n31842), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_7 (.CI(n31842), .I0(n2405), .I1(n2423), .CO(n31843));
    SB_LUT4 mod_5_add_1674_6_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n31841), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_6 (.CI(n31841), .I0(n2406), .I1(n2423), .CO(n31842));
    SB_LUT4 mod_5_add_1674_5_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n31840), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_5 (.CI(n31840), .I0(n2407), .I1(n2423), .CO(n31841));
    SB_LUT4 mod_5_add_1674_4_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n31839), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_4 (.CI(n31839), .I0(n2408), .I1(n2423), .CO(n31840));
    SB_LUT4 mod_5_add_1674_3_lut (.I0(n2409), .I1(n2409), .I2(n40639), 
            .I3(n31838), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_3 (.CI(n31838), .I0(n2409), .I1(n40639), .CO(n31839));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(bit_ctr[11]), .I1(bit_ctr[11]), .I2(n40639), 
            .I3(VCC_net), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(n40639), 
            .CO(n31838));
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n31837), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n31836), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_22 (.CI(n31836), .I0(n2490), .I1(n2522), .CO(n31837));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n31835), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_21 (.CI(n31835), .I0(n2491), .I1(n2522), .CO(n31836));
    SB_LUT4 mod_5_add_1741_20_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n31834), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_20 (.CI(n31834), .I0(n2492), .I1(n2522), .CO(n31835));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n31833), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_19 (.CI(n31833), .I0(n2493), .I1(n2522), .CO(n31834));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n31832), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_18 (.CI(n31832), .I0(n2494), .I1(n2522), .CO(n31833));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n31831), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_17 (.CI(n31831), .I0(n2495), .I1(n2522), .CO(n31832));
    SB_LUT4 add_21_14_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(n30659), .O(n255[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_16_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n31830), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n30973), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_16 (.CI(n31830), .I0(n2496), .I1(n2522), .CO(n31831));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n31829), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_15 (.CI(n31829), .I0(n2497), .I1(n2522), .CO(n31830));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n31828), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_14 (.CI(n31828), .I0(n2498), .I1(n2522), .CO(n31829));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n31827), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_13 (.CI(n31827), .I0(n2499), .I1(n2522), .CO(n31828));
    SB_LUT4 mod_5_add_1741_12_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n31826), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_12 (.CI(n31826), .I0(n2500), .I1(n2522), .CO(n31827));
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n31591), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_11_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n31825), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_11 (.CI(n31825), .I0(n2501), .I1(n2522), .CO(n31826));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n31824), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_10 (.CI(n31824), .I0(n2502), .I1(n2522), .CO(n31825));
    SB_LUT4 mod_5_add_1741_9_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n31823), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_669_6 (.CI(n30973), .I0(n906), .I1(VCC_net), .CO(n30974));
    SB_CARRY mod_5_add_1741_9 (.CI(n31823), .I0(n2503), .I1(n2522), .CO(n31824));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n31822), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_8 (.CI(n31822), .I0(n2504), .I1(n2522), .CO(n31823));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n31821), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_7 (.CI(n31821), .I0(n2505), .I1(n2522), .CO(n31822));
    SB_CARRY mod_5_add_2076_14 (.CI(n31591), .I0(n2998), .I1(n3017), .CO(n31592));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n31820), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_6 (.CI(n31820), .I0(n2506), .I1(n2522), .CO(n31821));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n31819), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_5 (.CI(n31819), .I0(n2507), .I1(n2522), .CO(n31820));
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n36488), .I2(VCC_net), 
            .I3(n30972), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_4_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n31818), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_6_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(n30651), .O(n255[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_4 (.CI(n31818), .I0(n2508), .I1(n2522), .CO(n31819));
    SB_CARRY mod_5_add_669_5 (.CI(n30972), .I0(n36488), .I1(VCC_net), 
            .CO(n30973));
    SB_LUT4 mod_5_add_1741_3_lut (.I0(n2509), .I1(n2509), .I2(n40640), 
            .I3(n31817), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n31590), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_3 (.CI(n31817), .I0(n2509), .I1(n40640), .CO(n31818));
    SB_LUT4 mod_5_add_1741_2_lut (.I0(bit_ctr[10]), .I1(bit_ctr[10]), .I2(n40640), 
            .I3(VCC_net), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(n40640), 
            .CO(n31817));
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n22070), .I2(VCC_net), 
            .I3(n30971), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_13 (.CI(n31590), .I0(n2999), .I1(n3017), .CO(n31591));
    SB_LUT4 i2_2_lut_adj_1619 (.I0(one_wire_N_520[5]), .I1(one_wire_N_520[7]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4824));
    defparam i2_2_lut_adj_1619.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_669_4 (.CI(n30971), .I0(n22070), .I1(VCC_net), 
            .CO(n30972));
    SB_CARRY add_21_14 (.CI(n30659), .I0(bit_ctr[12]), .I1(GND_net), .CO(n30660));
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n19296), .I2(GND_net), 
            .I3(n30970), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk32MHz), .D(n22291));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n31589), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i4_4_lut_adj_1620 (.I0(n7_adj_4824), .I1(\state[1] ), .I2(one_wire_N_520[11]), 
            .I3(n20_adj_4820), .O(n40929));
    defparam i4_4_lut_adj_1620.LUT_INIT = 16'hfeff;
    SB_CARRY mod_5_add_2076_12 (.CI(n31589), .I0(n3000), .I1(n3017), .CO(n31590));
    SB_LUT4 bit_ctr_0__bdd_4_lut_30678 (.I0(bit_ctr[0]), .I1(neopxl_color[6]), 
            .I2(neopxl_color[7]), .I3(bit_ctr[1]), .O(n40702));
    defparam bit_ctr_0__bdd_4_lut_30678.LUT_INIT = 16'he4aa;
    SB_CARRY add_21_6 (.CI(n30651), .I0(bit_ctr[4]), .I1(GND_net), .CO(n30652));
    SB_CARRY mod_5_add_669_3 (.CI(n30970), .I0(n19296), .I1(GND_net), 
            .CO(n30971));
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n31588), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 n40702_bdd_4_lut (.I0(n40702), .I1(neopxl_color[5]), .I2(neopxl_color[4]), 
            .I3(bit_ctr[1]), .O(n39869));
    defparam n40702_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut_adj_1621 (.I0(bit_ctr[22]), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(GND_net), .O(n30_adj_4825));
    defparam i2_2_lut_adj_1621.LUT_INIT = 16'heeee;
    SB_LUT4 i20_4_lut_adj_1622 (.I0(bit_ctr[20]), .I1(bit_ctr[7]), .I2(bit_ctr[16]), 
            .I3(bit_ctr[30]), .O(n48_adj_4826));
    defparam i20_4_lut_adj_1622.LUT_INIT = 16'hfffe;
    SB_LUT4 i30613_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40640));
    defparam i30613_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i18_4_lut_adj_1623 (.I0(bit_ctr[25]), .I1(bit_ctr[10]), .I2(bit_ctr[9]), 
            .I3(bit_ctr[27]), .O(n46_adj_4827));
    defparam i18_4_lut_adj_1623.LUT_INIT = 16'hfffe;
    SB_LUT4 i29359_3_lut_4_lut (.I0(n32422), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(n20592), .O(n39270));
    defparam i29359_3_lut_4_lut.LUT_INIT = 16'hcfdf;
    SB_LUT4 i3_2_lut_adj_1624 (.I0(n2491), .I1(n2504), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_4828));
    defparam i3_2_lut_adj_1624.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_1625 (.I0(n2496), .I1(n2505), .I2(n2500), .I3(n2499), 
            .O(n34_adj_4829));
    defparam i13_4_lut_adj_1625.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1626 (.I0(bit_ctr[10]), .I1(n2497), .I2(n2509), 
            .I3(GND_net), .O(n22_adj_4830));
    defparam i1_3_lut_adj_1626.LUT_INIT = 16'hecec;
    SB_LUT4 i19_4_lut_adj_1627 (.I0(bit_ctr[15]), .I1(bit_ctr[29]), .I2(bit_ctr[12]), 
            .I3(bit_ctr[23]), .O(n47_adj_4831));
    defparam i19_4_lut_adj_1627.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1628 (.I0(n2490), .I1(n34_adj_4829), .I2(n24_adj_4828), 
            .I3(n2494), .O(n38_adj_4832));
    defparam i17_4_lut_adj_1628.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1629 (.I0(n2501), .I1(n2502), .I2(n2506), .I3(n2492), 
            .O(n36_adj_4833));
    defparam i15_4_lut_adj_1629.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1630 (.I0(n2495), .I1(n2498), .I2(n2493), .I3(n22_adj_4830), 
            .O(n37_adj_4834));
    defparam i16_4_lut_adj_1630.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1631 (.I0(n2507), .I1(n2508), .I2(n2503), .I3(n2489), 
            .O(n35_adj_4835));
    defparam i14_4_lut_adj_1631.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1632 (.I0(bit_ctr[19]), .I1(bit_ctr[21]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[14]), .O(n45_adj_4836));
    defparam i17_4_lut_adj_1632.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1633 (.I0(bit_ctr[11]), .I1(bit_ctr[5]), .I2(bit_ctr[28]), 
            .I3(bit_ctr[6]), .O(n44_adj_4837));
    defparam i16_4_lut_adj_1633.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1634 (.I0(n35_adj_4835), .I1(n37_adj_4834), .I2(n36_adj_4833), 
            .I3(n38_adj_4832), .O(n2522));
    defparam i20_4_lut_adj_1634.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15_4_lut_adj_1635 (.I0(n2897), .I1(n2886), .I2(n2908), .I3(n2890), 
            .O(n40_adj_4838));
    defparam i15_4_lut_adj_1635.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1636 (.I0(n2903), .I1(bit_ctr[6]), .I2(n2909), 
            .I3(GND_net), .O(n27_adj_4839));
    defparam i2_3_lut_adj_1636.LUT_INIT = 16'heaea;
    SB_LUT4 i13_3_lut_adj_1637 (.I0(n2895), .I1(n2888), .I2(n2901), .I3(GND_net), 
            .O(n38_adj_4840));
    defparam i13_3_lut_adj_1637.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut_adj_1638 (.I0(n2900), .I1(n2891), .I2(n2899), .I3(n2902), 
            .O(n43_adj_4841));
    defparam i18_4_lut_adj_1638.LUT_INIT = 16'hfffe;
    SB_LUT4 i30612_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40639));
    defparam i30612_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17_4_lut_adj_1639 (.I0(n2885), .I1(n2904), .I2(n2906), .I3(n2887), 
            .O(n42_adj_4842));
    defparam i17_4_lut_adj_1639.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1640 (.I0(n2892), .I1(n2894), .I2(n2907), .I3(n2896), 
            .O(n41_adj_4843));
    defparam i16_4_lut_adj_1640.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1641 (.I0(bit_ctr[3]), .I1(n30_adj_4825), .I2(bit_ctr[13]), 
            .I3(bit_ctr[4]), .O(n43_adj_4844));
    defparam i15_4_lut_adj_1641.LUT_INIT = 16'hfefc;
    SB_LUT4 i20_4_lut_adj_1642 (.I0(n27_adj_4839), .I1(n40_adj_4838), .I2(n2898), 
            .I3(n2889), .O(n45_adj_4845));
    defparam i20_4_lut_adj_1642.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1643 (.I0(n43_adj_4841), .I1(n2905), .I2(n38_adj_4840), 
            .I3(n2893), .O(n47_adj_4846));
    defparam i22_4_lut_adj_1643.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut_adj_1644 (.I0(n47_adj_4846), .I1(n45_adj_4845), .I2(n41_adj_4843), 
            .I3(n42_adj_4842), .O(n2918));
    defparam i24_4_lut_adj_1644.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1645 (.I0(n45_adj_4836), .I1(n47_adj_4831), .I2(n46_adj_4827), 
            .I3(n48_adj_4826), .O(n54_adj_4847));
    defparam i26_4_lut_adj_1645.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1646 (.I0(bit_ctr[24]), .I1(bit_ctr[8]), .I2(bit_ctr[18]), 
            .I3(bit_ctr[26]), .O(n49_adj_4848));
    defparam i21_4_lut_adj_1646.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut_adj_1647 (.I0(n49_adj_4848), .I1(n54_adj_4847), .I2(n43_adj_4844), 
            .I3(n44_adj_4837), .O(\state_3__N_369[1] ));
    defparam i27_4_lut_adj_1647.LUT_INIT = 16'hfffe;
    SB_LUT4 bit_ctr_2__bdd_4_lut (.I0(bit_ctr[2]), .I1(n38446), .I2(n38449), 
            .I3(n41597), .O(n40654));
    defparam bit_ctr_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n40654_bdd_4_lut (.I0(n40654), .I1(n39869), .I2(n38455), .I3(n41597), 
            .O(n40657));
    defparam n40654_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1648 (.I0(one_wire_N_520[3]), .I1(one_wire_N_520[4]), 
            .I2(one_wire_N_520[2]), .I3(GND_net), .O(n32422));
    defparam i2_3_lut_adj_1648.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut (.I0(n14), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n36326));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 i29268_2_lut_3_lut (.I0(n28022), .I1(\neo_pixel_transmitter.done ), 
            .I2(state[0]), .I3(GND_net), .O(n39203));   // verilog/neopixel.v(35[12] 117[6])
    defparam i29268_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1649 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n20719));   // verilog/neopixel.v(52[18] 72[12])
    defparam i1_2_lut_adj_1649.LUT_INIT = 16'hbbbb;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut_adj_1650 (.I0(state[0]), .I1(\state[1] ), .I2(LED_c), 
            .I3(\state_3__N_369[1] ), .O(n22215));   // verilog/neopixel.v(35[12] 117[6])
    defparam i2_3_lut_4_lut_adj_1650.LUT_INIT = 16'h8000;
    SB_LUT4 i29552_3_lut_4_lut (.I0(\state[1] ), .I1(n39580), .I2(start), 
            .I3(n20592), .O(n39581));
    defparam i29552_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_3_lut_adj_1651 (.I0(bit_ctr[11]), .I1(n2403), .I2(n2409), 
            .I3(GND_net), .O(n27_adj_4849));
    defparam i7_3_lut_adj_1651.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut_adj_1652 (.I0(n2390), .I1(n2391), .I2(n2397), .I3(n2394), 
            .O(n33_adj_4850));
    defparam i13_4_lut_adj_1652.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1653 (.I0(n2392), .I1(n2405), .I2(n2400), .I3(n2398), 
            .O(n32_adj_4851));
    defparam i12_4_lut_adj_1653.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1654 (.I0(n2396), .I1(n2402), .I2(n2408), .I3(n2399), 
            .O(n31_adj_4852));
    defparam i11_4_lut_adj_1654.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1655 (.I0(n2393), .I1(n2406), .I2(n2395), .I3(n2407), 
            .O(n35_adj_4853));
    defparam i15_4_lut_adj_1655.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1656 (.I0(n33_adj_4850), .I1(n27_adj_4849), .I2(n2404), 
            .I3(n2401), .O(n37_adj_4854));
    defparam i17_4_lut_adj_1656.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1657 (.I0(n37_adj_4854), .I1(n35_adj_4853), .I2(n31_adj_4852), 
            .I3(n32_adj_4851), .O(n2423));
    defparam i19_4_lut_adj_1657.LUT_INIT = 16'hfffe;
    SB_LUT4 i30611_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40638));
    defparam i30611_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29549_3_lut_4_lut (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(n28022), .I3(start), .O(n39196));
    defparam i29549_3_lut_4_lut.LUT_INIT = 16'hff10;
    SB_LUT4 i2_3_lut_4_lut_adj_1658 (.I0(state[0]), .I1(\neo_pixel_transmitter.done ), 
            .I2(n28022), .I3(\state[1] ), .O(n36830));
    defparam i2_3_lut_4_lut_adj_1658.LUT_INIT = 16'h0100;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5024_2_lut_3_lut (.I0(bit_ctr[28]), .I1(n36524), .I2(bit_ctr[27]), 
            .I3(GND_net), .O(n9244));   // verilog/neopixel.v(22[26:36])
    defparam i5024_2_lut_3_lut.LUT_INIT = 16'h6060;
    SB_LUT4 i19445_2_lut_3_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(bit_ctr[29]), 
            .I3(GND_net), .O(n27850));
    defparam i19445_2_lut_3_lut.LUT_INIT = 16'h6464;
    SB_LUT4 i29429_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n36524), .I2(bit_ctr[27]), 
            .I3(n838), .O(n22070));
    defparam i29429_3_lut_4_lut.LUT_INIT = 16'h6696;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, \Ki[9] , \Ki[10] , \Ki[11] , \Kp[14] , 
            PWMLimit, \Kp[15] , \Ki[12] , \Kp[9] , \Kp[10] , \Ki[2] , 
            \Ki[13] , \Ki[14] , \Ki[15] , \Kp[7] , \Ki[1] , \Ki[0] , 
            \Kp[11] , \Ki[3] , \Ki[4] , \Ki[5] , \Ki[6] , \Ki[7] , 
            \Ki[8] , \Kp[1] , \Kp[0] , \Kp[2] , \Kp[12] , \Kp[3] , 
            \Kp[13] , \Kp[8] , \Kp[4] , \Kp[5] , IntegralLimit, \Kp[6] , 
            duty, clk32MHz, VCC_net, setpoint, motor_state, n40620) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input \Ki[9] ;
    input \Ki[10] ;
    input \Ki[11] ;
    input \Kp[14] ;
    input [23:0]PWMLimit;
    input \Kp[15] ;
    input \Ki[12] ;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Ki[2] ;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[15] ;
    input \Kp[7] ;
    input \Ki[1] ;
    input \Ki[0] ;
    input \Kp[11] ;
    input \Ki[3] ;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Kp[2] ;
    input \Kp[12] ;
    input \Kp[3] ;
    input \Kp[13] ;
    input \Kp[8] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input [23:0]IntegralLimit;
    input \Kp[6] ;
    output [23:0]duty;
    input clk32MHz;
    input VCC_net;
    input [23:0]setpoint;
    input [23:0]motor_state;
    output n40620;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n31507;
    wire [21:0]n9589;
    
    wire n658, n31508;
    wire [47:0]n106;
    
    wire n585, n31506;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3513 ;
    
    wire n679, n11;
    wire [23:0]n1;
    
    wire n30904;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(23[23:31])
    
    wire n752, n825, n512, n31505;
    wire [23:0]n28;
    
    wire n1023;
    wire [23:0]n1_adj_4704;
    
    wire \PID_CONTROLLER.integral_23__N_3561 ;
    wire [23:0]n3141;
    
    wire n1096, n439, n31504, n31033;
    wire [13:0]n12717;
    
    wire n463, n31034, n30905, n366, n31503, n898, n685, n758;
    wire [3:0]n9993;
    
    wire n30518;
    wire [4:0]n9986;
    
    wire n971, n1044, n1117, n533, n98, n29, n831, n171, n244, 
        n317, n390, n463_adj_4283, n536, n609, n107, n38, n682, 
        n755, n828, n180, n901, n974, n1047, n1120, n101, n32, 
        n174, n247, n320, n393, n904, n466, n539, n253, n612, 
        n685_adj_4288, n758_adj_4289, n831_adj_4290, n904_adj_4292, 
        n977, n977_adj_4293, n1050, n104, n35, n606, n177, n250, 
        n326, n323, n1050_adj_4295, n396, n469, n542, n399, n615, 
        n688, n679_adj_4297, n4, n761;
    wire [23:0]duty_23__N_3613;
    wire [23:0]n257;
    
    wire n256;
    wire [23:0]duty_23__N_3588;
    
    wire n293, n31502, duty_23__N_3612;
    wire [23:0]duty_23__N_3489;
    
    wire n834, n220, n31501, n147_adj_4298, n31500, n5, n74, n907, 
        n980;
    wire [20:0]n10450;
    
    wire n31499, n107_adj_4299, n38_adj_4300, n180_adj_4301, n253_adj_4302, 
        n326_adj_4303, n399_adj_4304, n472, n545, n618, n752_adj_4305, 
        n691, n825_adj_4306, n764, n837, n910, n31498, n110, n41, 
        n183, n256_adj_4307, n329, n402, n475, n898_adj_4308, n971_adj_4309, 
        n1044_adj_4310, n125, n56, n1117_adj_4311, n92, n23, n165, 
        n238, n311, n384, n457, n198, n548, n530, n603, n676, 
        n621, n749;
    wire [14:0]n12509;
    
    wire n390_adj_4315, n31032, n31497, n694, n767, n840, n9_adj_4316, 
        n30903, n113, n822, n44, n895, n186, n259, n968, n332, 
        n405, n478, n1041, n104_adj_4319, n35_adj_4321, n1114, n551, 
        n624, n116, n697, n47, n189, n262, n122, n335, n408, 
        n53, n481, n770, n116_adj_4322, n47_adj_4323, n189_adj_4324, 
        n262_adj_4325, n335_adj_4326, n408_adj_4327, n89, n20_adj_4329, 
        n162, n472_adj_4330, n481_adj_4331, n554, n627, n700, n235, 
        n308, n31496, n381, n454, n527, n119, n600, n673, n50, 
        n746, n819, n31495, n192, n265, n317_adj_4332, n31031, 
        n338, n411, n484, n892, n31494, n31493, n965, n1099, 
        n31492, n1038, n1111, n86, n17_adj_4334, n159, n232, n305, 
        n378, n451, n524, n597, n670, n743, n816, n889, n962, 
        n1035, n1108, n1026, n31491, n557, n630, n244_adj_4335, 
        n31030, n195, n7_adj_4336, n30902, n5_adj_4338, n30901, 
        n122_adj_4340, n53_adj_4341, n195_adj_4342, n953, n31490, 
        n880, n31489, n807, n31488, n734, n31487, n661, n31486, 
        n588, n31485, n515, n31484, n442, n31483, n369, n31482, 
        n296, n31481, n113_adj_4343, n44_adj_4344, n268, n186_adj_4345, 
        n268_adj_4346, n341, n414, n259_adj_4347, n341_adj_4348, n414_adj_4349, 
        n487, n332_adj_4350, n405_adj_4351, n478_adj_4352, n551_adj_4353, 
        n624_adj_4354, n697_adj_4355, n770_adj_4356, n83, n14_adj_4358, 
        n156, n229, n302, n375, n448, n521, n594, n223, n31480, 
        n150_adj_4359, n31479, n8_adj_4360, n77, n667, n740;
    wire [19:0]n10889;
    
    wire n31478, n31477, n813, n31476, n886, n959, n98_adj_4362, 
        n29_adj_4363, n560, n1032, n31475, n1105, n80, n11_adj_4364, 
        n125_adj_4365, n56_adj_4366, n171_adj_4367, n198_adj_4368, n271, 
        n344, n153_adj_4370, n417, n6_adj_4371, n554_adj_4372, n627_adj_4373;
    wire [1:0]n10004;
    
    wire n700_adj_4374, n4_adj_4375;
    wire [2:0]n9999;
    
    wire n490, n271_adj_4376, n12_adj_4377, n8_adj_4378, n11_adj_4379, 
        n6_adj_4380, n30620, n18_adj_4381, n13_adj_4382, n4_adj_4383, 
        n37896, n545_adj_4385, n31474, n487_adj_4388, n31473, n1102, 
        n31472, n1029, n31471, n956, n31470, n883, n31469, n810, 
        n31468, n737, n31467, n664, n31466, n591, n31465, n518, 
        n31464, n445, n31463, n372, n31462, n560_adj_4389, n299, 
        n31461, n226, n31460, n31459, n3, n30900, n31029;
    wire [18:0]n11287;
    
    wire n31458, n17_adj_4391, n9_adj_4392, n11_adj_4393, n39496, 
        n39493, n31457, n41474, n39867, n39746, n41456, n39744, 
        n39742, n31456, n41450, n27, n15_adj_4394, n13_adj_4395, 
        n39436, n21_adj_4396, n19_adj_4397, n17_adj_4398, n39442, 
        n43, n16_adj_4399, n31455, n39419, n8_adj_4400, n45, n24_adj_4401, 
        n39452, n31454, n39715, n39711, n25_adj_4402, n23_adj_4403, 
        n39988, n31, n29_adj_4404, n39835, n37, n35_adj_4405, n33, 
        n40042, n39748;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3564 ;
    
    wire n41443, n39736, n31453, n41437, n12_adj_4406, n31452, n39469, 
        n41461, n10_adj_4407, n31451, n31450, n30, n31449, n31448, 
        n39933, n39481, n41441, n31447, n39859, n41467, n39994, 
        n30899, n31446, n41432, n30898, n40064, n41429, n16_adj_4410, 
        n39454, n31445, n24_adj_4411, n6_adj_4412, n39873, n39874, 
        n31444, n39458, n30897, n31443, n8_adj_4413, n41427, n39851, 
        n31442, n39734, n4_adj_4414, n31441, n39966, n31440, n39967, 
        n344_adj_4415, n12_adj_4416, n39429, n10_adj_4417, n30_adj_4418, 
        n39431, n40048, n417_adj_4419, n6_adj_4420;
    wire [3:0]n13692;
    wire [4:0]n13668;
    
    wire n39908, n40099, n40100, n39, n40083, n6_adj_4421, n39974, 
        n39975, n39421, n39853, n39906, n41_adj_4422, n39423, n40004, 
        n40, n40006, n4_adj_4423, n39990, n39991, n39471, n40046, 
        n39902, n40097, n40098, n40085, n39461, n39998, n40_adj_4424, 
        \PID_CONTROLLER.integral_23__N_3563 , n40000, n177_adj_4425;
    wire [9:0]n13343;
    wire [8:0]n13442;
    
    wire n31439, n31438, n30896, n31437, n31436, n250_adj_4426;
    wire [1:0]n13712;
    
    wire n31435, n30895, n31434, n31433, n31432, n31431, n618_adj_4427;
    wire [17:0]n11646;
    
    wire n31430, n31429;
    wire [0:0]n7896;
    wire [0:0]n7900;
    
    wire n30739, n31428;
    wire [47:0]n155;
    
    wire n30738, n30894, n31427, n31426, n31425, n31424, n4_adj_4428;
    wire [2:0]n13707;
    
    wire n490_adj_4429, n31423, n12_adj_4431, n31422, n691_adj_4432, 
        n30893, n30737, n8_adj_4433, n11_adj_4434, n6_adj_4435, n31421, 
        n30411, n31420, n31419, n18_adj_4437, n13_adj_4438, n4_adj_4439, 
        n37173, n31418, n31417, n31416, n31415, n764_adj_4440, n31414, 
        n30736, n31413;
    wire [16:0]n11968;
    
    wire n31412, n31411, n31410, n31409, n31408, n837_adj_4442, 
        n30892, n30891, n31407, n31406, n31405, n31404, n31403, 
        n31402, n31401, n30890, n31400, n30889, n30888, n31399, 
        n30887, n30735, n30734, n30886, n31398, n31397, n31396, 
        n323_adj_4444;
    wire [11:0]n13080;
    wire [10:0]n13223;
    
    wire n910_adj_4445, n30772, n30885, n30733, n30884, n30771, 
        n30883, n30882, n30881, n30880, n30770, n30732, n30879, 
        n30945, n30731, n30944, n30878, n30769, n30943, n30877, 
        n30730, n30768, n30816, n30729, n30815;
    wire [6:0]n13585;
    wire [5:0]n13633;
    
    wire n31005, n31004, n30942, n396_adj_4451, n30814, n30767, 
        n41_adj_4452, n39_adj_4454, n45_adj_4455, n30941;
    wire [5:0]n9978;
    
    wire n32267, n32266, n32265, n32264, n32263;
    wire [6:0]n9969;
    
    wire n32262, n32261, n32260, n32259, n31003, n31002, n31001, 
        n32258, n32257, n31000;
    wire [7:0]n9959;
    
    wire n32256, n32255, n32254, n32253, n32252, n30940, n32251, 
        n32250;
    wire [8:0]n9948;
    
    wire n32249, n32248, n32247, n32246, n30766, n32245, n32244, 
        n30728, n32243, n32242;
    wire [9:0]n9936;
    
    wire n32241, n32240, n32239, n32238, n30939, n30938, n32237, 
        n32236, n32235, n32234, n32233;
    wire [10:0]n9923;
    
    wire n32232, n32231, n32230, n32229, n32228, n37_adj_4458, n29_adj_4459, 
        n31_adj_4460, n43_adj_4461, n23_adj_4462, n25_adj_4463, n35_adj_4464, 
        n11_adj_4465, n13_adj_4466, n15_adj_4467, n27_adj_4469, n33_adj_4470, 
        n9_adj_4471, n17_adj_4472, n19_adj_4473, n21_adj_4475, n39369, 
        n39361, n12_adj_4476, n10_adj_4477, n30_adj_4478, n32227, 
        n39379, n39650, n39646, n39972, n39803, n40038, n16_adj_4479, 
        n6_adj_4480, n39950, n39951, n8_adj_4481, n24_adj_4482, n39347, 
        n39345, n39857, n39918, n4_adj_4483, n39948, n39949, n39357, 
        n39355, n40052, n39920, n40103, n40104, n40079, n39349, 
        n40016, n40_adj_4484, n40018, n32226, n32225, n32224, n32223;
    wire [11:0]n9909;
    
    wire n32222, n32221, n32220, n32219, n32218, n32217, n32216, 
        n32215, n32214, n39_adj_4485, n32213, n41_adj_4486, n45_adj_4487, 
        n32212, n43_adj_4488, n30813, n37_adj_4489, n29_adj_4490, 
        n31_adj_4491, n23_adj_4492, n25_adj_4493, n35_adj_4494, n33_adj_4495, 
        n11_adj_4496, n13_adj_4497;
    wire [12:0]n9894;
    
    wire n32211, n15_adj_4498, n27_adj_4499, n9_adj_4500, n17_adj_4501, 
        n32210, n19_adj_4502, n21_adj_4503, n39407, n39399, n12_adj_4504, 
        n32209, n10_adj_4505, n30_adj_4506, n39417, n39683, n39679, 
        n39980, n39819, n32208, n40040, n16_adj_4507, n6_adj_4508, 
        n39956, n39957, n8_adj_4509, n24_adj_4510, n39383, n39381, 
        n39855, n39912, n4_adj_4511, n39954, n39955, n39394, n39392, 
        n40050, n39914, n40101, n40102, n40081, n39385, n40010, 
        n40_adj_4512, n40012, n32207, n32206, n30765, n32205, n32204, 
        n32203, n30937;
    wire [12:0]n12912;
    
    wire n30999, n32202, n30764, n32201, n32200, n30812, n30936;
    wire [13:0]n9878;
    
    wire n32199, n30998, n32198, n32197, n30935, n32196, n32195, 
        n30811, n32194, n32193, n30727, n30763, n32192, n32191, 
        n30934, n30997, n32190, n32189, n30810, n30933, n32188, 
        n32187, n30726;
    wire [14:0]n9861;
    
    wire n32186, n32185, n32184, n30809, n32183, n30762, n32182, 
        n32181, n32180, n30808, n32179, n32178, n32177, n30932, 
        n31521, n31520, n32176, n32175, n32174, n31519, n30807, 
        n32173, n31518, n30996, n30931, n31517, n31516;
    wire [15:0]n9843;
    
    wire n32172, n30930, n32171, n32170, n32169, n30995, n30994, 
        n32168, n31515, n31514, n30929, n31513, n30806, n30725, 
        n30928, n31512, n32167, n32166, n32165, n606_adj_4514, n32164, 
        n533_adj_4515, n32163, n460, n32162, n387, n32161, n314, 
        n32160, n241, n32159, n168, n32158, n26_adj_4516, n95;
    wire [16:0]n9824;
    
    wire n32157, n32156, n1114_adj_4517, n32155, n1041_adj_4518, n32154, 
        n612_adj_4519, n30993, n968_adj_4520, n32153, n895_adj_4521, 
        n32152, n822_adj_4522, n32151, n30927, n950, n31511, n749_adj_4524, 
        n32150, n676_adj_4525, n32149, n603_adj_4526, n32148, n530_adj_4527, 
        n32147, n457_adj_4528, n32146, n384_adj_4529, n32145, n311_adj_4530, 
        n32144, n238_adj_4531, n32143, n165_adj_4532, n32142, n23_adj_4533, 
        n92_adj_4534;
    wire [17:0]n9804;
    
    wire n32141, n32140, n32139, n1111_adj_4535, n32138, n1038_adj_4536, 
        n32137, n965_adj_4537, n32136, n539_adj_4538, n30992, n892_adj_4539, 
        n32135, n819_adj_4540, n32134, n746_adj_4541, n32133, n673_adj_4542, 
        n32132, n600_adj_4543, n32131, n527_adj_4544, n32130, n454_adj_4545, 
        n32129, n30805, n381_adj_4546, n32128, n30724, n308_adj_4548, 
        n32127, n235_adj_4549, n32126, n162_adj_4550, n32125, n20_adj_4551, 
        n89_adj_4552;
    wire [18:0]n9783;
    
    wire n32124, n32123, n32122, n32121, n1108_adj_4553, n32120, 
        n1035_adj_4554, n32119, n962_adj_4555, n32118, n889_adj_4556, 
        n32117, n30723, n816_adj_4557, n32116, n743_adj_4558, n32115, 
        n30926, n670_adj_4560, n32114, n597_adj_4561, n32113, n524_adj_4562, 
        n32112, n30804, n451_adj_4563, n32111, n30925, n378_adj_4565, 
        n32110, n469_adj_4566, n30803, n30924, n466_adj_4568, n30991, 
        n30722, n393_adj_4569, n30990, n30923, n30802, n30721, n305_adj_4573, 
        n32109, n232_adj_4574, n32108, n159_adj_4575, n32107, n17_adj_4576, 
        n86_adj_4577;
    wire [19:0]n9761;
    
    wire n32106, n32105, n32104, n32103, n32102, n1105_adj_4578, 
        n32101, n1032_adj_4579, n32100, n959_adj_4580, n32099, n886_adj_4581, 
        n32098, n813_adj_4582, n32097, n740_adj_4583, n32096, n667_adj_4584, 
        n32095, n594_adj_4585, n32094, n521_adj_4586, n32093, n448_adj_4587, 
        n32092, n30922, n375_adj_4589, n32091, n30921, n320_adj_4591, 
        n30989, n302_adj_4592, n32090, n229_adj_4593, n32089, n156_adj_4594, 
        n32088, n14_adj_4595, n83_adj_4596;
    wire [20:0]n9738;
    
    wire n32087, n32086, n32085, n32084, n32083, n32082, n1102_adj_4597, 
        n32081, n1029_adj_4598, n32080, n956_adj_4599, n32079, n883_adj_4600, 
        n32078, n810_adj_4601, n32077, n737_adj_4602, n32076, n664_adj_4603, 
        n32075, n591_adj_4604, n32074, n518_adj_4605, n32073, n445_adj_4606, 
        n32072, n372_adj_4607, n32071, n299_adj_4608, n32070, n247_adj_4609, 
        n30988, n226_adj_4610, n32069, n153_adj_4611, n32068, n30801, 
        n11_adj_4612, n80_adj_4613;
    wire [21:0]n9714;
    
    wire n32067, n32066, n32065, n32064, n174_adj_4614, n30987, 
        n32063, n32062, n32061, n32060, n1096_adj_4615, n32059, 
        n1023_adj_4616, n32058, n950_adj_4617, n32057, n877, n32056, 
        n804, n32055, n731, n32054, n30800, n658_adj_4618, n32053, 
        n585_adj_4619, n32052, n512_adj_4620, n32051, n439_adj_4621, 
        n32050, n366_adj_4622, n32049, n30720, n293_adj_4623, n32048, 
        n220_adj_4624, n32047, n147_adj_4625, n32046, n5_adj_4626, 
        n74_adj_4627, n32045, n32044, n32043, n32042, n32041, n32040, 
        n32039, n1099_adj_4628, n32038, n1026_adj_4629, n32037, n542_adj_4631, 
        n953_adj_4632, n32036, n880_adj_4633, n32035, n807_adj_4634, 
        n32034, n30920, n734_adj_4636, n32033, n32_adj_4637, n101_adj_4638, 
        n661_adj_4639, n32032, n588_adj_4640, n32031, n515_adj_4641, 
        n32030, n442_adj_4642, n32029, n369_adj_4643, n32028, n296_adj_4644, 
        n32027, n223_adj_4645, n32026, n30799, n150_adj_4646, n32025, 
        n30719, n8_adj_4647, n77_adj_4648, n30919, n30798, n30918, 
        n980_adj_4651, n30986, n30917, n615_adj_4653, n731_adj_4655, 
        n31509, n30797, n907_adj_4656, n30985, n834_adj_4657, n30984, 
        n688_adj_4658, n804_adj_4660, n31510, n877_adj_4661, n30916, 
        n30718, n840_adj_4663, n32002, n767_adj_4664, n32001, n694_adj_4665, 
        n32000, n621_adj_4666, n31999, n548_adj_4667, n31998, n475_adj_4668, 
        n31997, n402_adj_4669, n31996, n30915, n329_adj_4671, n31995, 
        n30796, n256_adj_4672, n31994, n183_adj_4673, n31993, n41_adj_4674, 
        n110_adj_4675, n761_adj_4676, n30983, n30914, n30982, n30913, 
        n30981, n30980, n30795, n30912, n30979, n30717, n30911, 
        n30794, n30978, n30910, n30977, n30909, n30845, n30976, 
        n30975, n30844, n30843, n30908, n30842;
    wire [7:0]n13522;
    
    wire n31088, n31087, n31086, n31085, n31084, n31083, n31082, 
        n31081;
    wire [15:0]n12255;
    
    wire n31080, n31079, n31078, n31077, n31076, n31075, n31074, 
        n31073, n31072, n31071, n31070, n30841, n31069, n31068, 
        n30907, n31067, n31066, n31065, n30906, n31064, n31063, 
        n31062, n31061, n536_adj_4677, n31060, n609_adj_4678, n682_adj_4679, 
        n31059, n755_adj_4680, n828_adj_4681, n31058, n31057, n31056, 
        n901_adj_4682, n31055, n974_adj_4683, n460_adj_4684, n31054, 
        n387_adj_4685, n31053, n314_adj_4686, n31052, n241_adj_4687, 
        n31051, n168_adj_4688, n31050, n26_adj_4689, n95_adj_4690, 
        n630_adj_4691, n31049, n557_adj_4692, n31048, n484_adj_4693, 
        n31047, n411_adj_4694, n31046, n338_adj_4696, n31045, n265_adj_4697, 
        n31044, n192_adj_4698, n31043, n50_adj_4699, n119_adj_4700, 
        n1047_adj_4701, n1120_adj_4702, n31042, n31041, n31040, n31039, 
        n31038, n31037, n31036, n31035, n4_adj_4703, n30468, n30427, 
        n30386, n30561, n30595;
    
    SB_CARRY mult_10_add_1225_10 (.CI(n31507), .I0(n9589[7]), .I1(n658), 
            .CO(n31508));
    SB_LUT4 mult_10_add_1225_9_lut (.I0(GND_net), .I1(n9589[6]), .I2(n585), 
            .I3(n31506), .O(n106[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1[5]), .I3(n30904), .O(n11)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_9 (.CI(n31506), .I0(n9589[6]), .I1(n585), 
            .CO(n31507));
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_8_lut (.I0(GND_net), .I1(n9589[5]), .I2(n512), 
            .I3(n31505), .O(n106[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[6]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_10_add_1225_8 (.CI(n31505), .I0(n9589[5]), .I1(n512), 
            .CO(n31506));
    SB_LUT4 i19140_2_lut (.I0(n28[13]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[13]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19140_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_7_lut (.I0(GND_net), .I1(n9589[4]), .I2(n439), 
            .I3(n31504), .O(n106[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_7 (.CI(n31504), .I0(n9589[4]), .I1(n439), 
            .CO(n31505));
    SB_CARRY add_5300_7 (.CI(n31033), .I0(n12717[4]), .I1(n463), .CO(n31034));
    SB_CARRY unary_minus_5_add_3_7 (.CI(n30904), .I0(GND_net), .I1(n1[5]), 
            .CO(n30905));
    SB_LUT4 mult_10_add_1225_6_lut (.I0(GND_net), .I1(n9589[3]), .I2(n366), 
            .I3(n31503), .O(n106[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[7]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [18]), 
            .I2(n9993[0]), .I3(n30518), .O(n9986[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[8]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[9]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19141_2_lut (.I0(n28[14]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[14]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19141_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[10]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_4283));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19142_2_lut (.I0(n28[15]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[15]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19142_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19143_2_lut (.I0(n28[16]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[16]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19143_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[11]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19144_2_lut (.I0(n28[17]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[17]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19144_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[12]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685_adj_4288));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19145_2_lut (.I0(n28[18]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[18]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19145_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758_adj_4289));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831_adj_4290));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[13]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_4292));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977_adj_4293));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[14]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19146_2_lut (.I0(n28[19]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[19]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19146_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050_adj_4295));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[15]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_6 (.CI(n31503), .I0(n9589[3]), .I1(n366), 
            .CO(n31504));
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_4297));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22150_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [18]), 
            .I2(n30518), .I3(n9993[0]), .O(n4));   // verilog/motorControl.v(34[25:36])
    defparam i22150_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i2_3_lut (.I0(duty_23__N_3613[1]), .I1(n257[1]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_add_1225_5_lut (.I0(GND_net), .I1(n9589[2]), .I2(n293), 
            .I3(n31502), .O(n106[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i2_3_lut (.I0(duty_23__N_3588[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_5 (.CI(n31502), .I0(n9589[2]), .I1(n293), 
            .CO(n31503));
    SB_LUT4 mult_10_add_1225_4_lut (.I0(GND_net), .I1(n9589[1]), .I2(n220), 
            .I3(n31501), .O(n106[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_4 (.CI(n31501), .I0(n9589[1]), .I1(n220), 
            .CO(n31502));
    SB_LUT4 mult_10_add_1225_3_lut (.I0(GND_net), .I1(n9589[0]), .I2(n147_adj_4298), 
            .I3(n31500), .O(n106[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_3 (.CI(n31500), .I0(n9589[0]), .I1(n147_adj_4298), 
            .CO(n31501));
    SB_LUT4 mult_10_add_1225_2_lut (.I0(GND_net), .I1(n5), .I2(n74), .I3(GND_net), 
            .O(n106[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5), .I1(n74), .CO(n31500));
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5070_23_lut (.I0(GND_net), .I1(n10450[20]), .I2(GND_net), 
            .I3(n31499), .O(n9589[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19147_2_lut (.I0(n28[20]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[20]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19147_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22139_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3513 [18]), .I3(\Ki[1] ), 
            .O(n30518));   // verilog/motorControl.v(34[25:36])
    defparam i22139_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_4299));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_4300));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_4301));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253_adj_4302));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_4303));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_4304));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_4305));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_4306));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5070_22_lut (.I0(GND_net), .I1(n10450[19]), .I2(GND_net), 
            .I3(n31498), .O(n9589[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_4307));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898_adj_4308));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971_adj_4309));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044_adj_4310));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(n28[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117_adj_4311));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5070_22 (.CI(n31498), .I0(n10450[19]), .I1(GND_net), 
            .CO(n31499));
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5300_6_lut (.I0(GND_net), .I1(n12717[3]), .I2(n390_adj_4315), 
            .I3(n31032), .O(n12509[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5070_21_lut (.I0(GND_net), .I1(n10450[18]), .I2(GND_net), 
            .I3(n31497), .O(n9589[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1[4]), .I3(n30903), .O(n9_adj_4316)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22137_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3513 [18]), .I3(\Ki[1] ), 
            .O(n9986[0]));   // verilog/motorControl.v(34[25:36])
    defparam i22137_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[16]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104_adj_4319));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[17]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4321));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_4322));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_4323));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_4324));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_4325));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_4326));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_4327));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(n28[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4329));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472_adj_4330));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_4331));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5070_21 (.CI(n31497), .I0(n10450[18]), .I1(GND_net), 
            .CO(n31498));
    SB_LUT4 add_5070_20_lut (.I0(GND_net), .I1(n10450[17]), .I2(GND_net), 
            .I3(n31496), .O(n9589[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5070_20 (.CI(n31496), .I0(n10450[17]), .I1(GND_net), 
            .CO(n31497));
    SB_CARRY add_5300_6 (.CI(n31032), .I0(n12717[3]), .I1(n390_adj_4315), 
            .CO(n31033));
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5070_19_lut (.I0(GND_net), .I1(n10450[16]), .I2(GND_net), 
            .I3(n31495), .O(n9589[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5070_19 (.CI(n31495), .I0(n10450[16]), .I1(GND_net), 
            .CO(n31496));
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5300_5_lut (.I0(GND_net), .I1(n12717[2]), .I2(n317_adj_4332), 
            .I3(n31031), .O(n12509[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[18]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5070_18_lut (.I0(GND_net), .I1(n10450[15]), .I2(GND_net), 
            .I3(n31494), .O(n9589[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_18 (.CI(n31494), .I0(n10450[15]), .I1(GND_net), 
            .CO(n31495));
    SB_LUT4 add_5070_17_lut (.I0(GND_net), .I1(n10450[14]), .I2(GND_net), 
            .I3(n31493), .O(n9589[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5070_17 (.CI(n31493), .I0(n10450[14]), .I1(GND_net), 
            .CO(n31494));
    SB_LUT4 add_5070_16_lut (.I0(GND_net), .I1(n10450[13]), .I2(n1099), 
            .I3(n31492), .O(n9589[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(n28[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4334));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n30903), .I0(GND_net), .I1(n1[4]), 
            .CO(n30904));
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5070_16 (.CI(n31492), .I0(n10450[13]), .I1(n1099), .CO(n31493));
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5070_15_lut (.I0(GND_net), .I1(n10450[12]), .I2(n1026), 
            .I3(n31491), .O(n9589[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5070_15 (.CI(n31491), .I0(n10450[12]), .I1(n1026), .CO(n31492));
    SB_CARRY add_5300_5 (.CI(n31031), .I0(n12717[2]), .I1(n317_adj_4332), 
            .CO(n31032));
    SB_LUT4 add_5300_4_lut (.I0(GND_net), .I1(n12717[1]), .I2(n244_adj_4335), 
            .I3(n31030), .O(n12509[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1[3]), .I3(n30902), .O(n7_adj_4336)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n30902), .I0(GND_net), .I1(n1[3]), 
            .CO(n30903));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1[2]), .I3(n30901), .O(n5_adj_4338)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_4340));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_4341));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_4342));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5070_14_lut (.I0(GND_net), .I1(n10450[11]), .I2(n953), 
            .I3(n31490), .O(n9589[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_14 (.CI(n31490), .I0(n10450[11]), .I1(n953), .CO(n31491));
    SB_LUT4 add_5070_13_lut (.I0(GND_net), .I1(n10450[10]), .I2(n880), 
            .I3(n31489), .O(n9589[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_13 (.CI(n31489), .I0(n10450[10]), .I1(n880), .CO(n31490));
    SB_LUT4 add_5070_12_lut (.I0(GND_net), .I1(n10450[9]), .I2(n807), 
            .I3(n31488), .O(n9589[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_12 (.CI(n31488), .I0(n10450[9]), .I1(n807), .CO(n31489));
    SB_LUT4 add_5070_11_lut (.I0(GND_net), .I1(n10450[8]), .I2(n734), 
            .I3(n31487), .O(n9589[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_11 (.CI(n31487), .I0(n10450[8]), .I1(n734), .CO(n31488));
    SB_LUT4 add_5070_10_lut (.I0(GND_net), .I1(n10450[7]), .I2(n661), 
            .I3(n31486), .O(n9589[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_10 (.CI(n31486), .I0(n10450[7]), .I1(n661), .CO(n31487));
    SB_LUT4 add_5070_9_lut (.I0(GND_net), .I1(n10450[6]), .I2(n588), .I3(n31485), 
            .O(n9589[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_9 (.CI(n31485), .I0(n10450[6]), .I1(n588), .CO(n31486));
    SB_LUT4 add_5070_8_lut (.I0(GND_net), .I1(n10450[5]), .I2(n515), .I3(n31484), 
            .O(n9589[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_8 (.CI(n31484), .I0(n10450[5]), .I1(n515), .CO(n31485));
    SB_LUT4 add_5070_7_lut (.I0(GND_net), .I1(n10450[4]), .I2(n442), .I3(n31483), 
            .O(n9589[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_7 (.CI(n31483), .I0(n10450[4]), .I1(n442), .CO(n31484));
    SB_LUT4 add_5070_6_lut (.I0(GND_net), .I1(n10450[3]), .I2(n369), .I3(n31482), 
            .O(n9589[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_6 (.CI(n31482), .I0(n10450[3]), .I1(n369), .CO(n31483));
    SB_LUT4 add_5070_5_lut (.I0(GND_net), .I1(n10450[2]), .I2(n296), .I3(n31481), 
            .O(n9589[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113_adj_4343));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44_adj_4344));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4345));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4346));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_4347));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_4348));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414_adj_4349));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_4350));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405_adj_4351));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4352));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4353));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_4354));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_4355));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_4356));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(n28[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4358));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5070_5 (.CI(n31481), .I0(n10450[2]), .I1(n296), .CO(n31482));
    SB_LUT4 add_5070_4_lut (.I0(GND_net), .I1(n10450[1]), .I2(n223), .I3(n31480), 
            .O(n9589[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_4 (.CI(n31480), .I0(n10450[1]), .I1(n223), .CO(n31481));
    SB_LUT4 add_5070_3_lut (.I0(GND_net), .I1(n10450[0]), .I2(n150_adj_4359), 
            .I3(n31479), .O(n9589[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_3 (.CI(n31479), .I0(n10450[0]), .I1(n150_adj_4359), 
            .CO(n31480));
    SB_LUT4 add_5070_2_lut (.I0(GND_net), .I1(n8_adj_4360), .I2(n77), 
            .I3(GND_net), .O(n9589[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5070_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5070_2 (.CI(GND_net), .I0(n8_adj_4360), .I1(n77), .CO(n31479));
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5195_22_lut (.I0(GND_net), .I1(n10889[19]), .I2(GND_net), 
            .I3(n31478), .O(n10450[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5195_21_lut (.I0(GND_net), .I1(n10889[18]), .I2(GND_net), 
            .I3(n31477), .O(n10450[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5195_21 (.CI(n31477), .I0(n10889[18]), .I1(GND_net), 
            .CO(n31478));
    SB_LUT4 add_5195_20_lut (.I0(GND_net), .I1(n10889[17]), .I2(GND_net), 
            .I3(n31476), .O(n10450[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_20 (.CI(n31476), .I0(n10889[17]), .I1(GND_net), 
            .CO(n31477));
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98_adj_4362));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4363));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5195_19_lut (.I0(GND_net), .I1(n10889[16]), .I2(GND_net), 
            .I3(n31475), .O(n10450[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(n28[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4364));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_4365));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_4366));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171_adj_4367));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_4368));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4370));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n6_adj_4371), .I1(\Ki[4] ), .I2(n9993[2]), .I3(\PID_CONTROLLER.integral_23__N_3513 [18]), 
            .O(n9986[3]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4372));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_4373));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22230_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3513 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3513 [21]), .O(n10004[0]));   // verilog/motorControl.v(34[25:36])
    defparam i22230_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(n28[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_4374));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1511 (.I0(n4_adj_4375), .I1(\Ki[3] ), .I2(n9999[1]), 
            .I3(\PID_CONTROLLER.integral_23__N_3513 [19]), .O(n9993[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1511.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_4376));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1512 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral_23__N_3513 [23]), 
            .I3(\PID_CONTROLLER.integral_23__N_3513 [20]), .O(n12_adj_4377));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1512.LUT_INIT = 16'h9c50;
    SB_LUT4 i22166_4_lut (.I0(n9993[2]), .I1(\Ki[4] ), .I2(n6_adj_4371), 
            .I3(\PID_CONTROLLER.integral_23__N_3513 [18]), .O(n8_adj_4378));   // verilog/motorControl.v(34[25:36])
    defparam i22166_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3513 [19]), 
            .I3(\PID_CONTROLLER.integral_23__N_3513 [21]), .O(n11_adj_4379));   // verilog/motorControl.v(34[25:36])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i22197_4_lut (.I0(n9999[1]), .I1(\Ki[3] ), .I2(n4_adj_4375), 
            .I3(\PID_CONTROLLER.integral_23__N_3513 [19]), .O(n6_adj_4380));   // verilog/motorControl.v(34[25:36])
    defparam i22197_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i22232_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3513 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3513 [21]), .O(n30620));   // verilog/motorControl.v(34[25:36])
    defparam i22232_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut (.I0(n6_adj_4380), .I1(n11_adj_4379), .I2(n8_adj_4378), 
            .I3(n12_adj_4377), .O(n18_adj_4381));   // verilog/motorControl.v(34[25:36])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3513 [18]), 
            .I3(\PID_CONTROLLER.integral_23__N_3513 [22]), .O(n13_adj_4382));   // verilog/motorControl.v(34[25:36])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut (.I0(n13_adj_4382), .I1(n18_adj_4381), .I2(n30620), 
            .I3(n4_adj_4383), .O(n37896));   // verilog/motorControl.v(34[25:36])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5195_19 (.CI(n31475), .I0(n10889[16]), .I1(GND_net), 
            .CO(n31476));
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[19]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545_adj_4385));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19148_2_lut (.I0(n28[21]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[21]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19148_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[20]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5195_18_lut (.I0(GND_net), .I1(n10889[15]), .I2(GND_net), 
            .I3(n31474), .O(n10450[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_4388));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5195_18 (.CI(n31474), .I0(n10889[15]), .I1(GND_net), 
            .CO(n31475));
    SB_LUT4 add_5195_17_lut (.I0(GND_net), .I1(n10889[14]), .I2(GND_net), 
            .I3(n31473), .O(n10450[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_17 (.CI(n31473), .I0(n10889[14]), .I1(GND_net), 
            .CO(n31474));
    SB_LUT4 add_5195_16_lut (.I0(GND_net), .I1(n10889[13]), .I2(n1102), 
            .I3(n31472), .O(n10450[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_16 (.CI(n31472), .I0(n10889[13]), .I1(n1102), .CO(n31473));
    SB_LUT4 add_5195_15_lut (.I0(GND_net), .I1(n10889[12]), .I2(n1029), 
            .I3(n31471), .O(n10450[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_15 (.CI(n31471), .I0(n10889[12]), .I1(n1029), .CO(n31472));
    SB_LUT4 add_5195_14_lut (.I0(GND_net), .I1(n10889[11]), .I2(n956), 
            .I3(n31470), .O(n10450[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_14 (.CI(n31470), .I0(n10889[11]), .I1(n956), .CO(n31471));
    SB_CARRY add_5300_4 (.CI(n31030), .I0(n12717[1]), .I1(n244_adj_4335), 
            .CO(n31031));
    SB_LUT4 add_5195_13_lut (.I0(GND_net), .I1(n10889[10]), .I2(n883), 
            .I3(n31469), .O(n10450[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_13 (.CI(n31469), .I0(n10889[10]), .I1(n883), .CO(n31470));
    SB_LUT4 add_5195_12_lut (.I0(GND_net), .I1(n10889[9]), .I2(n810), 
            .I3(n31468), .O(n10450[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3489[0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i0  (.Q(\PID_CONTROLLER.integral [0]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY unary_minus_5_add_3_4 (.CI(n30901), .I0(GND_net), .I1(n1[2]), 
            .CO(n30902));
    SB_CARRY add_5195_12 (.CI(n31468), .I0(n10889[9]), .I1(n810), .CO(n31469));
    SB_LUT4 add_5195_11_lut (.I0(GND_net), .I1(n10889[8]), .I2(n737), 
            .I3(n31467), .O(n10450[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_11 (.CI(n31467), .I0(n10889[8]), .I1(n737), .CO(n31468));
    SB_LUT4 add_5195_10_lut (.I0(GND_net), .I1(n10889[7]), .I2(n664), 
            .I3(n31466), .O(n10450[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_10 (.CI(n31466), .I0(n10889[7]), .I1(n664), .CO(n31467));
    SB_LUT4 add_5195_9_lut (.I0(GND_net), .I1(n10889[6]), .I2(n591), .I3(n31465), 
            .O(n10450[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_9 (.CI(n31465), .I0(n10889[6]), .I1(n591), .CO(n31466));
    SB_LUT4 add_5195_8_lut (.I0(GND_net), .I1(n10889[5]), .I2(n518), .I3(n31464), 
            .O(n10450[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_8 (.CI(n31464), .I0(n10889[5]), .I1(n518), .CO(n31465));
    SB_LUT4 add_5195_7_lut (.I0(GND_net), .I1(n10889[4]), .I2(n445), .I3(n31463), 
            .O(n10450[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_7 (.CI(n31463), .I0(n10889[4]), .I1(n445), .CO(n31464));
    SB_LUT4 add_5195_6_lut (.I0(GND_net), .I1(n10889[3]), .I2(n372), .I3(n31462), 
            .O(n10450[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_6 (.CI(n31462), .I0(n10889[3]), .I1(n372), .CO(n31463));
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_4389));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5195_5_lut (.I0(GND_net), .I1(n10889[2]), .I2(n299), .I3(n31461), 
            .O(n10450[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_5 (.CI(n31461), .I0(n10889[2]), .I1(n299), .CO(n31462));
    SB_LUT4 add_5195_4_lut (.I0(GND_net), .I1(n10889[1]), .I2(n226), .I3(n31460), 
            .O(n10450[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_4 (.CI(n31460), .I0(n10889[1]), .I1(n226), .CO(n31461));
    SB_LUT4 i19149_2_lut (.I0(n28[22]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[22]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5195_3_lut (.I0(GND_net), .I1(n10889[0]), .I2(n153_adj_4370), 
            .I3(n31459), .O(n10450[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_3 (.CI(n31459), .I0(n10889[0]), .I1(n153_adj_4370), 
            .CO(n31460));
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1[1]), .I3(n30900), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5300_3_lut (.I0(GND_net), .I1(n12717[0]), .I2(n171_adj_4367), 
            .I3(n31029), .O(n12509[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5195_2_lut (.I0(GND_net), .I1(n11_adj_4364), .I2(n80), 
            .I3(GND_net), .O(n10450[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5195_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5195_2 (.CI(GND_net), .I0(n11_adj_4364), .I1(n80), .CO(n31459));
    SB_LUT4 add_5215_21_lut (.I0(GND_net), .I1(n11287[18]), .I2(GND_net), 
            .I3(n31458), .O(n10889[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17_adj_4391));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_4392));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_4393));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29468_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n39496));
    defparam i29468_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i29465_3_lut (.I0(n11_adj_4393), .I1(n9_adj_4392), .I2(n39496), 
            .I3(GND_net), .O(n39493));
    defparam i29465_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 add_5215_20_lut (.I0(GND_net), .I1(n11287[17]), .I2(GND_net), 
            .I3(n31457), .O(n10889[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_196_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n41474));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_196_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29838_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n41474), 
            .I2(IntegralLimit[7]), .I3(n39493), .O(n39867));
    defparam i29838_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_5215_20 (.CI(n31457), .I0(n11287[17]), .I1(GND_net), 
            .CO(n31458));
    SB_LUT4 i29717_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4391), 
            .I2(IntegralLimit[9]), .I3(n39867), .O(n39746));
    defparam i29717_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_178_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n41456));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_178_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29715_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4391), 
            .I2(IntegralLimit[9]), .I3(n9_adj_4392), .O(n39744));
    defparam i29715_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i29713_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n41456), 
            .I2(IntegralLimit[11]), .I3(n39744), .O(n39742));
    defparam i29713_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 add_5215_19_lut (.I0(GND_net), .I1(n11287[16]), .I2(GND_net), 
            .I3(n31456), .O(n10889[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_172_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n41450));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_172_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29408_4_lut (.I0(n27), .I1(n15_adj_4394), .I2(n13_adj_4395), 
            .I3(n11), .O(n39436));
    defparam i29408_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29414_4_lut (.I0(n21_adj_4396), .I1(n19_adj_4397), .I2(n17_adj_4398), 
            .I3(n9_adj_4316), .O(n39442));
    defparam i29414_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_5215_19 (.CI(n31456), .I0(n11287[16]), .I1(GND_net), 
            .CO(n31457));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43), .I3(GND_net), 
            .O(n16_adj_4399));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 add_5215_18_lut (.I0(GND_net), .I1(n11287[15]), .I2(GND_net), 
            .I3(n31455), .O(n10889[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29391_2_lut (.I0(n43), .I1(n19_adj_4397), .I2(GND_net), .I3(GND_net), 
            .O(n39419));
    defparam i29391_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_4398), .I3(GND_net), 
            .O(n8_adj_4400));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_CARRY add_5215_18 (.CI(n31455), .I0(n11287[15]), .I1(GND_net), 
            .CO(n31456));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_4399), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45), .I3(GND_net), 
            .O(n24_adj_4401));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i29424_2_lut (.I0(n7_adj_4336), .I1(n5_adj_4338), .I2(GND_net), 
            .I3(GND_net), .O(n39452));
    defparam i29424_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n30900), .I0(GND_net), .I1(n1[1]), 
            .CO(n30901));
    SB_LUT4 add_5215_17_lut (.I0(GND_net), .I1(n11287[14]), .I2(GND_net), 
            .I3(n31454), .O(n10889[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29686_4_lut (.I0(n13_adj_4395), .I1(n11), .I2(n9_adj_4316), 
            .I3(n39452), .O(n39715));
    defparam i29686_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i29682_4_lut (.I0(n19_adj_4397), .I1(n17_adj_4398), .I2(n15_adj_4394), 
            .I3(n39715), .O(n39711));
    defparam i29682_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i29959_4_lut (.I0(n25_adj_4402), .I1(n23_adj_4403), .I2(n21_adj_4396), 
            .I3(n39711), .O(n39988));
    defparam i29959_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i29806_4_lut (.I0(n31), .I1(n29_adj_4404), .I2(n27), .I3(n39988), 
            .O(n39835));
    defparam i29806_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i30013_4_lut (.I0(n37), .I1(n35_adj_4405), .I2(n33), .I3(n39835), 
            .O(n40042));
    defparam i30013_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_5300_3 (.CI(n31029), .I0(n12717[0]), .I1(n171_adj_4367), 
            .CO(n31030));
    SB_CARRY add_5215_17 (.CI(n31454), .I0(n11287[14]), .I1(GND_net), 
            .CO(n31455));
    SB_LUT4 i29719_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n41474), 
            .I2(IntegralLimit[7]), .I3(n11_adj_4393), .O(n39748));
    defparam i29719_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3564 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_165_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n41443));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_165_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29707_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n41443), 
            .I2(IntegralLimit[14]), .I3(n39748), .O(n39736));
    defparam i29707_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 add_5215_16_lut (.I0(GND_net), .I1(n11287[13]), .I2(n1105), 
            .I3(n31453), .O(n10889[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_159_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n41437));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_159_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_4406));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5215_16 (.CI(n31453), .I0(n11287[13]), .I1(n1105), .CO(n31454));
    SB_LUT4 add_5215_15_lut (.I0(GND_net), .I1(n11287[12]), .I2(n1032), 
            .I3(n31452), .O(n10889[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5300_2_lut (.I0(GND_net), .I1(n29_adj_4363), .I2(n98_adj_4362), 
            .I3(GND_net), .O(n12509[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29441_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n39469));
    defparam i29441_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_183_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n41461));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_183_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_4407));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5215_15 (.CI(n31452), .I0(n11287[12]), .I1(n1032), .CO(n31453));
    SB_LUT4 add_5215_14_lut (.I0(GND_net), .I1(n11287[11]), .I2(n959), 
            .I3(n31451), .O(n10889[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5215_14 (.CI(n31451), .I0(n11287[11]), .I1(n959), .CO(n31452));
    SB_LUT4 add_5215_13_lut (.I0(GND_net), .I1(n11287[10]), .I2(n886), 
            .I3(n31450), .O(n10889[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_4406), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5215_13 (.CI(n31450), .I0(n11287[10]), .I1(n886), .CO(n31451));
    SB_LUT4 add_5215_12_lut (.I0(GND_net), .I1(n11287[9]), .I2(n813), 
            .I3(n31449), .O(n10889[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5215_12 (.CI(n31449), .I0(n11287[9]), .I1(n813), .CO(n31450));
    SB_LUT4 add_5215_11_lut (.I0(GND_net), .I1(n11287[8]), .I2(n740), 
            .I3(n31448), .O(n10889[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29904_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n41456), 
            .I2(IntegralLimit[11]), .I3(n39746), .O(n39933));
    defparam i29904_4_lut.LUT_INIT = 16'hffde;
    SB_CARRY add_5215_11 (.CI(n31448), .I0(n11287[8]), .I1(n740), .CO(n31449));
    SB_LUT4 i29453_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n41450), 
            .I2(IntegralLimit[13]), .I3(n39933), .O(n39481));
    defparam i29453_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_163_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n41441));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_163_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5215_10_lut (.I0(GND_net), .I1(n11287[7]), .I2(n667), 
            .I3(n31447), .O(n10889[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29830_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n41441), 
            .I2(IntegralLimit[15]), .I3(n39481), .O(n39859));
    defparam i29830_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_189_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n41467));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_189_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1[0]), 
            .CO(n30900));
    SB_LUT4 i29965_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n41467), 
            .I2(IntegralLimit[17]), .I3(n39859), .O(n39994));
    defparam i29965_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 sub_3_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(motor_state[23]), 
            .I3(n30899), .O(n28[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5215_10 (.CI(n31447), .I0(n11287[7]), .I1(n667), .CO(n31448));
    SB_LUT4 add_5215_9_lut (.I0(GND_net), .I1(n11287[6]), .I2(n594), .I3(n31446), 
            .O(n10889[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5300_2 (.CI(GND_net), .I0(n29_adj_4363), .I1(n98_adj_4362), 
            .CO(n31029));
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_154_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n41432));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_154_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5215_9 (.CI(n31446), .I0(n11287[6]), .I1(n594), .CO(n31447));
    SB_LUT4 sub_3_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(motor_state[22]), 
            .I3(n30898), .O(n28[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30035_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n41432), 
            .I2(IntegralLimit[19]), .I3(n39994), .O(n40064));
    defparam i30035_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_151_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n41429));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_151_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_4410));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29426_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n39454));
    defparam i29426_4_lut.LUT_INIT = 16'h7bde;
    SB_CARRY sub_3_add_2_24 (.CI(n30898), .I0(setpoint[22]), .I1(motor_state[22]), 
            .CO(n30899));
    SB_LUT4 add_5215_8_lut (.I0(GND_net), .I1(n11287[5]), .I2(n521), .I3(n31445), 
            .O(n10889[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_4410), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_4411));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_4412));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5215_8 (.CI(n31445), .I0(n11287[5]), .I1(n521), .CO(n31446));
    SB_LUT4 i29844_3_lut (.I0(n6_adj_4412), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n39873));   // verilog/motorControl.v(31[10:34])
    defparam i29844_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29845_3_lut (.I0(n39873), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n39874));   // verilog/motorControl.v(31[10:34])
    defparam i29845_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5215_7_lut (.I0(GND_net), .I1(n11287[4]), .I2(n448), .I3(n31444), 
            .O(n10889[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5215_7 (.CI(n31444), .I0(n11287[4]), .I1(n448), .CO(n31445));
    SB_LUT4 i29430_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n41450), 
            .I2(IntegralLimit[21]), .I3(n39742), .O(n39458));
    defparam i29430_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 sub_3_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(motor_state[21]), 
            .I3(n30897), .O(n28[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5215_6_lut (.I0(GND_net), .I1(n11287[3]), .I2(n375), .I3(n31443), 
            .O(n10889[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29822_4_lut (.I0(n24_adj_4411), .I1(n8_adj_4413), .I2(n41427), 
            .I3(n39454), .O(n39851));   // verilog/motorControl.v(31[10:34])
    defparam i29822_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_5215_6 (.CI(n31443), .I0(n11287[3]), .I1(n375), .CO(n31444));
    SB_LUT4 add_5215_5_lut (.I0(GND_net), .I1(n11287[2]), .I2(n302), .I3(n31442), 
            .O(n10889[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29705_3_lut (.I0(n39874), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n39734));   // verilog/motorControl.v(31[10:34])
    defparam i29705_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_5215_5 (.CI(n31442), .I0(n11287[2]), .I1(n302), .CO(n31443));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3564 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_4414));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 add_5215_4_lut (.I0(GND_net), .I1(n11287[1]), .I2(n229), .I3(n31441), 
            .O(n10889[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29937_3_lut (.I0(n4_adj_4414), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27), .I3(GND_net), .O(n39966));   // verilog/motorControl.v(31[38:63])
    defparam i29937_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5215_4 (.CI(n31441), .I0(n11287[1]), .I1(n229), .CO(n31442));
    SB_LUT4 add_5215_3_lut (.I0(GND_net), .I1(n11287[0]), .I2(n156), .I3(n31440), 
            .O(n10889[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29938_3_lut (.I0(n39966), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29_adj_4404), .I3(GND_net), .O(n39967));   // verilog/motorControl.v(31[38:63])
    defparam i29938_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY sub_3_add_2_23 (.CI(n30897), .I0(setpoint[21]), .I1(motor_state[21]), 
            .CO(n30898));
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4415));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33), .I3(GND_net), 
            .O(n12_adj_4416));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i29401_2_lut (.I0(n33), .I1(n15_adj_4394), .I2(GND_net), .I3(GND_net), 
            .O(n39429));
    defparam i29401_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_4395), .I3(GND_net), 
            .O(n10_adj_4417));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_4416), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35_adj_4405), .I3(GND_net), 
            .O(n30_adj_4418));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i29403_4_lut (.I0(n33), .I1(n31), .I2(n29_adj_4404), .I3(n39436), 
            .O(n39431));
    defparam i29403_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30019_4_lut (.I0(n30_adj_4418), .I1(n10_adj_4417), .I2(n35_adj_4405), 
            .I3(n39429), .O(n40048));   // verilog/motorControl.v(31[38:63])
    defparam i30019_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_4419));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1513 (.I0(n6_adj_4420), .I1(\Kp[4] ), .I2(n13692[2]), 
            .I3(n28[18]), .O(n13668[3]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1513.LUT_INIT = 16'h965a;
    SB_CARRY add_5215_3 (.CI(n31440), .I0(n11287[0]), .I1(n156), .CO(n31441));
    SB_LUT4 i29879_3_lut (.I0(n39967), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31), .I3(GND_net), .O(n39908));   // verilog/motorControl.v(31[38:63])
    defparam i29879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30070_4_lut (.I0(n39908), .I1(n40048), .I2(n35_adj_4405), 
            .I3(n39431), .O(n40099));   // verilog/motorControl.v(31[38:63])
    defparam i30070_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30071_3_lut (.I0(n40099), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37), .I3(GND_net), .O(n40100));   // verilog/motorControl.v(31[38:63])
    defparam i30071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30054_3_lut (.I0(n40100), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39), .I3(GND_net), .O(n40083));   // verilog/motorControl.v(31[38:63])
    defparam i30054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_4336), .I3(GND_net), 
            .O(n6_adj_4421));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i29945_3_lut (.I0(n6_adj_4421), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_4396), .I3(GND_net), .O(n39974));   // verilog/motorControl.v(31[38:63])
    defparam i29945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29946_3_lut (.I0(n39974), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_4403), .I3(GND_net), .O(n39975));   // verilog/motorControl.v(31[38:63])
    defparam i29946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29393_4_lut (.I0(n43), .I1(n25_adj_4402), .I2(n23_adj_4403), 
            .I3(n39442), .O(n39421));
    defparam i29393_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29824_4_lut (.I0(n24_adj_4401), .I1(n8_adj_4400), .I2(n45), 
            .I3(n39419), .O(n39853));   // verilog/motorControl.v(31[38:63])
    defparam i29824_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29877_3_lut (.I0(n39975), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_4402), .I3(GND_net), .O(n39906));   // verilog/motorControl.v(31[38:63])
    defparam i29877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29395_4_lut (.I0(n43), .I1(n41_adj_4422), .I2(n39), .I3(n40042), 
            .O(n39423));
    defparam i29395_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29975_4_lut (.I0(n39906), .I1(n39853), .I2(n45), .I3(n39421), 
            .O(n40004));   // verilog/motorControl.v(31[38:63])
    defparam i29975_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30040_3_lut (.I0(n40083), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41_adj_4422), .I3(GND_net), .O(n40));   // verilog/motorControl.v(31[38:63])
    defparam i30040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29977_4_lut (.I0(n40), .I1(n40004), .I2(n45), .I3(n39423), 
            .O(n40006));   // verilog/motorControl.v(31[38:63])
    defparam i29977_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_4423));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i29961_3_lut (.I0(n4_adj_4423), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n39990));   // verilog/motorControl.v(31[10:34])
    defparam i29961_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29962_3_lut (.I0(n39990), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n39991));   // verilog/motorControl.v(31[10:34])
    defparam i29962_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29443_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n41437), 
            .I2(IntegralLimit[16]), .I3(n39736), .O(n39471));
    defparam i29443_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i30017_4_lut (.I0(n30), .I1(n10_adj_4407), .I2(n41461), .I3(n39469), 
            .O(n40046));   // verilog/motorControl.v(31[10:34])
    defparam i30017_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29873_3_lut (.I0(n39991), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n39902));   // verilog/motorControl.v(31[10:34])
    defparam i29873_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i30068_4_lut (.I0(n39902), .I1(n40046), .I2(n41461), .I3(n39471), 
            .O(n40097));   // verilog/motorControl.v(31[10:34])
    defparam i30068_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30069_3_lut (.I0(n40097), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n40098));   // verilog/motorControl.v(31[10:34])
    defparam i30069_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i30056_3_lut (.I0(n40098), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n40085));   // verilog/motorControl.v(31[10:34])
    defparam i30056_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29433_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n41429), 
            .I2(IntegralLimit[21]), .I3(n40064), .O(n39461));
    defparam i29433_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_149_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n41427));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_149_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29969_4_lut (.I0(n39734), .I1(n39851), .I2(n41427), .I3(n39458), 
            .O(n39998));   // verilog/motorControl.v(31[10:34])
    defparam i29969_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30038_3_lut (.I0(n40085), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n40_adj_4424));   // verilog/motorControl.v(31[10:34])
    defparam i30038_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29978_3_lut (.I0(n40006), .I1(\PID_CONTROLLER.integral_23__N_3564 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3563 ));   // verilog/motorControl.v(31[38:63])
    defparam i29978_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29971_4_lut (.I0(n40_adj_4424), .I1(n39998), .I2(n41427), 
            .I3(n39461), .O(n40000));   // verilog/motorControl.v(31[10:34])
    defparam i29971_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_830_4_lut  (.I0(n40000), .I1(\PID_CONTROLLER.integral_23__N_3563 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3561 ));   // verilog/motorControl.v(31[10:63])
    defparam \PID_CONTROLLER.integral_23__I_830_4_lut .LUT_INIT = 16'h80c8;
    SB_LUT4 add_5215_2_lut (.I0(GND_net), .I1(n14_adj_4358), .I2(n83), 
            .I3(GND_net), .O(n10889[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5215_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177_adj_4425));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5215_2 (.CI(GND_net), .I0(n14_adj_4358), .I1(n83), .CO(n31440));
    SB_LUT4 add_5359_11_lut (.I0(GND_net), .I1(n13442[8]), .I2(n770_adj_4356), 
            .I3(n31439), .O(n13343[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5359_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5359_10_lut (.I0(GND_net), .I1(n13442[7]), .I2(n697_adj_4355), 
            .I3(n31438), .O(n13343[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5359_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(motor_state[20]), 
            .I3(n30896), .O(n28[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5359_10 (.CI(n31438), .I0(n13442[7]), .I1(n697_adj_4355), 
            .CO(n31439));
    SB_LUT4 add_5359_9_lut (.I0(GND_net), .I1(n13442[6]), .I2(n624_adj_4354), 
            .I3(n31437), .O(n13343[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5359_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_22 (.CI(n30896), .I0(setpoint[20]), .I1(motor_state[20]), 
            .CO(n30897));
    SB_CARRY add_5359_9 (.CI(n31437), .I0(n13442[6]), .I1(n624_adj_4354), 
            .CO(n31438));
    SB_LUT4 add_5359_8_lut (.I0(GND_net), .I1(n13442[5]), .I2(n551_adj_4353), 
            .I3(n31436), .O(n13343[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5359_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250_adj_4426));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5359_8 (.CI(n31436), .I0(n13442[5]), .I1(n551_adj_4353), 
            .CO(n31437));
    SB_LUT4 i22038_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n28[22]), .I3(n28[21]), 
            .O(n13712[0]));   // verilog/motorControl.v(34[16:22])
    defparam i22038_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_5359_7_lut (.I0(GND_net), .I1(n13442[4]), .I2(n478_adj_4352), 
            .I3(n31435), .O(n13343[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5359_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(motor_state[19]), 
            .I3(n30895), .O(n28[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5359_7 (.CI(n31435), .I0(n13442[4]), .I1(n478_adj_4352), 
            .CO(n31436));
    SB_LUT4 i19150_2_lut (.I0(n28[23]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[23]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19150_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5359_6_lut (.I0(GND_net), .I1(n13442[3]), .I2(n405_adj_4351), 
            .I3(n31434), .O(n13343[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5359_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5359_6 (.CI(n31434), .I0(n13442[3]), .I1(n405_adj_4351), 
            .CO(n31435));
    SB_LUT4 add_5359_5_lut (.I0(GND_net), .I1(n13442[2]), .I2(n332_adj_4350), 
            .I3(n31433), .O(n13343[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5359_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5359_5 (.CI(n31433), .I0(n13442[2]), .I1(n332_adj_4350), 
            .CO(n31434));
    SB_LUT4 add_5359_4_lut (.I0(GND_net), .I1(n13442[1]), .I2(n259_adj_4347), 
            .I3(n31432), .O(n13343[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5359_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5359_4 (.CI(n31432), .I0(n13442[1]), .I1(n259_adj_4347), 
            .CO(n31433));
    SB_CARRY sub_3_add_2_21 (.CI(n30895), .I0(setpoint[19]), .I1(motor_state[19]), 
            .CO(n30896));
    SB_LUT4 add_5359_3_lut (.I0(GND_net), .I1(n13442[0]), .I2(n186_adj_4345), 
            .I3(n31431), .O(n13343[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5359_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618_adj_4427));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5359_3 (.CI(n31431), .I0(n13442[0]), .I1(n186_adj_4345), 
            .CO(n31432));
    SB_LUT4 add_5359_2_lut (.I0(GND_net), .I1(n44_adj_4344), .I2(n113_adj_4343), 
            .I3(GND_net), .O(n13343[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5359_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5359_2 (.CI(GND_net), .I0(n44_adj_4344), .I1(n113_adj_4343), 
            .CO(n31431));
    SB_LUT4 add_5234_20_lut (.I0(GND_net), .I1(n11646[17]), .I2(GND_net), 
            .I3(n31430), .O(n11287[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5234_19_lut (.I0(GND_net), .I1(n11646[16]), .I2(GND_net), 
            .I3(n31429), .O(n11287[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_19 (.CI(n31429), .I0(n11646[16]), .I1(GND_net), 
            .CO(n31430));
    SB_LUT4 add_12_25_lut (.I0(GND_net), .I1(n7896[0]), .I2(n7900[0]), 
            .I3(n30739), .O(duty_23__N_3613[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5234_18_lut (.I0(GND_net), .I1(n11646[15]), .I2(GND_net), 
            .I3(n31428), .O(n11287[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_24_lut (.I0(GND_net), .I1(n106[22]), .I2(n155[22]), 
            .I3(n30738), .O(duty_23__N_3613[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(motor_state[18]), 
            .I3(n30894), .O(n28[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_18 (.CI(n31428), .I0(n11646[15]), .I1(GND_net), 
            .CO(n31429));
    SB_LUT4 add_5234_17_lut (.I0(GND_net), .I1(n11646[14]), .I2(GND_net), 
            .I3(n31427), .O(n11287[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_17 (.CI(n31427), .I0(n11646[14]), .I1(GND_net), 
            .CO(n31428));
    SB_LUT4 add_5234_16_lut (.I0(GND_net), .I1(n11646[13]), .I2(n1108), 
            .I3(n31426), .O(n11287[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_16 (.CI(n31426), .I0(n11646[13]), .I1(n1108), .CO(n31427));
    SB_LUT4 add_5234_15_lut (.I0(GND_net), .I1(n11646[12]), .I2(n1035), 
            .I3(n31425), .O(n11287[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_15 (.CI(n31425), .I0(n11646[12]), .I1(n1035), .CO(n31426));
    SB_LUT4 add_5234_14_lut (.I0(GND_net), .I1(n11646[11]), .I2(n962), 
            .I3(n31424), .O(n11287[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_14 (.CI(n31424), .I0(n11646[11]), .I1(n962), .CO(n31425));
    SB_LUT4 i2_4_lut_adj_1514 (.I0(n4_adj_4428), .I1(\Kp[3] ), .I2(n13707[1]), 
            .I3(n28[19]), .O(n13692[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1514.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(n28[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_4429));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[21]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5234_13_lut (.I0(GND_net), .I1(n11646[10]), .I2(n889), 
            .I3(n31423), .O(n11287[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_24 (.CI(n30738), .I0(n106[22]), .I1(n155[22]), .CO(n30739));
    SB_CARRY add_5234_13 (.CI(n31423), .I0(n11646[10]), .I1(n889), .CO(n31424));
    SB_LUT4 i2_4_lut_adj_1515 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(n28[23]), 
            .I3(n28[20]), .O(n12_adj_4431));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1515.LUT_INIT = 16'h9c50;
    SB_LUT4 add_5234_12_lut (.I0(GND_net), .I1(n11646[9]), .I2(n816), 
            .I3(n31422), .O(n11287[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691_adj_4432));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5234_12 (.CI(n31422), .I0(n11646[9]), .I1(n816), .CO(n31423));
    SB_CARRY sub_3_add_2_20 (.CI(n30894), .I0(setpoint[18]), .I1(motor_state[18]), 
            .CO(n30895));
    SB_LUT4 sub_3_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(motor_state[17]), 
            .I3(n30893), .O(n28[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_23_lut (.I0(GND_net), .I1(n106[21]), .I2(n155[21]), 
            .I3(n30737), .O(duty_23__N_3613[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22120_4_lut (.I0(n13692[2]), .I1(\Kp[4] ), .I2(n6_adj_4420), 
            .I3(n28[18]), .O(n8_adj_4433));   // verilog/motorControl.v(34[16:22])
    defparam i22120_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_1516 (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(n28[19]), 
            .I3(n28[21]), .O(n11_adj_4434));   // verilog/motorControl.v(34[16:22])
    defparam i1_4_lut_adj_1516.LUT_INIT = 16'h6ca0;
    SB_LUT4 i22074_4_lut (.I0(n13707[1]), .I1(\Kp[3] ), .I2(n4_adj_4428), 
            .I3(n28[19]), .O(n6_adj_4435));   // verilog/motorControl.v(34[16:22])
    defparam i22074_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 add_5234_11_lut (.I0(GND_net), .I1(n11646[8]), .I2(n743), 
            .I3(n31421), .O(n11287[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_11 (.CI(n31421), .I0(n11646[8]), .I1(n743), .CO(n31422));
    SB_LUT4 i22040_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n28[22]), .I3(n28[21]), 
            .O(n30411));   // verilog/motorControl.v(34[16:22])
    defparam i22040_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_5234_10_lut (.I0(GND_net), .I1(n11646[7]), .I2(n670), 
            .I3(n31420), .O(n11287[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_10 (.CI(n31420), .I0(n11646[7]), .I1(n670), .CO(n31421));
    SB_LUT4 add_5234_9_lut (.I0(GND_net), .I1(n11646[6]), .I2(n597), .I3(n31419), 
            .O(n11287[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_19 (.CI(n30893), .I0(setpoint[17]), .I1(motor_state[17]), 
            .CO(n30894));
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[22]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[23]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_4_lut_adj_1517 (.I0(n6_adj_4435), .I1(n11_adj_4434), .I2(n8_adj_4433), 
            .I3(n12_adj_4431), .O(n18_adj_4437));   // verilog/motorControl.v(34[16:22])
    defparam i8_4_lut_adj_1517.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1518 (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(n28[18]), 
            .I3(n28[22]), .O(n13_adj_4438));   // verilog/motorControl.v(34[16:22])
    defparam i3_4_lut_adj_1518.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut_adj_1519 (.I0(n13_adj_4438), .I1(n18_adj_4437), .I2(n30411), 
            .I3(n4_adj_4439), .O(n37173));   // verilog/motorControl.v(34[16:22])
    defparam i9_4_lut_adj_1519.LUT_INIT = 16'h6996;
    SB_CARRY add_5234_9 (.CI(n31419), .I0(n11646[6]), .I1(n597), .CO(n31420));
    SB_LUT4 add_5234_8_lut (.I0(GND_net), .I1(n11646[5]), .I2(n524), .I3(n31418), 
            .O(n11287[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_8 (.CI(n31418), .I0(n11646[5]), .I1(n524), .CO(n31419));
    SB_LUT4 add_5234_7_lut (.I0(GND_net), .I1(n11646[4]), .I2(n451), .I3(n31417), 
            .O(n11287[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_7 (.CI(n31417), .I0(n11646[4]), .I1(n451), .CO(n31418));
    SB_LUT4 add_5234_6_lut (.I0(GND_net), .I1(n11646[3]), .I2(n378), .I3(n31416), 
            .O(n11287[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_6 (.CI(n31416), .I0(n11646[3]), .I1(n378), .CO(n31417));
    SB_LUT4 add_5234_5_lut (.I0(GND_net), .I1(n11646[2]), .I2(n305), .I3(n31415), 
            .O(n11287[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764_adj_4440));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5234_5 (.CI(n31415), .I0(n11646[2]), .I1(n305), .CO(n31416));
    SB_LUT4 add_5234_4_lut (.I0(GND_net), .I1(n11646[1]), .I2(n232), .I3(n31414), 
            .O(n11287[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_23 (.CI(n30737), .I0(n106[21]), .I1(n155[21]), .CO(n30738));
    SB_LUT4 add_12_22_lut (.I0(GND_net), .I1(n106[20]), .I2(n155[20]), 
            .I3(n30736), .O(duty_23__N_3613[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_4 (.CI(n31414), .I0(n11646[1]), .I1(n232), .CO(n31415));
    SB_LUT4 add_5234_3_lut (.I0(GND_net), .I1(n11646[0]), .I2(n159), .I3(n31413), 
            .O(n11287[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_3 (.CI(n31413), .I0(n11646[0]), .I1(n159), .CO(n31414));
    SB_LUT4 add_5234_2_lut (.I0(GND_net), .I1(n17_adj_4334), .I2(n86), 
            .I3(GND_net), .O(n11287[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5234_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5234_2 (.CI(GND_net), .I0(n17_adj_4334), .I1(n86), .CO(n31413));
    SB_LUT4 add_5252_19_lut (.I0(GND_net), .I1(n11968[16]), .I2(GND_net), 
            .I3(n31412), .O(n11646[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5252_18_lut (.I0(GND_net), .I1(n11968[15]), .I2(GND_net), 
            .I3(n31411), .O(n11646[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_18 (.CI(n31411), .I0(n11968[15]), .I1(GND_net), 
            .CO(n31412));
    SB_LUT4 add_5252_17_lut (.I0(GND_net), .I1(n11968[14]), .I2(GND_net), 
            .I3(n31410), .O(n11646[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_17 (.CI(n31410), .I0(n11968[14]), .I1(GND_net), 
            .CO(n31411));
    SB_LUT4 add_5252_16_lut (.I0(GND_net), .I1(n11968[13]), .I2(n1111), 
            .I3(n31409), .O(n11646[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_16 (.CI(n31409), .I0(n11968[13]), .I1(n1111), .CO(n31410));
    SB_LUT4 add_5252_15_lut (.I0(GND_net), .I1(n11968[12]), .I2(n1038), 
            .I3(n31408), .O(n11646[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_15 (.CI(n31408), .I0(n11968[12]), .I1(n1038), .CO(n31409));
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837_adj_4442));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(motor_state[16]), 
            .I3(n30892), .O(n28[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_18 (.CI(n30892), .I0(setpoint[16]), .I1(motor_state[16]), 
            .CO(n30893));
    SB_LUT4 sub_3_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(motor_state[15]), 
            .I3(n30891), .O(n28[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5252_14_lut (.I0(GND_net), .I1(n11968[11]), .I2(n965), 
            .I3(n31407), .O(n11646[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_14 (.CI(n31407), .I0(n11968[11]), .I1(n965), .CO(n31408));
    SB_LUT4 add_5252_13_lut (.I0(GND_net), .I1(n11968[10]), .I2(n892), 
            .I3(n31406), .O(n11646[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_13 (.CI(n31406), .I0(n11968[10]), .I1(n892), .CO(n31407));
    SB_LUT4 add_5252_12_lut (.I0(GND_net), .I1(n11968[9]), .I2(n819), 
            .I3(n31405), .O(n11646[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_12 (.CI(n31405), .I0(n11968[9]), .I1(n819), .CO(n31406));
    SB_CARRY sub_3_add_2_17 (.CI(n30891), .I0(setpoint[15]), .I1(motor_state[15]), 
            .CO(n30892));
    SB_LUT4 add_5252_11_lut (.I0(GND_net), .I1(n11968[8]), .I2(n746), 
            .I3(n31404), .O(n11646[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_11 (.CI(n31404), .I0(n11968[8]), .I1(n746), .CO(n31405));
    SB_LUT4 add_5252_10_lut (.I0(GND_net), .I1(n11968[7]), .I2(n673), 
            .I3(n31403), .O(n11646[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_10 (.CI(n31403), .I0(n11968[7]), .I1(n673), .CO(n31404));
    SB_LUT4 add_5252_9_lut (.I0(GND_net), .I1(n11968[6]), .I2(n600), .I3(n31402), 
            .O(n11646[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_9 (.CI(n31402), .I0(n11968[6]), .I1(n600), .CO(n31403));
    SB_LUT4 add_5252_8_lut (.I0(GND_net), .I1(n11968[5]), .I2(n527), .I3(n31401), 
            .O(n11646[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(motor_state[14]), 
            .I3(n30890), .O(n28[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_8 (.CI(n31401), .I0(n11968[5]), .I1(n527), .CO(n31402));
    SB_LUT4 add_5252_7_lut (.I0(GND_net), .I1(n11968[4]), .I2(n454), .I3(n31400), 
            .O(n11646[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_7 (.CI(n31400), .I0(n11968[4]), .I1(n454), .CO(n31401));
    SB_CARRY sub_3_add_2_16 (.CI(n30890), .I0(setpoint[14]), .I1(motor_state[14]), 
            .CO(n30891));
    SB_LUT4 sub_3_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(motor_state[13]), 
            .I3(n30889), .O(n28[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_15 (.CI(n30889), .I0(setpoint[13]), .I1(motor_state[13]), 
            .CO(n30890));
    SB_LUT4 sub_3_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(motor_state[12]), 
            .I3(n30888), .O(n28[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5252_6_lut (.I0(GND_net), .I1(n11968[3]), .I2(n381), .I3(n31399), 
            .O(n11646[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_22 (.CI(n30736), .I0(n106[20]), .I1(n155[20]), .CO(n30737));
    SB_CARRY sub_3_add_2_14 (.CI(n30888), .I0(setpoint[12]), .I1(motor_state[12]), 
            .CO(n30889));
    SB_LUT4 sub_3_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(motor_state[11]), 
            .I3(n30887), .O(n28[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_21_lut (.I0(GND_net), .I1(n106[19]), .I2(n155[19]), 
            .I3(n30735), .O(duty_23__N_3613[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_13 (.CI(n30887), .I0(setpoint[11]), .I1(motor_state[11]), 
            .CO(n30888));
    SB_CARRY add_12_21 (.CI(n30735), .I0(n106[19]), .I1(n155[19]), .CO(n30736));
    SB_LUT4 add_12_20_lut (.I0(GND_net), .I1(n106[18]), .I2(n155[18]), 
            .I3(n30734), .O(duty_23__N_3613[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(motor_state[10]), 
            .I3(n30886), .O(n28[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_6 (.CI(n31399), .I0(n11968[3]), .I1(n381), .CO(n31400));
    SB_LUT4 add_5252_5_lut (.I0(GND_net), .I1(n11968[2]), .I2(n308), .I3(n31398), 
            .O(n11646[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_12 (.CI(n30886), .I0(setpoint[10]), .I1(motor_state[10]), 
            .CO(n30887));
    SB_CARRY add_12_20 (.CI(n30734), .I0(n106[18]), .I1(n155[18]), .CO(n30735));
    SB_CARRY add_5252_5 (.CI(n31398), .I0(n11968[2]), .I1(n308), .CO(n31399));
    SB_LUT4 add_5252_4_lut (.I0(GND_net), .I1(n11968[1]), .I2(n235), .I3(n31397), 
            .O(n11646[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5252_4 (.CI(n31397), .I0(n11968[1]), .I1(n235), .CO(n31398));
    SB_LUT4 add_5252_3_lut (.I0(GND_net), .I1(n11968[0]), .I2(n162), .I3(n31396), 
            .O(n11646[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_3 (.CI(n31396), .I0(n11968[0]), .I1(n162), .CO(n31397));
    SB_LUT4 add_5252_2_lut (.I0(GND_net), .I1(n20_adj_4329), .I2(n89), 
            .I3(GND_net), .O(n11646[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5252_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5252_2 (.CI(GND_net), .I0(n20_adj_4329), .I1(n89), .CO(n31396));
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323_adj_4444));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i18684_2_lut (.I0(n28[0]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[0]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i18684_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5338_13_lut (.I0(GND_net), .I1(n13223[10]), .I2(n910_adj_4445), 
            .I3(n30772), .O(n13080[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(motor_state[9]), 
            .I3(n30885), .O(n28[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_19_lut (.I0(GND_net), .I1(n106[17]), .I2(n155[17]), 
            .I3(n30733), .O(duty_23__N_3613[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_11 (.CI(n30885), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n30886));
    SB_LUT4 sub_3_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(motor_state[8]), 
            .I3(n30884), .O(n28[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5338_12_lut (.I0(GND_net), .I1(n13223[9]), .I2(n837_adj_4442), 
            .I3(n30771), .O(n13080[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_10 (.CI(n30884), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n30885));
    SB_CARRY add_5338_12 (.CI(n30771), .I0(n13223[9]), .I1(n837_adj_4442), 
            .CO(n30772));
    SB_LUT4 sub_3_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(motor_state[7]), 
            .I3(n30883), .O(n28[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_9 (.CI(n30883), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n30884));
    SB_LUT4 sub_3_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(motor_state[6]), 
            .I3(n30882), .O(n28[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_19 (.CI(n30733), .I0(n106[17]), .I1(n155[17]), .CO(n30734));
    SB_CARRY sub_3_add_2_8 (.CI(n30882), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n30883));
    SB_LUT4 sub_3_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(motor_state[5]), 
            .I3(n30881), .O(n28[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_7 (.CI(n30881), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n30882));
    SB_LUT4 sub_3_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(motor_state[4]), 
            .I3(n30880), .O(n28[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5338_11_lut (.I0(GND_net), .I1(n13223[8]), .I2(n764_adj_4440), 
            .I3(n30770), .O(n13080[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_18_lut (.I0(GND_net), .I1(n106[16]), .I2(n155[16]), 
            .I3(n30732), .O(duty_23__N_3613[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_6 (.CI(n30880), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n30881));
    SB_LUT4 sub_3_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(motor_state[3]), 
            .I3(n30879), .O(n28[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5338_11 (.CI(n30770), .I0(n13223[8]), .I1(n764_adj_4440), 
            .CO(n30771));
    SB_CARRY sub_3_add_2_5 (.CI(n30879), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n30880));
    SB_CARRY add_12_18 (.CI(n30732), .I0(n106[16]), .I1(n155[16]), .CO(n30733));
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[23]), 
            .I3(n30945), .O(n257[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_17_lut (.I0(GND_net), .I1(n106[15]), .I2(n155[15]), 
            .I3(n30731), .O(duty_23__N_3613[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[22]), 
            .I3(n30944), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(motor_state[2]), 
            .I3(n30878), .O(n28[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5338_10_lut (.I0(GND_net), .I1(n13223[7]), .I2(n691_adj_4432), 
            .I3(n30769), .O(n13080[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_4 (.CI(n30878), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n30879));
    SB_CARRY unary_minus_16_add_3_24 (.CI(n30944), .I0(GND_net), .I1(n1_adj_4704[22]), 
            .CO(n30945));
    SB_CARRY add_12_17 (.CI(n30731), .I0(n106[15]), .I1(n155[15]), .CO(n30732));
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[21]), 
            .I3(n30943), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(motor_state[1]), 
            .I3(n30877), .O(n28[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_3 (.CI(n30877), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n30878));
    SB_LUT4 sub_3_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(motor_state[0]), 
            .I3(VCC_net), .O(n28[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_16_lut (.I0(GND_net), .I1(n106[14]), .I2(n155[14]), 
            .I3(n30730), .O(duty_23__N_3613[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n30877));
    SB_CARRY add_5338_10 (.CI(n30769), .I0(n13223[7]), .I1(n691_adj_4432), 
            .CO(n30770));
    SB_LUT4 add_5338_9_lut (.I0(GND_net), .I1(n13223[6]), .I2(n618_adj_4427), 
            .I3(n30768), .O(n13080[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_16 (.CI(n30730), .I0(n106[14]), .I1(n155[14]), .CO(n30731));
    SB_LUT4 add_723_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n3141[23]), .I3(n30816), .O(\PID_CONTROLLER.integral_23__N_3513 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_12_15_lut (.I0(GND_net), .I1(n106[13]), .I2(n155[13]), 
            .I3(n30729), .O(duty_23__N_3613[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_723_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n3141[22]), .I3(n30815), .O(\PID_CONTROLLER.integral_23__N_3513 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5383_8_lut (.I0(GND_net), .I1(n13633[5]), .I2(n560_adj_4389), 
            .I3(n31005), .O(n13585[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n30943), .I0(GND_net), .I1(n1_adj_4704[21]), 
            .CO(n30944));
    SB_CARRY add_723_24 (.CI(n30815), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n3141[22]), .CO(n30816));
    SB_CARRY add_5338_9 (.CI(n30768), .I0(n13223[6]), .I1(n618_adj_4427), 
            .CO(n30769));
    SB_CARRY add_12_15 (.CI(n30729), .I0(n106[13]), .I1(n155[13]), .CO(n30730));
    SB_LUT4 add_5383_7_lut (.I0(GND_net), .I1(n13633[4]), .I2(n487_adj_4388), 
            .I3(n31004), .O(n13585[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[20]), 
            .I3(n30942), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396_adj_4451));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5383_7 (.CI(n31004), .I0(n13633[4]), .I1(n487_adj_4388), 
            .CO(n31005));
    SB_CARRY unary_minus_16_add_3_22 (.CI(n30942), .I0(GND_net), .I1(n1_adj_4704[20]), 
            .CO(n30943));
    SB_LUT4 add_723_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n3141[21]), .I3(n30814), .O(\PID_CONTROLLER.integral_23__N_3513 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5338_8_lut (.I0(GND_net), .I1(n13223[5]), .I2(n545_adj_4385), 
            .I3(n30767), .O(n13080[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty_23__N_3613[20]), .I1(n257[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4452));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty_23__N_3613[19]), .I1(n257[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4454));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty_23__N_3613[22]), .I1(n257[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4455));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_11_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n155[0]));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n106[0]));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[19]), 
            .I3(n30941), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(n28[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910_adj_4445));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19128_2_lut (.I0(n28[1]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[1]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5167_7_lut (.I0(GND_net), .I1(n37896), .I2(n490), .I3(n32267), 
            .O(n9978[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5167_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5167_6_lut (.I0(GND_net), .I1(n9986[3]), .I2(n417), .I3(n32266), 
            .O(n9978[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5167_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5167_6 (.CI(n32266), .I0(n9986[3]), .I1(n417), .CO(n32267));
    SB_LUT4 add_5167_5_lut (.I0(GND_net), .I1(n9986[2]), .I2(n344), .I3(n32265), 
            .O(n9978[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5167_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5167_5 (.CI(n32265), .I0(n9986[2]), .I1(n344), .CO(n32266));
    SB_LUT4 add_5167_4_lut (.I0(GND_net), .I1(n9986[1]), .I2(n271), .I3(n32264), 
            .O(n9978[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5167_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5167_4 (.CI(n32264), .I0(n9986[1]), .I1(n271), .CO(n32265));
    SB_LUT4 add_5167_3_lut (.I0(GND_net), .I1(n9986[0]), .I2(n198_adj_4368), 
            .I3(n32263), .O(n9978[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5167_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5167_3 (.CI(n32263), .I0(n9986[0]), .I1(n198_adj_4368), 
            .CO(n32264));
    SB_LUT4 add_5167_2_lut (.I0(GND_net), .I1(n56_adj_4366), .I2(n125_adj_4365), 
            .I3(GND_net), .O(n9978[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5167_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i30593_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40620));   // verilog/motorControl.v(29[14] 48[8])
    defparam i30593_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5167_2 (.CI(GND_net), .I0(n56_adj_4366), .I1(n125_adj_4365), 
            .CO(n32263));
    SB_LUT4 add_5166_8_lut (.I0(GND_net), .I1(n9978[5]), .I2(n560), .I3(n32262), 
            .O(n9969[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5166_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5166_7_lut (.I0(GND_net), .I1(n9978[4]), .I2(n487), .I3(n32261), 
            .O(n9969[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5166_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5166_7 (.CI(n32261), .I0(n9978[4]), .I1(n487), .CO(n32262));
    SB_LUT4 add_5166_6_lut (.I0(GND_net), .I1(n9978[3]), .I2(n414_adj_4349), 
            .I3(n32260), .O(n9969[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5166_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5166_6 (.CI(n32260), .I0(n9978[3]), .I1(n414_adj_4349), 
            .CO(n32261));
    SB_LUT4 add_5166_5_lut (.I0(GND_net), .I1(n9978[2]), .I2(n341_adj_4348), 
            .I3(n32259), .O(n9969[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5166_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5166_5 (.CI(n32259), .I0(n9978[2]), .I1(n341_adj_4348), 
            .CO(n32260));
    SB_LUT4 add_5383_6_lut (.I0(GND_net), .I1(n13633[3]), .I2(n414), .I3(n31003), 
            .O(n13585[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5383_6 (.CI(n31003), .I0(n13633[3]), .I1(n414), .CO(n31004));
    SB_CARRY unary_minus_16_add_3_21 (.CI(n30941), .I0(GND_net), .I1(n1_adj_4704[19]), 
            .CO(n30942));
    SB_LUT4 add_5383_5_lut (.I0(GND_net), .I1(n13633[2]), .I2(n341), .I3(n31002), 
            .O(n13585[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5383_5 (.CI(n31002), .I0(n13633[2]), .I1(n341), .CO(n31003));
    SB_LUT4 add_5383_4_lut (.I0(GND_net), .I1(n13633[1]), .I2(n268_adj_4346), 
            .I3(n31001), .O(n13585[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5383_4 (.CI(n31001), .I0(n13633[1]), .I1(n268_adj_4346), 
            .CO(n31002));
    SB_LUT4 add_5166_4_lut (.I0(GND_net), .I1(n9978[1]), .I2(n268), .I3(n32258), 
            .O(n9969[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5166_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5166_4 (.CI(n32258), .I0(n9978[1]), .I1(n268), .CO(n32259));
    SB_LUT4 add_5166_3_lut (.I0(GND_net), .I1(n9978[0]), .I2(n195_adj_4342), 
            .I3(n32257), .O(n9969[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5166_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5166_3 (.CI(n32257), .I0(n9978[0]), .I1(n195_adj_4342), 
            .CO(n32258));
    SB_LUT4 add_5166_2_lut (.I0(GND_net), .I1(n53_adj_4341), .I2(n122_adj_4340), 
            .I3(GND_net), .O(n9969[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5166_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5383_3_lut (.I0(GND_net), .I1(n13633[0]), .I2(n195), .I3(n31000), 
            .O(n13585[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5166_2 (.CI(GND_net), .I0(n53_adj_4341), .I1(n122_adj_4340), 
            .CO(n32257));
    SB_LUT4 add_5165_9_lut (.I0(GND_net), .I1(n9969[6]), .I2(n630), .I3(n32256), 
            .O(n9959[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5165_8_lut (.I0(GND_net), .I1(n9969[5]), .I2(n557), .I3(n32255), 
            .O(n9959[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_8 (.CI(n32255), .I0(n9969[5]), .I1(n557), .CO(n32256));
    SB_LUT4 add_5165_7_lut (.I0(GND_net), .I1(n9969[4]), .I2(n484), .I3(n32254), 
            .O(n9959[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_7 (.CI(n32254), .I0(n9969[4]), .I1(n484), .CO(n32255));
    SB_LUT4 add_5165_6_lut (.I0(GND_net), .I1(n9969[3]), .I2(n411), .I3(n32253), 
            .O(n9959[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_6 (.CI(n32253), .I0(n9969[3]), .I1(n411), .CO(n32254));
    SB_LUT4 add_5165_5_lut (.I0(GND_net), .I1(n9969[2]), .I2(n338), .I3(n32252), 
            .O(n9959[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_5 (.CI(n32252), .I0(n9969[2]), .I1(n338), .CO(n32253));
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[18]), 
            .I3(n30940), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5165_4_lut (.I0(GND_net), .I1(n9969[1]), .I2(n265), .I3(n32251), 
            .O(n9959[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_4 (.CI(n32251), .I0(n9969[1]), .I1(n265), .CO(n32252));
    SB_CARRY unary_minus_16_add_3_20 (.CI(n30940), .I0(GND_net), .I1(n1_adj_4704[18]), 
            .CO(n30941));
    SB_LUT4 add_5165_3_lut (.I0(GND_net), .I1(n9969[0]), .I2(n192), .I3(n32250), 
            .O(n9959[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_3 (.CI(n32250), .I0(n9969[0]), .I1(n192), .CO(n32251));
    SB_LUT4 add_5165_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n9959[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5165_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5165_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n32250));
    SB_CARRY add_5383_3 (.CI(n31000), .I0(n13633[0]), .I1(n195), .CO(n31001));
    SB_CARRY add_5338_8 (.CI(n30767), .I0(n13223[5]), .I1(n545_adj_4385), 
            .CO(n30768));
    SB_LUT4 add_5164_10_lut (.I0(GND_net), .I1(n9959[7]), .I2(n700), .I3(n32249), 
            .O(n9948[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5164_9_lut (.I0(GND_net), .I1(n9959[6]), .I2(n627), .I3(n32248), 
            .O(n9948[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5164_9 (.CI(n32248), .I0(n9959[6]), .I1(n627), .CO(n32249));
    SB_LUT4 add_5164_8_lut (.I0(GND_net), .I1(n9959[5]), .I2(n554), .I3(n32247), 
            .O(n9948[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5164_8 (.CI(n32247), .I0(n9959[5]), .I1(n554), .CO(n32248));
    SB_LUT4 add_5164_7_lut (.I0(GND_net), .I1(n9959[4]), .I2(n481_adj_4331), 
            .I3(n32246), .O(n9948[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_723_23 (.CI(n30814), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n3141[21]), .CO(n30815));
    SB_CARRY add_5164_7 (.CI(n32246), .I0(n9959[4]), .I1(n481_adj_4331), 
            .CO(n32247));
    SB_LUT4 add_5338_7_lut (.I0(GND_net), .I1(n13223[4]), .I2(n472_adj_4330), 
            .I3(n30766), .O(n13080[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5164_6_lut (.I0(GND_net), .I1(n9959[3]), .I2(n408_adj_4327), 
            .I3(n32245), .O(n9948[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5164_6 (.CI(n32245), .I0(n9959[3]), .I1(n408_adj_4327), 
            .CO(n32246));
    SB_LUT4 add_5164_5_lut (.I0(GND_net), .I1(n9959[2]), .I2(n335_adj_4326), 
            .I3(n32244), .O(n9948[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_14_lut (.I0(GND_net), .I1(n106[12]), .I2(n155[12]), 
            .I3(n30728), .O(duty_23__N_3613[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5164_5 (.CI(n32244), .I0(n9959[2]), .I1(n335_adj_4326), 
            .CO(n32245));
    SB_LUT4 add_5164_4_lut (.I0(GND_net), .I1(n9959[1]), .I2(n262_adj_4325), 
            .I3(n32243), .O(n9948[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5164_4 (.CI(n32243), .I0(n9959[1]), .I1(n262_adj_4325), 
            .CO(n32244));
    SB_LUT4 add_5164_3_lut (.I0(GND_net), .I1(n9959[0]), .I2(n189_adj_4324), 
            .I3(n32242), .O(n9948[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5164_3 (.CI(n32242), .I0(n9959[0]), .I1(n189_adj_4324), 
            .CO(n32243));
    SB_LUT4 add_5164_2_lut (.I0(GND_net), .I1(n47_adj_4323), .I2(n116_adj_4322), 
            .I3(GND_net), .O(n9948[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5164_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5164_2 (.CI(GND_net), .I0(n47_adj_4323), .I1(n116_adj_4322), 
            .CO(n32242));
    SB_LUT4 add_5163_11_lut (.I0(GND_net), .I1(n9948[8]), .I2(n770), .I3(n32241), 
            .O(n9936[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5163_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5383_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n13585[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5383_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5163_10_lut (.I0(GND_net), .I1(n9948[7]), .I2(n697), .I3(n32240), 
            .O(n9936[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5163_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5163_10 (.CI(n32240), .I0(n9948[7]), .I1(n697), .CO(n32241));
    SB_LUT4 add_5163_9_lut (.I0(GND_net), .I1(n9948[6]), .I2(n624), .I3(n32239), 
            .O(n9936[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5163_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5163_9 (.CI(n32239), .I0(n9948[6]), .I1(n624), .CO(n32240));
    SB_LUT4 add_5163_8_lut (.I0(GND_net), .I1(n9948[5]), .I2(n551), .I3(n32238), 
            .O(n9936[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5163_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[17]), 
            .I3(n30939), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_19 (.CI(n30939), .I0(GND_net), .I1(n1_adj_4704[17]), 
            .CO(n30940));
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[16]), 
            .I3(n30938), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5163_8 (.CI(n32238), .I0(n9948[5]), .I1(n551), .CO(n32239));
    SB_LUT4 add_5163_7_lut (.I0(GND_net), .I1(n9948[4]), .I2(n478), .I3(n32237), 
            .O(n9936[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5163_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5163_7 (.CI(n32237), .I0(n9948[4]), .I1(n478), .CO(n32238));
    SB_LUT4 add_5163_6_lut (.I0(GND_net), .I1(n9948[3]), .I2(n405), .I3(n32236), 
            .O(n9936[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5163_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5163_6 (.CI(n32236), .I0(n9948[3]), .I1(n405), .CO(n32237));
    SB_LUT4 add_5163_5_lut (.I0(GND_net), .I1(n9948[2]), .I2(n332), .I3(n32235), 
            .O(n9936[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5163_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5163_5 (.CI(n32235), .I0(n9948[2]), .I1(n332), .CO(n32236));
    SB_LUT4 add_5163_4_lut (.I0(GND_net), .I1(n9948[1]), .I2(n259), .I3(n32234), 
            .O(n9936[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5163_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5163_4 (.CI(n32234), .I0(n9948[1]), .I1(n259), .CO(n32235));
    SB_LUT4 add_5163_3_lut (.I0(GND_net), .I1(n9948[0]), .I2(n186), .I3(n32233), 
            .O(n9936[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5163_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5163_3 (.CI(n32233), .I0(n9948[0]), .I1(n186), .CO(n32234));
    SB_LUT4 add_5163_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n9936[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5163_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5163_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n32233));
    SB_LUT4 add_5162_12_lut (.I0(GND_net), .I1(n9936[9]), .I2(n840), .I3(n32232), 
            .O(n9923[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5162_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5162_11_lut (.I0(GND_net), .I1(n9936[8]), .I2(n767), .I3(n32231), 
            .O(n9923[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5162_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5162_11 (.CI(n32231), .I0(n9936[8]), .I1(n767), .CO(n32232));
    SB_LUT4 add_5162_10_lut (.I0(GND_net), .I1(n9936[7]), .I2(n694), .I3(n32230), 
            .O(n9923[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5162_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5162_10 (.CI(n32230), .I0(n9936[7]), .I1(n694), .CO(n32231));
    SB_LUT4 add_5162_9_lut (.I0(GND_net), .I1(n9936[6]), .I2(n621), .I3(n32229), 
            .O(n9923[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5162_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5162_9 (.CI(n32229), .I0(n9936[6]), .I1(n621), .CO(n32230));
    SB_LUT4 add_5162_8_lut (.I0(GND_net), .I1(n9936[5]), .I2(n548), .I3(n32228), 
            .O(n9923[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5162_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty_23__N_3613[18]), .I1(n257[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4458));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5162_8 (.CI(n32228), .I0(n9936[5]), .I1(n548), .CO(n32229));
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty_23__N_3613[14]), .I1(n257[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4459));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty_23__N_3613[15]), .I1(n257[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4460));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty_23__N_3613[21]), .I1(n257[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4461));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty_23__N_3613[11]), .I1(n257[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4462));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty_23__N_3613[12]), .I1(n257[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4463));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty_23__N_3613[17]), .I1(n257[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4464));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty_23__N_3613[5]), .I1(n257[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4465));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty_23__N_3613[6]), .I1(n257[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4466));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty_23__N_3613[7]), .I1(n257[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4467));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty_23__N_3613[13]), .I1(n257[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4469));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty_23__N_3613[16]), .I1(n257[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4470));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty_23__N_3613[4]), .I1(n257[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4471));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty_23__N_3613[8]), .I1(n257[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4472));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty_23__N_3613[9]), .I1(n257[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4473));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty_23__N_3613[10]), .I1(n257[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4475));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29341_4_lut (.I0(n21_adj_4475), .I1(n19_adj_4473), .I2(n17_adj_4472), 
            .I3(n9_adj_4471), .O(n39369));
    defparam i29341_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29333_4_lut (.I0(n27_adj_4469), .I1(n15_adj_4467), .I2(n13_adj_4466), 
            .I3(n11_adj_4465), .O(n39361));
    defparam i29333_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_4470), 
            .I3(GND_net), .O(n12_adj_4476));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_4466), 
            .I3(GND_net), .O(n10_adj_4477));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_4476), .I1(n257[17]), .I2(n35_adj_4464), 
            .I3(GND_net), .O(n30_adj_4478));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5162_7_lut (.I0(GND_net), .I1(n9936[4]), .I2(n475), .I3(n32227), 
            .O(n9923[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5162_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29621_4_lut (.I0(n13_adj_4466), .I1(n11_adj_4465), .I2(n9_adj_4471), 
            .I3(n39379), .O(n39650));
    defparam i29621_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_5162_7 (.CI(n32227), .I0(n9936[4]), .I1(n475), .CO(n32228));
    SB_LUT4 i29617_4_lut (.I0(n19_adj_4473), .I1(n17_adj_4472), .I2(n15_adj_4467), 
            .I3(n39650), .O(n39646));
    defparam i29617_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i29943_4_lut (.I0(n25_adj_4463), .I1(n23_adj_4462), .I2(n21_adj_4475), 
            .I3(n39646), .O(n39972));
    defparam i29943_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i29774_4_lut (.I0(n31_adj_4460), .I1(n29_adj_4459), .I2(n27_adj_4469), 
            .I3(n39972), .O(n39803));
    defparam i29774_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i30009_4_lut (.I0(n37_adj_4458), .I1(n35_adj_4464), .I2(n33_adj_4470), 
            .I3(n39803), .O(n40038));
    defparam i30009_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_4461), 
            .I3(GND_net), .O(n16_adj_4479));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29921_3_lut (.I0(n6_adj_4480), .I1(n257[10]), .I2(n21_adj_4475), 
            .I3(GND_net), .O(n39950));   // verilog/motorControl.v(38[19:35])
    defparam i29921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29922_3_lut (.I0(n39950), .I1(n257[11]), .I2(n23_adj_4462), 
            .I3(GND_net), .O(n39951));   // verilog/motorControl.v(38[19:35])
    defparam i29922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_4472), 
            .I3(GND_net), .O(n8_adj_4481));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_4479), .I1(n257[22]), .I2(n45_adj_4455), 
            .I3(GND_net), .O(n24_adj_4482));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29319_4_lut (.I0(n43_adj_4461), .I1(n25_adj_4463), .I2(n23_adj_4462), 
            .I3(n39369), .O(n39347));
    defparam i29319_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29828_4_lut (.I0(n24_adj_4482), .I1(n8_adj_4481), .I2(n45_adj_4455), 
            .I3(n39345), .O(n39857));   // verilog/motorControl.v(38[19:35])
    defparam i29828_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29889_3_lut (.I0(n39951), .I1(n257[12]), .I2(n25_adj_4463), 
            .I3(GND_net), .O(n39918));   // verilog/motorControl.v(38[19:35])
    defparam i29889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_4_lut (.I0(duty_23__N_3613[0]), .I1(n257[1]), 
            .I2(duty_23__N_3613[1]), .I3(n257[0]), .O(n4_adj_4483));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i29919_3_lut (.I0(n4_adj_4483), .I1(n257[13]), .I2(n27_adj_4469), 
            .I3(GND_net), .O(n39948));   // verilog/motorControl.v(38[19:35])
    defparam i29919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29920_3_lut (.I0(n39948), .I1(n257[14]), .I2(n29_adj_4459), 
            .I3(GND_net), .O(n39949));   // verilog/motorControl.v(38[19:35])
    defparam i29920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29329_4_lut (.I0(n33_adj_4470), .I1(n31_adj_4460), .I2(n29_adj_4459), 
            .I3(n39361), .O(n39357));
    defparam i29329_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30023_4_lut (.I0(n30_adj_4478), .I1(n10_adj_4477), .I2(n35_adj_4464), 
            .I3(n39355), .O(n40052));   // verilog/motorControl.v(38[19:35])
    defparam i30023_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29891_3_lut (.I0(n39949), .I1(n257[15]), .I2(n31_adj_4460), 
            .I3(GND_net), .O(n39920));   // verilog/motorControl.v(38[19:35])
    defparam i29891_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30074_4_lut (.I0(n39920), .I1(n40052), .I2(n35_adj_4464), 
            .I3(n39357), .O(n40103));   // verilog/motorControl.v(38[19:35])
    defparam i30074_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30075_3_lut (.I0(n40103), .I1(n257[18]), .I2(n37_adj_4458), 
            .I3(GND_net), .O(n40104));   // verilog/motorControl.v(38[19:35])
    defparam i30075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30050_3_lut (.I0(n40104), .I1(n257[19]), .I2(n39_adj_4454), 
            .I3(GND_net), .O(n40079));   // verilog/motorControl.v(38[19:35])
    defparam i30050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29321_4_lut (.I0(n43_adj_4461), .I1(n41_adj_4452), .I2(n39_adj_4454), 
            .I3(n40038), .O(n39349));
    defparam i29321_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29987_4_lut (.I0(n39918), .I1(n39857), .I2(n45_adj_4455), 
            .I3(n39347), .O(n40016));   // verilog/motorControl.v(38[19:35])
    defparam i29987_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30044_3_lut (.I0(n40079), .I1(n257[20]), .I2(n41_adj_4452), 
            .I3(GND_net), .O(n40_adj_4484));   // verilog/motorControl.v(38[19:35])
    defparam i30044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29989_4_lut (.I0(n40_adj_4484), .I1(n40016), .I2(n45_adj_4455), 
            .I3(n39349), .O(n40018));   // verilog/motorControl.v(38[19:35])
    defparam i29989_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i29990_3_lut (.I0(n40018), .I1(duty_23__N_3613[23]), .I2(n257[23]), 
            .I3(GND_net), .O(n256));   // verilog/motorControl.v(38[19:35])
    defparam i29990_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5162_6_lut (.I0(GND_net), .I1(n9936[3]), .I2(n402), .I3(n32226), 
            .O(n9923[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5162_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5162_6 (.CI(n32226), .I0(n9936[3]), .I1(n402), .CO(n32227));
    SB_LUT4 add_5162_5_lut (.I0(GND_net), .I1(n9936[2]), .I2(n329), .I3(n32225), 
            .O(n9923[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5162_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5162_5 (.CI(n32225), .I0(n9936[2]), .I1(n329), .CO(n32226));
    SB_LUT4 add_5162_4_lut (.I0(GND_net), .I1(n9936[1]), .I2(n256_adj_4307), 
            .I3(n32224), .O(n9923[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5162_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5162_4 (.CI(n32224), .I0(n9936[1]), .I1(n256_adj_4307), 
            .CO(n32225));
    SB_LUT4 add_5162_3_lut (.I0(GND_net), .I1(n9936[0]), .I2(n183), .I3(n32223), 
            .O(n9923[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5162_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5162_3 (.CI(n32223), .I0(n9936[0]), .I1(n183), .CO(n32224));
    SB_LUT4 add_5162_2_lut (.I0(GND_net), .I1(n41), .I2(n110), .I3(GND_net), 
            .O(n9923[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5162_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5162_2 (.CI(GND_net), .I0(n41), .I1(n110), .CO(n32223));
    SB_LUT4 add_5161_13_lut (.I0(GND_net), .I1(n9923[10]), .I2(n910), 
            .I3(n32222), .O(n9909[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5161_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5161_12_lut (.I0(GND_net), .I1(n9923[9]), .I2(n837), .I3(n32221), 
            .O(n9909[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5161_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5161_12 (.CI(n32221), .I0(n9923[9]), .I1(n837), .CO(n32222));
    SB_LUT4 add_5161_11_lut (.I0(GND_net), .I1(n9923[8]), .I2(n764), .I3(n32220), 
            .O(n9909[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5161_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5161_11 (.CI(n32220), .I0(n9923[8]), .I1(n764), .CO(n32221));
    SB_LUT4 add_5161_10_lut (.I0(GND_net), .I1(n9923[7]), .I2(n691), .I3(n32219), 
            .O(n9909[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5161_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5161_10 (.CI(n32219), .I0(n9923[7]), .I1(n691), .CO(n32220));
    SB_LUT4 add_5161_9_lut (.I0(GND_net), .I1(n9923[6]), .I2(n618), .I3(n32218), 
            .O(n9909[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5161_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5161_9 (.CI(n32218), .I0(n9923[6]), .I1(n618), .CO(n32219));
    SB_LUT4 add_5161_8_lut (.I0(GND_net), .I1(n9923[5]), .I2(n545), .I3(n32217), 
            .O(n9909[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5161_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5161_8 (.CI(n32217), .I0(n9923[5]), .I1(n545), .CO(n32218));
    SB_LUT4 add_5161_7_lut (.I0(GND_net), .I1(n9923[4]), .I2(n472), .I3(n32216), 
            .O(n9909[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5161_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5161_7 (.CI(n32216), .I0(n9923[4]), .I1(n472), .CO(n32217));
    SB_LUT4 add_5161_6_lut (.I0(GND_net), .I1(n9923[3]), .I2(n399_adj_4304), 
            .I3(n32215), .O(n9909[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5161_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5161_6 (.CI(n32215), .I0(n9923[3]), .I1(n399_adj_4304), 
            .CO(n32216));
    SB_LUT4 add_5161_5_lut (.I0(GND_net), .I1(n9923[2]), .I2(n326_adj_4303), 
            .I3(n32214), .O(n9909[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5161_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5161_5 (.CI(n32214), .I0(n9923[2]), .I1(n326_adj_4303), 
            .CO(n32215));
    SB_LUT4 duty_23__I_831_i39_2_lut (.I0(PWMLimit[19]), .I1(duty_23__N_3613[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4485));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5161_4_lut (.I0(GND_net), .I1(n9923[1]), .I2(n253_adj_4302), 
            .I3(n32213), .O(n9909[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5161_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i41_2_lut (.I0(PWMLimit[20]), .I1(duty_23__N_3613[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4486));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i41_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5161_4 (.CI(n32213), .I0(n9923[1]), .I1(n253_adj_4302), 
            .CO(n32214));
    SB_LUT4 duty_23__I_831_i45_2_lut (.I0(PWMLimit[22]), .I1(duty_23__N_3613[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4487));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5161_3_lut (.I0(GND_net), .I1(n9923[0]), .I2(n180_adj_4301), 
            .I3(n32212), .O(n9909[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5161_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i43_2_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3613[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4488));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i43_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5161_3 (.CI(n32212), .I0(n9923[0]), .I1(n180_adj_4301), 
            .CO(n32213));
    SB_LUT4 add_5161_2_lut (.I0(GND_net), .I1(n38_adj_4300), .I2(n107_adj_4299), 
            .I3(GND_net), .O(n9909[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5161_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_723_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n3141[20]), .I3(n30813), .O(\PID_CONTROLLER.integral_23__N_3513 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_723_22 (.CI(n30813), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n3141[20]), .CO(n30814));
    SB_LUT4 duty_23__I_831_i37_2_lut (.I0(PWMLimit[18]), .I1(duty_23__N_3613[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4489));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5161_2 (.CI(GND_net), .I0(n38_adj_4300), .I1(n107_adj_4299), 
            .CO(n32212));
    SB_LUT4 duty_23__I_831_i29_2_lut (.I0(PWMLimit[14]), .I1(duty_23__N_3613[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4490));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i31_2_lut (.I0(PWMLimit[15]), .I1(duty_23__N_3613[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4491));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i23_2_lut (.I0(PWMLimit[11]), .I1(duty_23__N_3613[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4492));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i25_2_lut (.I0(PWMLimit[12]), .I1(duty_23__N_3613[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4493));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i35_2_lut (.I0(PWMLimit[17]), .I1(duty_23__N_3613[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4494));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i33_2_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3613[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4495));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i11_2_lut (.I0(PWMLimit[5]), .I1(duty_23__N_3613[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4496));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i13_2_lut (.I0(PWMLimit[6]), .I1(duty_23__N_3613[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4497));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5160_14_lut (.I0(GND_net), .I1(n9909[11]), .I2(n980), 
            .I3(n32211), .O(n9894[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5160_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i15_2_lut (.I0(PWMLimit[7]), .I1(duty_23__N_3613[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4498));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i27_2_lut (.I0(PWMLimit[13]), .I1(duty_23__N_3613[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4499));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i9_2_lut (.I0(PWMLimit[4]), .I1(duty_23__N_3613[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4500));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i17_2_lut (.I0(PWMLimit[8]), .I1(duty_23__N_3613[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4501));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_5160_13_lut (.I0(GND_net), .I1(n9909[10]), .I2(n907), 
            .I3(n32210), .O(n9894[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5160_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5160_13 (.CI(n32210), .I0(n9909[10]), .I1(n907), .CO(n32211));
    SB_LUT4 duty_23__I_831_i19_2_lut (.I0(PWMLimit[9]), .I1(duty_23__N_3613[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4502));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_831_i21_2_lut (.I0(PWMLimit[10]), .I1(duty_23__N_3613[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4503));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i29379_4_lut (.I0(n21_adj_4503), .I1(n19_adj_4502), .I2(n17_adj_4501), 
            .I3(n9_adj_4500), .O(n39407));
    defparam i29379_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29371_4_lut (.I0(n27_adj_4499), .I1(n15_adj_4498), .I2(n13_adj_4497), 
            .I3(n11_adj_4496), .O(n39399));
    defparam i29371_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_831_i12_3_lut (.I0(duty_23__N_3613[7]), .I1(duty_23__N_3613[16]), 
            .I2(n33_adj_4495), .I3(GND_net), .O(n12_adj_4504));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5160_12_lut (.I0(GND_net), .I1(n9909[9]), .I2(n834), .I3(n32209), 
            .O(n9894[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5160_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i10_3_lut (.I0(duty_23__N_3613[5]), .I1(duty_23__N_3613[6]), 
            .I2(n13_adj_4497), .I3(GND_net), .O(n10_adj_4505));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_831_i30_3_lut (.I0(n12_adj_4504), .I1(duty_23__N_3613[17]), 
            .I2(n35_adj_4494), .I3(GND_net), .O(n30_adj_4506));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3489[1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 i29654_4_lut (.I0(n13_adj_4497), .I1(n11_adj_4496), .I2(n9_adj_4500), 
            .I3(n39417), .O(n39683));
    defparam i29654_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_5160_12 (.CI(n32209), .I0(n9909[9]), .I1(n834), .CO(n32210));
    SB_LUT4 i29650_4_lut (.I0(n19_adj_4502), .I1(n17_adj_4501), .I2(n15_adj_4498), 
            .I3(n39683), .O(n39679));
    defparam i29650_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i29951_4_lut (.I0(n25_adj_4493), .I1(n23_adj_4492), .I2(n21_adj_4503), 
            .I3(n39679), .O(n39980));
    defparam i29951_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i29790_4_lut (.I0(n31_adj_4491), .I1(n29_adj_4490), .I2(n27_adj_4499), 
            .I3(n39980), .O(n39819));
    defparam i29790_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 add_5160_11_lut (.I0(GND_net), .I1(n9909[8]), .I2(n761), .I3(n32208), 
            .O(n9894[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5160_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30011_4_lut (.I0(n37_adj_4489), .I1(n35_adj_4494), .I2(n33_adj_4495), 
            .I3(n39819), .O(n40040));
    defparam i30011_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 duty_23__I_831_i16_3_lut (.I0(duty_23__N_3613[9]), .I1(duty_23__N_3613[21]), 
            .I2(n43_adj_4488), .I3(GND_net), .O(n16_adj_4507));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29927_3_lut (.I0(n6_adj_4508), .I1(duty_23__N_3613[10]), .I2(n21_adj_4503), 
            .I3(GND_net), .O(n39956));   // verilog/motorControl.v(36[10:25])
    defparam i29927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29928_3_lut (.I0(n39956), .I1(duty_23__N_3613[11]), .I2(n23_adj_4492), 
            .I3(GND_net), .O(n39957));   // verilog/motorControl.v(36[10:25])
    defparam i29928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_831_i8_3_lut (.I0(duty_23__N_3613[4]), .I1(duty_23__N_3613[8]), 
            .I2(n17_adj_4501), .I3(GND_net), .O(n8_adj_4509));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5160_11 (.CI(n32208), .I0(n9909[8]), .I1(n761), .CO(n32209));
    SB_LUT4 duty_23__I_831_i24_3_lut (.I0(n16_adj_4507), .I1(duty_23__N_3613[22]), 
            .I2(n45_adj_4487), .I3(GND_net), .O(n24_adj_4510));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29355_4_lut (.I0(n43_adj_4488), .I1(n25_adj_4493), .I2(n23_adj_4492), 
            .I3(n39407), .O(n39383));
    defparam i29355_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29826_4_lut (.I0(n24_adj_4510), .I1(n8_adj_4509), .I2(n45_adj_4487), 
            .I3(n39381), .O(n39855));   // verilog/motorControl.v(36[10:25])
    defparam i29826_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29883_3_lut (.I0(n39957), .I1(duty_23__N_3613[12]), .I2(n25_adj_4493), 
            .I3(GND_net), .O(n39912));   // verilog/motorControl.v(36[10:25])
    defparam i29883_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_831_i4_4_lut (.I0(duty_23__N_3613[0]), .I1(duty_23__N_3613[1]), 
            .I2(PWMLimit[1]), .I3(PWMLimit[0]), .O(n4_adj_4511));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i29925_3_lut (.I0(n4_adj_4511), .I1(duty_23__N_3613[13]), .I2(n27_adj_4499), 
            .I3(GND_net), .O(n39954));   // verilog/motorControl.v(36[10:25])
    defparam i29925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29926_3_lut (.I0(n39954), .I1(duty_23__N_3613[14]), .I2(n29_adj_4490), 
            .I3(GND_net), .O(n39955));   // verilog/motorControl.v(36[10:25])
    defparam i29926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29366_4_lut (.I0(n33_adj_4495), .I1(n31_adj_4491), .I2(n29_adj_4490), 
            .I3(n39399), .O(n39394));
    defparam i29366_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i30021_4_lut (.I0(n30_adj_4506), .I1(n10_adj_4505), .I2(n35_adj_4494), 
            .I3(n39392), .O(n40050));   // verilog/motorControl.v(36[10:25])
    defparam i30021_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i29885_3_lut (.I0(n39955), .I1(duty_23__N_3613[15]), .I2(n31_adj_4491), 
            .I3(GND_net), .O(n39914));   // verilog/motorControl.v(36[10:25])
    defparam i29885_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30072_4_lut (.I0(n39914), .I1(n40050), .I2(n35_adj_4494), 
            .I3(n39394), .O(n40101));   // verilog/motorControl.v(36[10:25])
    defparam i30072_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30073_3_lut (.I0(n40101), .I1(duty_23__N_3613[18]), .I2(n37_adj_4489), 
            .I3(GND_net), .O(n40102));   // verilog/motorControl.v(36[10:25])
    defparam i30073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30052_3_lut (.I0(n40102), .I1(duty_23__N_3613[19]), .I2(n39_adj_4485), 
            .I3(GND_net), .O(n40081));   // verilog/motorControl.v(36[10:25])
    defparam i30052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29357_4_lut (.I0(n43_adj_4488), .I1(n41_adj_4486), .I2(n39_adj_4485), 
            .I3(n40040), .O(n39385));
    defparam i29357_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i29981_4_lut (.I0(n39912), .I1(n39855), .I2(n45_adj_4487), 
            .I3(n39383), .O(n40010));   // verilog/motorControl.v(36[10:25])
    defparam i29981_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i30042_3_lut (.I0(n40081), .I1(duty_23__N_3613[20]), .I2(n41_adj_4486), 
            .I3(GND_net), .O(n40_adj_4512));   // verilog/motorControl.v(36[10:25])
    defparam i30042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29983_4_lut (.I0(n40_adj_4512), .I1(n40010), .I2(n45_adj_4487), 
            .I3(n39385), .O(n40012));   // verilog/motorControl.v(36[10:25])
    defparam i29983_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i29984_3_lut (.I0(n40012), .I1(PWMLimit[23]), .I2(duty_23__N_3613[23]), 
            .I3(GND_net), .O(duty_23__N_3612));   // verilog/motorControl.v(36[10:25])
    defparam i29984_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5160_10_lut (.I0(GND_net), .I1(n9909[7]), .I2(n688), .I3(n32207), 
            .O(n9894[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5160_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5160_10 (.CI(n32207), .I0(n9909[7]), .I1(n688), .CO(n32208));
    SB_CARRY add_5338_7 (.CI(n30766), .I0(n13223[4]), .I1(n472_adj_4330), 
            .CO(n30767));
    SB_LUT4 add_5160_9_lut (.I0(GND_net), .I1(n9909[6]), .I2(n615), .I3(n32206), 
            .O(n9894[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5160_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5338_6_lut (.I0(GND_net), .I1(n13223[3]), .I2(n399), .I3(n30765), 
            .O(n13080[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5338_6 (.CI(n30765), .I0(n13223[3]), .I1(n399), .CO(n30766));
    SB_CARRY add_5160_9 (.CI(n32206), .I0(n9909[6]), .I1(n615), .CO(n32207));
    SB_LUT4 add_5160_8_lut (.I0(GND_net), .I1(n9909[5]), .I2(n542), .I3(n32205), 
            .O(n9894[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5160_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5160_8 (.CI(n32205), .I0(n9909[5]), .I1(n542), .CO(n32206));
    SB_LUT4 add_5160_7_lut (.I0(GND_net), .I1(n9909[4]), .I2(n469), .I3(n32204), 
            .O(n9894[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5160_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5160_7 (.CI(n32204), .I0(n9909[4]), .I1(n469), .CO(n32205));
    SB_LUT4 mux_17_i1_3_lut (.I0(duty_23__N_3613[0]), .I1(n257[0]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i1_3_lut (.I0(duty_23__N_3588[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_18 (.CI(n30938), .I0(GND_net), .I1(n1_adj_4704[16]), 
            .CO(n30939));
    SB_LUT4 add_5160_6_lut (.I0(GND_net), .I1(n9909[3]), .I2(n396), .I3(n32203), 
            .O(n9894[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5160_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[15]), 
            .I3(n30937), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5383_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n31000));
    SB_LUT4 add_5313_15_lut (.I0(GND_net), .I1(n12912[12]), .I2(n1050_adj_4295), 
            .I3(n30999), .O(n12717[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5313_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5160_6 (.CI(n32203), .I0(n9909[3]), .I1(n396), .CO(n32204));
    SB_LUT4 add_5160_5_lut (.I0(GND_net), .I1(n9909[2]), .I2(n323), .I3(n32202), 
            .O(n9894[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5160_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5160_5 (.CI(n32202), .I0(n9909[2]), .I1(n323), .CO(n32203));
    SB_CARRY add_12_14 (.CI(n30728), .I0(n106[12]), .I1(n155[12]), .CO(n30729));
    SB_LUT4 add_5338_5_lut (.I0(GND_net), .I1(n13223[2]), .I2(n326), .I3(n30764), 
            .O(n13080[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5160_4_lut (.I0(GND_net), .I1(n9909[1]), .I2(n250), .I3(n32201), 
            .O(n9894[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5160_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5160_4 (.CI(n32201), .I0(n9909[1]), .I1(n250), .CO(n32202));
    SB_LUT4 add_5160_3_lut (.I0(GND_net), .I1(n9909[0]), .I2(n177), .I3(n32200), 
            .O(n9894[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5160_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5160_3 (.CI(n32200), .I0(n9909[0]), .I1(n177), .CO(n32201));
    SB_LUT4 add_723_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n3141[19]), .I3(n30812), .O(\PID_CONTROLLER.integral_23__N_3513 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5160_2_lut (.I0(GND_net), .I1(n35), .I2(n104), .I3(GND_net), 
            .O(n9894[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5160_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5160_2 (.CI(GND_net), .I0(n35), .I1(n104), .CO(n32200));
    SB_CARRY unary_minus_16_add_3_17 (.CI(n30937), .I0(GND_net), .I1(n1_adj_4704[15]), 
            .CO(n30938));
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[14]), 
            .I3(n30936), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5159_15_lut (.I0(GND_net), .I1(n9894[12]), .I2(n1050), 
            .I3(n32199), .O(n9878[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5313_14_lut (.I0(GND_net), .I1(n12912[11]), .I2(n977_adj_4293), 
            .I3(n30998), .O(n12717[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5313_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5159_14_lut (.I0(GND_net), .I1(n9894[11]), .I2(n977), 
            .I3(n32198), .O(n9878[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_16 (.CI(n30936), .I0(GND_net), .I1(n1_adj_4704[14]), 
            .CO(n30937));
    SB_CARRY add_5313_14 (.CI(n30998), .I0(n12912[11]), .I1(n977_adj_4293), 
            .CO(n30999));
    SB_CARRY add_5159_14 (.CI(n32198), .I0(n9894[11]), .I1(n977), .CO(n32199));
    SB_LUT4 add_5159_13_lut (.I0(GND_net), .I1(n9894[10]), .I2(n904_adj_4292), 
            .I3(n32197), .O(n9878[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_13 (.CI(n32197), .I0(n9894[10]), .I1(n904_adj_4292), 
            .CO(n32198));
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[13]), 
            .I3(n30935), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5159_12_lut (.I0(GND_net), .I1(n9894[9]), .I2(n831_adj_4290), 
            .I3(n32196), .O(n9878[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_723_21 (.CI(n30812), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n3141[19]), .CO(n30813));
    SB_CARRY add_5159_12 (.CI(n32196), .I0(n9894[9]), .I1(n831_adj_4290), 
            .CO(n32197));
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5159_11_lut (.I0(GND_net), .I1(n9894[8]), .I2(n758_adj_4289), 
            .I3(n32195), .O(n9878[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_723_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n3141[18]), .I3(n30811), .O(\PID_CONTROLLER.integral_23__N_3513 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_723_20 (.CI(n30811), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n3141[18]), .CO(n30812));
    SB_CARRY add_5338_5 (.CI(n30764), .I0(n13223[2]), .I1(n326), .CO(n30765));
    SB_CARRY add_5159_11 (.CI(n32195), .I0(n9894[8]), .I1(n758_adj_4289), 
            .CO(n32196));
    SB_LUT4 add_5159_10_lut (.I0(GND_net), .I1(n9894[7]), .I2(n685_adj_4288), 
            .I3(n32194), .O(n9878[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n30935), .I0(GND_net), .I1(n1_adj_4704[13]), 
            .CO(n30936));
    SB_CARRY add_5159_10 (.CI(n32194), .I0(n9894[7]), .I1(n685_adj_4288), 
            .CO(n32195));
    SB_LUT4 add_5159_9_lut (.I0(GND_net), .I1(n9894[6]), .I2(n612), .I3(n32193), 
            .O(n9878[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_13_lut (.I0(GND_net), .I1(n106[11]), .I2(n155[11]), 
            .I3(n30727), .O(duty_23__N_3613[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5338_4_lut (.I0(GND_net), .I1(n13223[1]), .I2(n253), .I3(n30763), 
            .O(n13080[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_13 (.CI(n30727), .I0(n106[11]), .I1(n155[11]), .CO(n30728));
    SB_CARRY add_5159_9 (.CI(n32193), .I0(n9894[6]), .I1(n612), .CO(n32194));
    SB_LUT4 add_5159_8_lut (.I0(GND_net), .I1(n9894[5]), .I2(n539), .I3(n32192), 
            .O(n9878[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_8 (.CI(n32192), .I0(n9894[5]), .I1(n539), .CO(n32193));
    SB_LUT4 add_5159_7_lut (.I0(GND_net), .I1(n9894[4]), .I2(n466), .I3(n32191), 
            .O(n9878[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_7 (.CI(n32191), .I0(n9894[4]), .I1(n466), .CO(n32192));
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[12]), 
            .I3(n30934), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n30934), .I0(GND_net), .I1(n1_adj_4704[12]), 
            .CO(n30935));
    SB_LUT4 add_5313_13_lut (.I0(GND_net), .I1(n12912[10]), .I2(n904), 
            .I3(n30997), .O(n12717[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5313_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5159_6_lut (.I0(GND_net), .I1(n9894[3]), .I2(n393), .I3(n32190), 
            .O(n9878[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_6 (.CI(n32190), .I0(n9894[3]), .I1(n393), .CO(n32191));
    SB_LUT4 add_5159_5_lut (.I0(GND_net), .I1(n9894[2]), .I2(n320), .I3(n32189), 
            .O(n9878[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_723_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n3141[17]), .I3(n30810), .O(\PID_CONTROLLER.integral_23__N_3513 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_5 (.CI(n32189), .I0(n9894[2]), .I1(n320), .CO(n32190));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[11]), 
            .I3(n30933), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5159_4_lut (.I0(GND_net), .I1(n9894[1]), .I2(n247), .I3(n32188), 
            .O(n9878[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5159_4 (.CI(n32188), .I0(n9894[1]), .I1(n247), .CO(n32189));
    SB_LUT4 add_5159_3_lut (.I0(GND_net), .I1(n9894[0]), .I2(n174), .I3(n32187), 
            .O(n9878[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_723_19 (.CI(n30810), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n3141[17]), .CO(n30811));
    SB_CARRY add_5159_3 (.CI(n32187), .I0(n9894[0]), .I1(n174), .CO(n32188));
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(n28[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4360));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4359));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5159_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n9878[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5159_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5338_4 (.CI(n30763), .I0(n13223[1]), .I1(n253), .CO(n30764));
    SB_CARRY add_5159_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n32187));
    SB_LUT4 add_12_12_lut (.I0(GND_net), .I1(n106[10]), .I2(n155[10]), 
            .I3(n30726), .O(duty_23__N_3613[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5158_16_lut (.I0(GND_net), .I1(n9878[13]), .I2(n1120), 
            .I3(n32186), .O(n9861[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5158_15_lut (.I0(GND_net), .I1(n9878[12]), .I2(n1047), 
            .I3(n32185), .O(n9861[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5158_15 (.CI(n32185), .I0(n9878[12]), .I1(n1047), .CO(n32186));
    SB_LUT4 add_5158_14_lut (.I0(GND_net), .I1(n9878[11]), .I2(n974), 
            .I3(n32184), .O(n9861[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5158_14 (.CI(n32184), .I0(n9878[11]), .I1(n974), .CO(n32185));
    SB_LUT4 add_723_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n3141[16]), .I3(n30809), .O(\PID_CONTROLLER.integral_23__N_3513 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5158_13_lut (.I0(GND_net), .I1(n9878[10]), .I2(n901), 
            .I3(n32183), .O(n9861[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5158_13 (.CI(n32183), .I0(n9878[10]), .I1(n901), .CO(n32184));
    SB_LUT4 add_5338_3_lut (.I0(GND_net), .I1(n13223[0]), .I2(n180), .I3(n30762), 
            .O(n13080[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5158_12_lut (.I0(GND_net), .I1(n9878[9]), .I2(n828), .I3(n32182), 
            .O(n9861[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5158_12 (.CI(n32182), .I0(n9878[9]), .I1(n828), .CO(n32183));
    SB_CARRY add_723_18 (.CI(n30809), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n3141[16]), .CO(n30810));
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244_adj_4335));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317_adj_4332));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5338_3 (.CI(n30762), .I0(n13223[0]), .I1(n180), .CO(n30763));
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390_adj_4315));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5158_11_lut (.I0(GND_net), .I1(n9878[8]), .I2(n755), .I3(n32181), 
            .O(n9861[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5158_11 (.CI(n32181), .I0(n9878[8]), .I1(n755), .CO(n32182));
    SB_CARRY unary_minus_16_add_3_13 (.CI(n30933), .I0(GND_net), .I1(n1_adj_4704[11]), 
            .CO(n30934));
    SB_LUT4 add_5158_10_lut (.I0(GND_net), .I1(n9878[7]), .I2(n682), .I3(n32180), 
            .O(n9861[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_12 (.CI(n30726), .I0(n106[10]), .I1(n155[10]), .CO(n30727));
    SB_LUT4 add_723_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n3141[15]), .I3(n30808), .O(\PID_CONTROLLER.integral_23__N_3513 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5338_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n13080[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5338_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5313_13 (.CI(n30997), .I0(n12912[10]), .I1(n904), .CO(n30998));
    SB_CARRY add_5158_10 (.CI(n32180), .I0(n9878[7]), .I1(n682), .CO(n32181));
    SB_LUT4 add_5158_9_lut (.I0(GND_net), .I1(n9878[6]), .I2(n609), .I3(n32179), 
            .O(n9861[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5158_9 (.CI(n32179), .I0(n9878[6]), .I1(n609), .CO(n32180));
    SB_LUT4 add_5158_8_lut (.I0(GND_net), .I1(n9878[5]), .I2(n536), .I3(n32178), 
            .O(n9861[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5158_8 (.CI(n32178), .I0(n9878[5]), .I1(n536), .CO(n32179));
    SB_LUT4 add_5158_7_lut (.I0(GND_net), .I1(n9878[4]), .I2(n463_adj_4283), 
            .I3(n32177), .O(n9861[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(n28[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4298));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[10]), 
            .I3(n30932), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_24_lut (.I0(n28[23]), .I1(n9589[21]), .I2(GND_net), 
            .I3(n31521), .O(n7896[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_723_17 (.CI(n30808), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n3141[15]), .CO(n30809));
    SB_CARRY add_5158_7 (.CI(n32177), .I0(n9878[4]), .I1(n463_adj_4283), 
            .CO(n32178));
    SB_LUT4 mult_10_add_1225_23_lut (.I0(GND_net), .I1(n9589[20]), .I2(GND_net), 
            .I3(n31520), .O(n106[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5158_6_lut (.I0(GND_net), .I1(n9878[3]), .I2(n390), .I3(n32176), 
            .O(n9861[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_23 (.CI(n31520), .I0(n9589[20]), .I1(GND_net), 
            .CO(n31521));
    SB_CARRY add_5158_6 (.CI(n32176), .I0(n9878[3]), .I1(n390), .CO(n32177));
    SB_LUT4 add_5158_5_lut (.I0(GND_net), .I1(n9878[2]), .I2(n317), .I3(n32175), 
            .O(n9861[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5158_5 (.CI(n32175), .I0(n9878[2]), .I1(n317), .CO(n32176));
    SB_LUT4 add_5158_4_lut (.I0(GND_net), .I1(n9878[1]), .I2(n244), .I3(n32174), 
            .O(n9861[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n30932), .I0(GND_net), .I1(n1_adj_4704[10]), 
            .CO(n30933));
    SB_LUT4 mult_10_add_1225_22_lut (.I0(GND_net), .I1(n9589[19]), .I2(GND_net), 
            .I3(n31519), .O(n106[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_22 (.CI(n31519), .I0(n9589[19]), .I1(GND_net), 
            .CO(n31520));
    SB_LUT4 add_723_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n3141[14]), .I3(n30807), .O(\PID_CONTROLLER.integral_23__N_3513 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5158_4 (.CI(n32174), .I0(n9878[1]), .I1(n244), .CO(n32175));
    SB_CARRY add_723_16 (.CI(n30807), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n3141[14]), .CO(n30808));
    SB_LUT4 add_5158_3_lut (.I0(GND_net), .I1(n9878[0]), .I2(n171), .I3(n32173), 
            .O(n9861[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_21_lut (.I0(GND_net), .I1(n9589[18]), .I2(GND_net), 
            .I3(n31518), .O(n106[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5313_12_lut (.I0(GND_net), .I1(n12912[9]), .I2(n831), 
            .I3(n30996), .O(n12717[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5313_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_21 (.CI(n31518), .I0(n9589[18]), .I1(GND_net), 
            .CO(n31519));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[9]), 
            .I3(n30931), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_20_lut (.I0(GND_net), .I1(n9589[17]), .I2(GND_net), 
            .I3(n31517), .O(n106[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5338_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n30762));
    SB_CARRY add_5158_3 (.CI(n32173), .I0(n9878[0]), .I1(n171), .CO(n32174));
    SB_CARRY mult_10_add_1225_20 (.CI(n31517), .I0(n9589[17]), .I1(GND_net), 
            .CO(n31518));
    SB_LUT4 add_5158_2_lut (.I0(GND_net), .I1(n29), .I2(n98), .I3(GND_net), 
            .O(n9861[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5158_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_19_lut (.I0(GND_net), .I1(n9589[16]), .I2(GND_net), 
            .I3(n31516), .O(n106[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5158_2 (.CI(GND_net), .I0(n29), .I1(n98), .CO(n32173));
    SB_CARRY unary_minus_16_add_3_11 (.CI(n30931), .I0(GND_net), .I1(n1_adj_4704[9]), 
            .CO(n30932));
    SB_LUT4 add_5157_17_lut (.I0(GND_net), .I1(n9861[14]), .I2(GND_net), 
            .I3(n32172), .O(n9843[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5157_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[8]), 
            .I3(n30930), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5157_16_lut (.I0(GND_net), .I1(n9861[13]), .I2(n1117), 
            .I3(n32171), .O(n9843[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5157_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n30930), .I0(GND_net), .I1(n1_adj_4704[8]), 
            .CO(n30931));
    SB_CARRY add_5157_16 (.CI(n32171), .I0(n9861[13]), .I1(n1117), .CO(n32172));
    SB_CARRY add_5313_12 (.CI(n30996), .I0(n12912[9]), .I1(n831), .CO(n30997));
    SB_LUT4 add_5157_15_lut (.I0(GND_net), .I1(n9861[12]), .I2(n1044), 
            .I3(n32170), .O(n9843[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5157_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_19 (.CI(n31516), .I0(n9589[16]), .I1(GND_net), 
            .CO(n31517));
    SB_CARRY add_5157_15 (.CI(n32170), .I0(n9861[12]), .I1(n1044), .CO(n32171));
    SB_LUT4 add_5157_14_lut (.I0(GND_net), .I1(n9861[11]), .I2(n971), 
            .I3(n32169), .O(n9843[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5157_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5313_11_lut (.I0(GND_net), .I1(n12912[8]), .I2(n758), 
            .I3(n30995), .O(n12717[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5313_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5313_11 (.CI(n30995), .I0(n12912[8]), .I1(n758), .CO(n30996));
    SB_CARRY add_5157_14 (.CI(n32169), .I0(n9861[11]), .I1(n971), .CO(n32170));
    SB_LUT4 add_5313_10_lut (.I0(GND_net), .I1(n12912[7]), .I2(n685), 
            .I3(n30994), .O(n12717[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5313_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5157_13_lut (.I0(GND_net), .I1(n9861[10]), .I2(n898), 
            .I3(n32168), .O(n9843[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5157_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_18_lut (.I0(GND_net), .I1(n9589[15]), .I2(GND_net), 
            .I3(n31515), .O(n106[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_18 (.CI(n31515), .I0(n9589[15]), .I1(GND_net), 
            .CO(n31516));
    SB_LUT4 mult_10_add_1225_17_lut (.I0(GND_net), .I1(n9589[14]), .I2(GND_net), 
            .I3(n31514), .O(n106[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_17 (.CI(n31514), .I0(n9589[14]), .I1(GND_net), 
            .CO(n31515));
    SB_CARRY add_5313_10 (.CI(n30994), .I0(n12912[7]), .I1(n685), .CO(n30995));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[7]), 
            .I3(n30929), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_16_lut (.I0(GND_net), .I1(n9589[13]), .I2(n1096), 
            .I3(n31513), .O(n106[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_723_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n3141[13]), .I3(n30806), .O(\PID_CONTROLLER.integral_23__N_3513 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_16 (.CI(n31513), .I0(n9589[13]), .I1(n1096), 
            .CO(n31514));
    SB_CARRY unary_minus_16_add_3_9 (.CI(n30929), .I0(GND_net), .I1(n1_adj_4704[7]), 
            .CO(n30930));
    SB_LUT4 add_12_11_lut (.I0(GND_net), .I1(n106[9]), .I2(n155[9]), .I3(n30725), 
            .O(duty_23__N_3613[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[6]), 
            .I3(n30928), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5157_13 (.CI(n32168), .I0(n9861[10]), .I1(n898), .CO(n32169));
    SB_LUT4 mult_10_add_1225_15_lut (.I0(GND_net), .I1(n9589[12]), .I2(n1023), 
            .I3(n31512), .O(n106[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5157_12_lut (.I0(GND_net), .I1(n9861[9]), .I2(n825), .I3(n32167), 
            .O(n9843[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5157_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5157_12 (.CI(n32167), .I0(n9861[9]), .I1(n825), .CO(n32168));
    SB_LUT4 add_5157_11_lut (.I0(GND_net), .I1(n9861[8]), .I2(n752), .I3(n32166), 
            .O(n9843[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5157_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5157_11 (.CI(n32166), .I0(n9861[8]), .I1(n752), .CO(n32167));
    SB_LUT4 add_5157_10_lut (.I0(GND_net), .I1(n9861[7]), .I2(n679), .I3(n32165), 
            .O(n9843[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5157_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5157_10 (.CI(n32165), .I0(n9861[7]), .I1(n679), .CO(n32166));
    SB_LUT4 add_5157_9_lut (.I0(GND_net), .I1(n9861[6]), .I2(n606_adj_4514), 
            .I3(n32164), .O(n9843[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5157_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5157_9 (.CI(n32164), .I0(n9861[6]), .I1(n606_adj_4514), 
            .CO(n32165));
    SB_LUT4 add_5157_8_lut (.I0(GND_net), .I1(n9861[5]), .I2(n533_adj_4515), 
            .I3(n32163), .O(n9843[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5157_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_15 (.CI(n31512), .I0(n9589[12]), .I1(n1023), 
            .CO(n31513));
    SB_CARRY add_5157_8 (.CI(n32163), .I0(n9861[5]), .I1(n533_adj_4515), 
            .CO(n32164));
    SB_LUT4 add_5157_7_lut (.I0(GND_net), .I1(n9861[4]), .I2(n460), .I3(n32162), 
            .O(n9843[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5157_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5157_7 (.CI(n32162), .I0(n9861[4]), .I1(n460), .CO(n32163));
    SB_LUT4 add_5157_6_lut (.I0(GND_net), .I1(n9861[3]), .I2(n387), .I3(n32161), 
            .O(n9843[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5157_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5157_6 (.CI(n32161), .I0(n9861[3]), .I1(n387), .CO(n32162));
    SB_LUT4 add_5157_5_lut (.I0(GND_net), .I1(n9861[2]), .I2(n314), .I3(n32160), 
            .O(n9843[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5157_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5157_5 (.CI(n32160), .I0(n9861[2]), .I1(n314), .CO(n32161));
    SB_LUT4 add_5157_4_lut (.I0(GND_net), .I1(n9861[1]), .I2(n241), .I3(n32159), 
            .O(n9843[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5157_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5157_4 (.CI(n32159), .I0(n9861[1]), .I1(n241), .CO(n32160));
    SB_LUT4 add_5157_3_lut (.I0(GND_net), .I1(n9861[0]), .I2(n168), .I3(n32158), 
            .O(n9843[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5157_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5157_3 (.CI(n32158), .I0(n9861[0]), .I1(n168), .CO(n32159));
    SB_LUT4 add_5157_2_lut (.I0(GND_net), .I1(n26_adj_4516), .I2(n95), 
            .I3(GND_net), .O(n9843[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5157_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5157_2 (.CI(GND_net), .I0(n26_adj_4516), .I1(n95), .CO(n32158));
    SB_LUT4 add_5156_18_lut (.I0(GND_net), .I1(n9843[15]), .I2(GND_net), 
            .I3(n32157), .O(n9824[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5156_17_lut (.I0(GND_net), .I1(n9843[14]), .I2(GND_net), 
            .I3(n32156), .O(n9824[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_17 (.CI(n32156), .I0(n9843[14]), .I1(GND_net), .CO(n32157));
    SB_LUT4 add_5156_16_lut (.I0(GND_net), .I1(n9843[13]), .I2(n1114_adj_4517), 
            .I3(n32155), .O(n9824[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_16 (.CI(n32155), .I0(n9843[13]), .I1(n1114_adj_4517), 
            .CO(n32156));
    SB_LUT4 add_5156_15_lut (.I0(GND_net), .I1(n9843[12]), .I2(n1041_adj_4518), 
            .I3(n32154), .O(n9824[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_11 (.CI(n30725), .I0(n106[9]), .I1(n155[9]), .CO(n30726));
    SB_LUT4 add_5313_9_lut (.I0(GND_net), .I1(n12912[6]), .I2(n612_adj_4519), 
            .I3(n30993), .O(n12717[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5313_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_15 (.CI(n32154), .I0(n9843[12]), .I1(n1041_adj_4518), 
            .CO(n32155));
    SB_LUT4 add_5156_14_lut (.I0(GND_net), .I1(n9843[11]), .I2(n968_adj_4520), 
            .I3(n32153), .O(n9824[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_14 (.CI(n32153), .I0(n9843[11]), .I1(n968_adj_4520), 
            .CO(n32154));
    SB_LUT4 add_5156_13_lut (.I0(GND_net), .I1(n9843[10]), .I2(n895_adj_4521), 
            .I3(n32152), .O(n9824[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_13 (.CI(n32152), .I0(n9843[10]), .I1(n895_adj_4521), 
            .CO(n32153));
    SB_CARRY unary_minus_16_add_3_8 (.CI(n30928), .I0(GND_net), .I1(n1_adj_4704[6]), 
            .CO(n30929));
    SB_LUT4 add_5156_12_lut (.I0(GND_net), .I1(n9843[9]), .I2(n822_adj_4522), 
            .I3(n32151), .O(n9824[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[5]), 
            .I3(n30927), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_12 (.CI(n32151), .I0(n9843[9]), .I1(n822_adj_4522), 
            .CO(n32152));
    SB_LUT4 mult_10_add_1225_14_lut (.I0(GND_net), .I1(n9589[11]), .I2(n950), 
            .I3(n31511), .O(n106[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5156_11_lut (.I0(GND_net), .I1(n9843[8]), .I2(n749_adj_4524), 
            .I3(n32150), .O(n9824[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_11 (.CI(n32150), .I0(n9843[8]), .I1(n749_adj_4524), 
            .CO(n32151));
    SB_LUT4 add_5156_10_lut (.I0(GND_net), .I1(n9843[7]), .I2(n676_adj_4525), 
            .I3(n32149), .O(n9824[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_10 (.CI(n32149), .I0(n9843[7]), .I1(n676_adj_4525), 
            .CO(n32150));
    SB_LUT4 add_5156_9_lut (.I0(GND_net), .I1(n9843[6]), .I2(n603_adj_4526), 
            .I3(n32148), .O(n9824[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_9 (.CI(n32148), .I0(n9843[6]), .I1(n603_adj_4526), 
            .CO(n32149));
    SB_LUT4 add_5156_8_lut (.I0(GND_net), .I1(n9843[5]), .I2(n530_adj_4527), 
            .I3(n32147), .O(n9824[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_8 (.CI(n32147), .I0(n9843[5]), .I1(n530_adj_4527), 
            .CO(n32148));
    SB_LUT4 add_5156_7_lut (.I0(GND_net), .I1(n9843[4]), .I2(n457_adj_4528), 
            .I3(n32146), .O(n9824[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_7 (.CI(n32146), .I0(n9843[4]), .I1(n457_adj_4528), 
            .CO(n32147));
    SB_LUT4 add_5156_6_lut (.I0(GND_net), .I1(n9843[3]), .I2(n384_adj_4529), 
            .I3(n32145), .O(n9824[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_6 (.CI(n32145), .I0(n9843[3]), .I1(n384_adj_4529), 
            .CO(n32146));
    SB_LUT4 add_5156_5_lut (.I0(GND_net), .I1(n9843[2]), .I2(n311_adj_4530), 
            .I3(n32144), .O(n9824[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_5 (.CI(n32144), .I0(n9843[2]), .I1(n311_adj_4530), 
            .CO(n32145));
    SB_LUT4 add_5156_4_lut (.I0(GND_net), .I1(n9843[1]), .I2(n238_adj_4531), 
            .I3(n32143), .O(n9824[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_4 (.CI(n32143), .I0(n9843[1]), .I1(n238_adj_4531), 
            .CO(n32144));
    SB_LUT4 add_5156_3_lut (.I0(GND_net), .I1(n9843[0]), .I2(n165_adj_4532), 
            .I3(n32142), .O(n9824[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5313_9 (.CI(n30993), .I0(n12912[6]), .I1(n612_adj_4519), 
            .CO(n30994));
    SB_CARRY add_5156_3 (.CI(n32142), .I0(n9843[0]), .I1(n165_adj_4532), 
            .CO(n32143));
    SB_LUT4 add_5156_2_lut (.I0(GND_net), .I1(n23_adj_4533), .I2(n92_adj_4534), 
            .I3(GND_net), .O(n9824[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5156_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5156_2 (.CI(GND_net), .I0(n23_adj_4533), .I1(n92_adj_4534), 
            .CO(n32142));
    SB_LUT4 add_5155_19_lut (.I0(GND_net), .I1(n9824[16]), .I2(GND_net), 
            .I3(n32141), .O(n9804[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5155_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5155_18_lut (.I0(GND_net), .I1(n9824[15]), .I2(GND_net), 
            .I3(n32140), .O(n9804[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5155_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5155_18 (.CI(n32140), .I0(n9824[15]), .I1(GND_net), .CO(n32141));
    SB_LUT4 add_5155_17_lut (.I0(GND_net), .I1(n9824[14]), .I2(GND_net), 
            .I3(n32139), .O(n9804[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5155_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5155_17 (.CI(n32139), .I0(n9824[14]), .I1(GND_net), .CO(n32140));
    SB_LUT4 add_5155_16_lut (.I0(GND_net), .I1(n9824[13]), .I2(n1111_adj_4535), 
            .I3(n32138), .O(n9804[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5155_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5155_16 (.CI(n32138), .I0(n9824[13]), .I1(n1111_adj_4535), 
            .CO(n32139));
    SB_LUT4 add_5155_15_lut (.I0(GND_net), .I1(n9824[12]), .I2(n1038_adj_4536), 
            .I3(n32137), .O(n9804[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5155_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5155_15 (.CI(n32137), .I0(n9824[12]), .I1(n1038_adj_4536), 
            .CO(n32138));
    SB_LUT4 add_5155_14_lut (.I0(GND_net), .I1(n9824[11]), .I2(n965_adj_4537), 
            .I3(n32136), .O(n9804[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5155_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5155_14 (.CI(n32136), .I0(n9824[11]), .I1(n965_adj_4537), 
            .CO(n32137));
    SB_LUT4 add_5313_8_lut (.I0(GND_net), .I1(n12912[5]), .I2(n539_adj_4538), 
            .I3(n30992), .O(n12717[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5313_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5155_13_lut (.I0(GND_net), .I1(n9824[10]), .I2(n892_adj_4539), 
            .I3(n32135), .O(n9804[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5155_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5155_13 (.CI(n32135), .I0(n9824[10]), .I1(n892_adj_4539), 
            .CO(n32136));
    SB_LUT4 add_5155_12_lut (.I0(GND_net), .I1(n9824[9]), .I2(n819_adj_4540), 
            .I3(n32134), .O(n9804[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5155_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5155_12 (.CI(n32134), .I0(n9824[9]), .I1(n819_adj_4540), 
            .CO(n32135));
    SB_LUT4 add_5155_11_lut (.I0(GND_net), .I1(n9824[8]), .I2(n746_adj_4541), 
            .I3(n32133), .O(n9804[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5155_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5155_11 (.CI(n32133), .I0(n9824[8]), .I1(n746_adj_4541), 
            .CO(n32134));
    SB_LUT4 add_5155_10_lut (.I0(GND_net), .I1(n9824[7]), .I2(n673_adj_4542), 
            .I3(n32132), .O(n9804[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5155_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5155_10 (.CI(n32132), .I0(n9824[7]), .I1(n673_adj_4542), 
            .CO(n32133));
    SB_LUT4 add_5155_9_lut (.I0(GND_net), .I1(n9824[6]), .I2(n600_adj_4543), 
            .I3(n32131), .O(n9804[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5155_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5155_9 (.CI(n32131), .I0(n9824[6]), .I1(n600_adj_4543), 
            .CO(n32132));
    SB_LUT4 add_5155_8_lut (.I0(GND_net), .I1(n9824[5]), .I2(n527_adj_4544), 
            .I3(n32130), .O(n9804[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5155_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5155_8 (.CI(n32130), .I0(n9824[5]), .I1(n527_adj_4544), 
            .CO(n32131));
    SB_LUT4 add_5155_7_lut (.I0(GND_net), .I1(n9824[4]), .I2(n454_adj_4545), 
            .I3(n32129), .O(n9804[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5155_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_723_15 (.CI(n30806), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n3141[13]), .CO(n30807));
    SB_CARRY add_5155_7 (.CI(n32129), .I0(n9824[4]), .I1(n454_adj_4545), 
            .CO(n32130));
    SB_LUT4 add_723_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n3141[12]), .I3(n30805), .O(\PID_CONTROLLER.integral_23__N_3513 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5155_6_lut (.I0(GND_net), .I1(n9824[3]), .I2(n381_adj_4546), 
            .I3(n32128), .O(n9804[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5155_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_10_lut (.I0(GND_net), .I1(n106[8]), .I2(n155[8]), .I3(n30724), 
            .O(duty_23__N_3613[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5155_6 (.CI(n32128), .I0(n9824[3]), .I1(n381_adj_4546), 
            .CO(n32129));
    SB_LUT4 add_5155_5_lut (.I0(GND_net), .I1(n9824[2]), .I2(n308_adj_4548), 
            .I3(n32127), .O(n9804[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5155_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5155_5 (.CI(n32127), .I0(n9824[2]), .I1(n308_adj_4548), 
            .CO(n32128));
    SB_LUT4 add_5155_4_lut (.I0(GND_net), .I1(n9824[1]), .I2(n235_adj_4549), 
            .I3(n32126), .O(n9804[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5155_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5155_4 (.CI(n32126), .I0(n9824[1]), .I1(n235_adj_4549), 
            .CO(n32127));
    SB_LUT4 add_5155_3_lut (.I0(GND_net), .I1(n9824[0]), .I2(n162_adj_4550), 
            .I3(n32125), .O(n9804[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5155_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5155_3 (.CI(n32125), .I0(n9824[0]), .I1(n162_adj_4550), 
            .CO(n32126));
    SB_LUT4 add_5155_2_lut (.I0(GND_net), .I1(n20_adj_4551), .I2(n89_adj_4552), 
            .I3(GND_net), .O(n9804[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5155_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5155_2 (.CI(GND_net), .I0(n20_adj_4551), .I1(n89_adj_4552), 
            .CO(n32125));
    SB_LUT4 add_5154_20_lut (.I0(GND_net), .I1(n9804[17]), .I2(GND_net), 
            .I3(n32124), .O(n9783[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5154_19_lut (.I0(GND_net), .I1(n9804[16]), .I2(GND_net), 
            .I3(n32123), .O(n9783[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5154_19 (.CI(n32123), .I0(n9804[16]), .I1(GND_net), .CO(n32124));
    SB_CARRY unary_minus_16_add_3_7 (.CI(n30927), .I0(GND_net), .I1(n1_adj_4704[5]), 
            .CO(n30928));
    SB_LUT4 add_5154_18_lut (.I0(GND_net), .I1(n9804[15]), .I2(GND_net), 
            .I3(n32122), .O(n9783[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5154_18 (.CI(n32122), .I0(n9804[15]), .I1(GND_net), .CO(n32123));
    SB_LUT4 add_5154_17_lut (.I0(GND_net), .I1(n9804[14]), .I2(GND_net), 
            .I3(n32121), .O(n9783[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5154_17 (.CI(n32121), .I0(n9804[14]), .I1(GND_net), .CO(n32122));
    SB_LUT4 add_5154_16_lut (.I0(GND_net), .I1(n9804[13]), .I2(n1108_adj_4553), 
            .I3(n32120), .O(n9783[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5154_16 (.CI(n32120), .I0(n9804[13]), .I1(n1108_adj_4553), 
            .CO(n32121));
    SB_CARRY add_12_10 (.CI(n30724), .I0(n106[8]), .I1(n155[8]), .CO(n30725));
    SB_LUT4 add_5154_15_lut (.I0(GND_net), .I1(n9804[12]), .I2(n1035_adj_4554), 
            .I3(n32119), .O(n9783[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5154_15 (.CI(n32119), .I0(n9804[12]), .I1(n1035_adj_4554), 
            .CO(n32120));
    SB_LUT4 add_5154_14_lut (.I0(GND_net), .I1(n9804[11]), .I2(n962_adj_4555), 
            .I3(n32118), .O(n9783[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5154_14 (.CI(n32118), .I0(n9804[11]), .I1(n962_adj_4555), 
            .CO(n32119));
    SB_CARRY add_5313_8 (.CI(n30992), .I0(n12912[5]), .I1(n539_adj_4538), 
            .CO(n30993));
    SB_LUT4 add_5154_13_lut (.I0(GND_net), .I1(n9804[10]), .I2(n889_adj_4556), 
            .I3(n32117), .O(n9783[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5154_13 (.CI(n32117), .I0(n9804[10]), .I1(n889_adj_4556), 
            .CO(n32118));
    SB_LUT4 add_12_9_lut (.I0(GND_net), .I1(n106[7]), .I2(n155[7]), .I3(n30723), 
            .O(duty_23__N_3613[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5154_12_lut (.I0(GND_net), .I1(n9804[9]), .I2(n816_adj_4557), 
            .I3(n32116), .O(n9783[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5154_12 (.CI(n32116), .I0(n9804[9]), .I1(n816_adj_4557), 
            .CO(n32117));
    SB_LUT4 add_5154_11_lut (.I0(GND_net), .I1(n9804[8]), .I2(n743_adj_4558), 
            .I3(n32115), .O(n9783[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5154_11 (.CI(n32115), .I0(n9804[8]), .I1(n743_adj_4558), 
            .CO(n32116));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[4]), 
            .I3(n30926), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5154_10_lut (.I0(GND_net), .I1(n9804[7]), .I2(n670_adj_4560), 
            .I3(n32114), .O(n9783[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5154_10 (.CI(n32114), .I0(n9804[7]), .I1(n670_adj_4560), 
            .CO(n32115));
    SB_LUT4 add_5154_9_lut (.I0(GND_net), .I1(n9804[6]), .I2(n597_adj_4561), 
            .I3(n32113), .O(n9783[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n30926), .I0(GND_net), .I1(n1_adj_4704[4]), 
            .CO(n30927));
    SB_CARRY add_5154_9 (.CI(n32113), .I0(n9804[6]), .I1(n597_adj_4561), 
            .CO(n32114));
    SB_CARRY add_723_14 (.CI(n30805), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n3141[12]), .CO(n30806));
    SB_LUT4 add_5154_8_lut (.I0(GND_net), .I1(n9804[5]), .I2(n524_adj_4562), 
            .I3(n32112), .O(n9783[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5154_8 (.CI(n32112), .I0(n9804[5]), .I1(n524_adj_4562), 
            .CO(n32113));
    SB_LUT4 add_723_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n3141[11]), .I3(n30804), .O(\PID_CONTROLLER.integral_23__N_3513 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5154_7_lut (.I0(GND_net), .I1(n9804[4]), .I2(n451_adj_4563), 
            .I3(n32111), .O(n9783[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5154_7 (.CI(n32111), .I0(n9804[4]), .I1(n451_adj_4563), 
            .CO(n32112));
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[3]), 
            .I3(n30925), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5154_6_lut (.I0(GND_net), .I1(n9804[3]), .I2(n378_adj_4565), 
            .I3(n32110), .O(n9783[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5154_6 (.CI(n32110), .I0(n9804[3]), .I1(n378_adj_4565), 
            .CO(n32111));
    SB_CARRY add_723_13 (.CI(n30804), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n3141[11]), .CO(n30805));
    SB_CARRY add_12_9 (.CI(n30723), .I0(n106[7]), .I1(n155[7]), .CO(n30724));
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469_adj_4566));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_723_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n3141[10]), .I3(n30803), .O(\PID_CONTROLLER.integral_23__N_3513 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n30925), .I0(GND_net), .I1(n1_adj_4704[3]), 
            .CO(n30926));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[2]), 
            .I3(n30924), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5313_7_lut (.I0(GND_net), .I1(n12912[4]), .I2(n466_adj_4568), 
            .I3(n30991), .O(n12717[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5313_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_723_12 (.CI(n30803), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n3141[10]), .CO(n30804));
    SB_LUT4 add_12_8_lut (.I0(GND_net), .I1(n106[6]), .I2(n155[6]), .I3(n30722), 
            .O(duty_23__N_3613[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5313_7 (.CI(n30991), .I0(n12912[4]), .I1(n466_adj_4568), 
            .CO(n30992));
    SB_CARRY unary_minus_16_add_3_4 (.CI(n30924), .I0(GND_net), .I1(n1_adj_4704[2]), 
            .CO(n30925));
    SB_LUT4 add_5313_6_lut (.I0(GND_net), .I1(n12912[3]), .I2(n393_adj_4569), 
            .I3(n30990), .O(n12717[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5313_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_8 (.CI(n30722), .I0(n106[6]), .I1(n155[6]), .CO(n30723));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[1]), 
            .I3(n30923), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n30923), .I0(GND_net), .I1(n1_adj_4704[1]), 
            .CO(n30924));
    SB_LUT4 mult_10_add_1225_10_lut (.I0(GND_net), .I1(n9589[7]), .I2(n658), 
            .I3(n31507), .O(n106[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_723_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n3141[9]), .I3(n30802), .O(\PID_CONTROLLER.integral_23__N_3513 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_7_lut (.I0(GND_net), .I1(n106[5]), .I2(n155[5]), .I3(n30721), 
            .O(duty_23__N_3613[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5313_6 (.CI(n30990), .I0(n12912[3]), .I1(n393_adj_4569), 
            .CO(n30991));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4704[0]), 
            .I3(VCC_net), .O(n257[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4704[0]), 
            .CO(n30923));
    SB_LUT4 add_5154_5_lut (.I0(GND_net), .I1(n9804[2]), .I2(n305_adj_4573), 
            .I3(n32109), .O(n9783[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5154_5 (.CI(n32109), .I0(n9804[2]), .I1(n305_adj_4573), 
            .CO(n32110));
    SB_LUT4 add_5154_4_lut (.I0(GND_net), .I1(n9804[1]), .I2(n232_adj_4574), 
            .I3(n32108), .O(n9783[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5154_4 (.CI(n32108), .I0(n9804[1]), .I1(n232_adj_4574), 
            .CO(n32109));
    SB_LUT4 add_5154_3_lut (.I0(GND_net), .I1(n9804[0]), .I2(n159_adj_4575), 
            .I3(n32107), .O(n9783[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5154_3 (.CI(n32107), .I0(n9804[0]), .I1(n159_adj_4575), 
            .CO(n32108));
    SB_LUT4 add_5154_2_lut (.I0(GND_net), .I1(n17_adj_4576), .I2(n86_adj_4577), 
            .I3(GND_net), .O(n9783[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5154_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5154_2 (.CI(GND_net), .I0(n17_adj_4576), .I1(n86_adj_4577), 
            .CO(n32107));
    SB_LUT4 add_5153_21_lut (.I0(GND_net), .I1(n9783[18]), .I2(GND_net), 
            .I3(n32106), .O(n9761[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5153_20_lut (.I0(GND_net), .I1(n9783[17]), .I2(GND_net), 
            .I3(n32105), .O(n9761[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_20 (.CI(n32105), .I0(n9783[17]), .I1(GND_net), .CO(n32106));
    SB_LUT4 add_5153_19_lut (.I0(GND_net), .I1(n9783[16]), .I2(GND_net), 
            .I3(n32104), .O(n9761[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_19 (.CI(n32104), .I0(n9783[16]), .I1(GND_net), .CO(n32105));
    SB_LUT4 add_5153_18_lut (.I0(GND_net), .I1(n9783[15]), .I2(GND_net), 
            .I3(n32103), .O(n9761[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_18 (.CI(n32103), .I0(n9783[15]), .I1(GND_net), .CO(n32104));
    SB_LUT4 add_5153_17_lut (.I0(GND_net), .I1(n9783[14]), .I2(GND_net), 
            .I3(n32102), .O(n9761[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_17 (.CI(n32102), .I0(n9783[14]), .I1(GND_net), .CO(n32103));
    SB_LUT4 add_5153_16_lut (.I0(GND_net), .I1(n9783[13]), .I2(n1105_adj_4578), 
            .I3(n32101), .O(n9761[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_16 (.CI(n32101), .I0(n9783[13]), .I1(n1105_adj_4578), 
            .CO(n32102));
    SB_LUT4 add_5153_15_lut (.I0(GND_net), .I1(n9783[12]), .I2(n1032_adj_4579), 
            .I3(n32100), .O(n9761[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_15 (.CI(n32100), .I0(n9783[12]), .I1(n1032_adj_4579), 
            .CO(n32101));
    SB_LUT4 add_5153_14_lut (.I0(GND_net), .I1(n9783[11]), .I2(n959_adj_4580), 
            .I3(n32099), .O(n9761[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_14 (.CI(n32099), .I0(n9783[11]), .I1(n959_adj_4580), 
            .CO(n32100));
    SB_LUT4 add_5153_13_lut (.I0(GND_net), .I1(n9783[10]), .I2(n886_adj_4581), 
            .I3(n32098), .O(n9761[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_13 (.CI(n32098), .I0(n9783[10]), .I1(n886_adj_4581), 
            .CO(n32099));
    SB_LUT4 add_5153_12_lut (.I0(GND_net), .I1(n9783[9]), .I2(n813_adj_4582), 
            .I3(n32097), .O(n9761[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_12 (.CI(n32097), .I0(n9783[9]), .I1(n813_adj_4582), 
            .CO(n32098));
    SB_LUT4 add_5153_11_lut (.I0(GND_net), .I1(n9783[8]), .I2(n740_adj_4583), 
            .I3(n32096), .O(n9761[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_11 (.CI(n32096), .I0(n9783[8]), .I1(n740_adj_4583), 
            .CO(n32097));
    SB_LUT4 add_5153_10_lut (.I0(GND_net), .I1(n9783[7]), .I2(n667_adj_4584), 
            .I3(n32095), .O(n9761[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_10_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3489[2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_5153_10 (.CI(n32095), .I0(n9783[7]), .I1(n667_adj_4584), 
            .CO(n32096));
    SB_LUT4 add_5153_9_lut (.I0(GND_net), .I1(n9783[6]), .I2(n594_adj_4585), 
            .I3(n32094), .O(n9761[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_9 (.CI(n32094), .I0(n9783[6]), .I1(n594_adj_4585), 
            .CO(n32095));
    SB_LUT4 add_5153_8_lut (.I0(GND_net), .I1(n9783[5]), .I2(n521_adj_4586), 
            .I3(n32093), .O(n9761[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_8 (.CI(n32093), .I0(n9783[5]), .I1(n521_adj_4586), 
            .CO(n32094));
    SB_LUT4 add_5153_7_lut (.I0(GND_net), .I1(n9783[4]), .I2(n448_adj_4587), 
            .I3(n32092), .O(n9761[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1[23]), 
            .I3(n30922), .O(\PID_CONTROLLER.integral_23__N_3564 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_7 (.CI(n32092), .I0(n9783[4]), .I1(n448_adj_4587), 
            .CO(n32093));
    SB_LUT4 add_5153_6_lut (.I0(GND_net), .I1(n9783[3]), .I2(n375_adj_4589), 
            .I3(n32091), .O(n9761[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1[22]), .I3(n30921), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5313_5_lut (.I0(GND_net), .I1(n12912[2]), .I2(n320_adj_4591), 
            .I3(n30989), .O(n12717[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5313_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5313_5 (.CI(n30989), .I0(n12912[2]), .I1(n320_adj_4591), 
            .CO(n30990));
    SB_CARRY add_5153_6 (.CI(n32091), .I0(n9783[3]), .I1(n375_adj_4589), 
            .CO(n32092));
    SB_LUT4 add_5153_5_lut (.I0(GND_net), .I1(n9783[2]), .I2(n302_adj_4592), 
            .I3(n32090), .O(n9761[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_5 (.CI(n32090), .I0(n9783[2]), .I1(n302_adj_4592), 
            .CO(n32091));
    SB_LUT4 add_5153_4_lut (.I0(GND_net), .I1(n9783[1]), .I2(n229_adj_4593), 
            .I3(n32089), .O(n9761[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_4 (.CI(n32089), .I0(n9783[1]), .I1(n229_adj_4593), 
            .CO(n32090));
    SB_LUT4 add_5153_3_lut (.I0(GND_net), .I1(n9783[0]), .I2(n156_adj_4594), 
            .I3(n32088), .O(n9761[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_3 (.CI(n32088), .I0(n9783[0]), .I1(n156_adj_4594), 
            .CO(n32089));
    SB_LUT4 add_5153_2_lut (.I0(GND_net), .I1(n14_adj_4595), .I2(n83_adj_4596), 
            .I3(GND_net), .O(n9761[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5153_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5153_2 (.CI(GND_net), .I0(n14_adj_4595), .I1(n83_adj_4596), 
            .CO(n32088));
    SB_LUT4 add_5152_22_lut (.I0(GND_net), .I1(n9761[19]), .I2(GND_net), 
            .I3(n32087), .O(n9738[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5152_21_lut (.I0(GND_net), .I1(n9761[18]), .I2(GND_net), 
            .I3(n32086), .O(n9738[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_21 (.CI(n32086), .I0(n9761[18]), .I1(GND_net), .CO(n32087));
    SB_LUT4 add_5152_20_lut (.I0(GND_net), .I1(n9761[17]), .I2(GND_net), 
            .I3(n32085), .O(n9738[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_20 (.CI(n32085), .I0(n9761[17]), .I1(GND_net), .CO(n32086));
    SB_LUT4 add_5152_19_lut (.I0(GND_net), .I1(n9761[16]), .I2(GND_net), 
            .I3(n32084), .O(n9738[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_19 (.CI(n32084), .I0(n9761[16]), .I1(GND_net), .CO(n32085));
    SB_LUT4 add_5152_18_lut (.I0(GND_net), .I1(n9761[15]), .I2(GND_net), 
            .I3(n32083), .O(n9738[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_18 (.CI(n32083), .I0(n9761[15]), .I1(GND_net), .CO(n32084));
    SB_LUT4 add_5152_17_lut (.I0(GND_net), .I1(n9761[14]), .I2(GND_net), 
            .I3(n32082), .O(n9738[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_17 (.CI(n32082), .I0(n9761[14]), .I1(GND_net), .CO(n32083));
    SB_LUT4 add_5152_16_lut (.I0(GND_net), .I1(n9761[13]), .I2(n1102_adj_4597), 
            .I3(n32081), .O(n9738[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_16 (.CI(n32081), .I0(n9761[13]), .I1(n1102_adj_4597), 
            .CO(n32082));
    SB_LUT4 add_5152_15_lut (.I0(GND_net), .I1(n9761[12]), .I2(n1029_adj_4598), 
            .I3(n32080), .O(n9738[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_15 (.CI(n32080), .I0(n9761[12]), .I1(n1029_adj_4598), 
            .CO(n32081));
    SB_LUT4 add_5152_14_lut (.I0(GND_net), .I1(n9761[11]), .I2(n956_adj_4599), 
            .I3(n32079), .O(n9738[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_14 (.CI(n32079), .I0(n9761[11]), .I1(n956_adj_4599), 
            .CO(n32080));
    SB_LUT4 add_5152_13_lut (.I0(GND_net), .I1(n9761[10]), .I2(n883_adj_4600), 
            .I3(n32078), .O(n9738[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_13 (.CI(n32078), .I0(n9761[10]), .I1(n883_adj_4600), 
            .CO(n32079));
    SB_LUT4 add_5152_12_lut (.I0(GND_net), .I1(n9761[9]), .I2(n810_adj_4601), 
            .I3(n32077), .O(n9738[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_12 (.CI(n32077), .I0(n9761[9]), .I1(n810_adj_4601), 
            .CO(n32078));
    SB_LUT4 add_5152_11_lut (.I0(GND_net), .I1(n9761[8]), .I2(n737_adj_4602), 
            .I3(n32076), .O(n9738[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_11 (.CI(n32076), .I0(n9761[8]), .I1(n737_adj_4602), 
            .CO(n32077));
    SB_LUT4 add_5152_10_lut (.I0(GND_net), .I1(n9761[7]), .I2(n664_adj_4603), 
            .I3(n32075), .O(n9738[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_10 (.CI(n32075), .I0(n9761[7]), .I1(n664_adj_4603), 
            .CO(n32076));
    SB_LUT4 add_5152_9_lut (.I0(GND_net), .I1(n9761[6]), .I2(n591_adj_4604), 
            .I3(n32074), .O(n9738[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_9 (.CI(n32074), .I0(n9761[6]), .I1(n591_adj_4604), 
            .CO(n32075));
    SB_LUT4 add_5152_8_lut (.I0(GND_net), .I1(n9761[5]), .I2(n518_adj_4605), 
            .I3(n32073), .O(n9738[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_8 (.CI(n32073), .I0(n9761[5]), .I1(n518_adj_4605), 
            .CO(n32074));
    SB_LUT4 add_5152_7_lut (.I0(GND_net), .I1(n9761[4]), .I2(n445_adj_4606), 
            .I3(n32072), .O(n9738[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_7 (.CI(n32072), .I0(n9761[4]), .I1(n445_adj_4606), 
            .CO(n32073));
    SB_LUT4 add_5152_6_lut (.I0(GND_net), .I1(n9761[3]), .I2(n372_adj_4607), 
            .I3(n32071), .O(n9738[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_6 (.CI(n32071), .I0(n9761[3]), .I1(n372_adj_4607), 
            .CO(n32072));
    SB_LUT4 add_5152_5_lut (.I0(GND_net), .I1(n9761[2]), .I2(n299_adj_4608), 
            .I3(n32070), .O(n9738[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_5 (.CI(n32070), .I0(n9761[2]), .I1(n299_adj_4608), 
            .CO(n32071));
    SB_LUT4 add_5313_4_lut (.I0(GND_net), .I1(n12912[1]), .I2(n247_adj_4609), 
            .I3(n30988), .O(n12717[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5313_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5152_4_lut (.I0(GND_net), .I1(n9761[1]), .I2(n226_adj_4610), 
            .I3(n32069), .O(n9738[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_4 (.CI(n32069), .I0(n9761[1]), .I1(n226_adj_4610), 
            .CO(n32070));
    SB_CARRY add_723_11 (.CI(n30802), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n3141[9]), .CO(n30803));
    SB_LUT4 add_5152_3_lut (.I0(GND_net), .I1(n9761[0]), .I2(n153_adj_4611), 
            .I3(n32068), .O(n9738[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_3 (.CI(n32068), .I0(n9761[0]), .I1(n153_adj_4611), 
            .CO(n32069));
    SB_LUT4 add_723_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n3141[8]), .I3(n30801), .O(\PID_CONTROLLER.integral_23__N_3513 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5152_2_lut (.I0(GND_net), .I1(n11_adj_4612), .I2(n80_adj_4613), 
            .I3(GND_net), .O(n9738[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5152_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5152_2 (.CI(GND_net), .I0(n11_adj_4612), .I1(n80_adj_4613), 
            .CO(n32068));
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3513 [23]), 
            .I1(n9714[21]), .I2(GND_net), .I3(n32067), .O(n7900[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5313_4 (.CI(n30988), .I0(n12912[1]), .I1(n247_adj_4609), 
            .CO(n30989));
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n9714[20]), .I2(GND_net), 
            .I3(n32066), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_23 (.CI(n32066), .I0(n9714[20]), .I1(GND_net), 
            .CO(n32067));
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n9714[19]), .I2(GND_net), 
            .I3(n32065), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_22 (.CI(n32065), .I0(n9714[19]), .I1(GND_net), 
            .CO(n32066));
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n9714[18]), .I2(GND_net), 
            .I3(n32064), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_21 (.CI(n32064), .I0(n9714[18]), .I1(GND_net), 
            .CO(n32065));
    SB_LUT4 add_5313_3_lut (.I0(GND_net), .I1(n12912[0]), .I2(n174_adj_4614), 
            .I3(n30987), .O(n12717[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5313_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n9714[17]), .I2(GND_net), 
            .I3(n32063), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n30921), .I0(GND_net), .I1(n1[22]), 
            .CO(n30922));
    SB_CARRY mult_11_add_1225_20 (.CI(n32063), .I0(n9714[17]), .I1(GND_net), 
            .CO(n32064));
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n9714[16]), .I2(GND_net), 
            .I3(n32062), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_19 (.CI(n32062), .I0(n9714[16]), .I1(GND_net), 
            .CO(n32063));
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n9714[15]), .I2(GND_net), 
            .I3(n32061), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5313_3 (.CI(n30987), .I0(n12912[0]), .I1(n174_adj_4614), 
            .CO(n30988));
    SB_CARRY mult_11_add_1225_18 (.CI(n32061), .I0(n9714[15]), .I1(GND_net), 
            .CO(n32062));
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n9714[14]), .I2(GND_net), 
            .I3(n32060), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_17 (.CI(n32060), .I0(n9714[14]), .I1(GND_net), 
            .CO(n32061));
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n9714[13]), .I2(n1096_adj_4615), 
            .I3(n32059), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_16 (.CI(n32059), .I0(n9714[13]), .I1(n1096_adj_4615), 
            .CO(n32060));
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n9714[12]), .I2(n1023_adj_4616), 
            .I3(n32058), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_723_10 (.CI(n30801), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n3141[8]), .CO(n30802));
    SB_CARRY mult_11_add_1225_15 (.CI(n32058), .I0(n9714[12]), .I1(n1023_adj_4616), 
            .CO(n32059));
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n9714[11]), .I2(n950_adj_4617), 
            .I3(n32057), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_7 (.CI(n30721), .I0(n106[5]), .I1(n155[5]), .CO(n30722));
    SB_CARRY mult_11_add_1225_14 (.CI(n32057), .I0(n9714[11]), .I1(n950_adj_4617), 
            .CO(n32058));
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n9714[10]), .I2(n877), 
            .I3(n32056), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_13 (.CI(n32056), .I0(n9714[10]), .I1(n877), 
            .CO(n32057));
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n9714[9]), .I2(n804), 
            .I3(n32055), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_12 (.CI(n32055), .I0(n9714[9]), .I1(n804), 
            .CO(n32056));
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n9714[8]), .I2(n731), 
            .I3(n32054), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_11 (.CI(n32054), .I0(n9714[8]), .I1(n731), 
            .CO(n32055));
    SB_LUT4 add_723_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n3141[7]), .I3(n30800), .O(\PID_CONTROLLER.integral_23__N_3513 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n9714[7]), .I2(n658_adj_4618), 
            .I3(n32053), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n32053), .I0(n9714[7]), .I1(n658_adj_4618), 
            .CO(n32054));
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n9714[6]), .I2(n585_adj_4619), 
            .I3(n32052), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_9 (.CI(n32052), .I0(n9714[6]), .I1(n585_adj_4619), 
            .CO(n32053));
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n9714[5]), .I2(n512_adj_4620), 
            .I3(n32051), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_8 (.CI(n32051), .I0(n9714[5]), .I1(n512_adj_4620), 
            .CO(n32052));
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n9714[4]), .I2(n439_adj_4621), 
            .I3(n32050), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_7 (.CI(n32050), .I0(n9714[4]), .I1(n439_adj_4621), 
            .CO(n32051));
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n9714[3]), .I2(n366_adj_4622), 
            .I3(n32049), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_6_lut (.I0(GND_net), .I1(n106[4]), .I2(n155[4]), .I3(n30720), 
            .O(duty_23__N_3613[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_6 (.CI(n32049), .I0(n9714[3]), .I1(n366_adj_4622), 
            .CO(n32050));
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n9714[2]), .I2(n293_adj_4623), 
            .I3(n32048), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_5 (.CI(n32048), .I0(n9714[2]), .I1(n293_adj_4623), 
            .CO(n32049));
    SB_CARRY add_12_6 (.CI(n30720), .I0(n106[4]), .I1(n155[4]), .CO(n30721));
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n9714[1]), .I2(n220_adj_4624), 
            .I3(n32047), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_4 (.CI(n32047), .I0(n9714[1]), .I1(n220_adj_4624), 
            .CO(n32048));
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n9714[0]), .I2(n147_adj_4625), 
            .I3(n32046), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n32046), .I0(n9714[0]), .I1(n147_adj_4625), 
            .CO(n32047));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4626), .I2(n74_adj_4627), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_4626), .I1(n74_adj_4627), 
            .CO(n32046));
    SB_LUT4 add_5151_23_lut (.I0(GND_net), .I1(n9738[20]), .I2(GND_net), 
            .I3(n32045), .O(n9714[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5151_22_lut (.I0(GND_net), .I1(n9738[19]), .I2(GND_net), 
            .I3(n32044), .O(n9714[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_22 (.CI(n32044), .I0(n9738[19]), .I1(GND_net), .CO(n32045));
    SB_LUT4 add_5151_21_lut (.I0(GND_net), .I1(n9738[18]), .I2(GND_net), 
            .I3(n32043), .O(n9714[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_21 (.CI(n32043), .I0(n9738[18]), .I1(GND_net), .CO(n32044));
    SB_LUT4 add_5151_20_lut (.I0(GND_net), .I1(n9738[17]), .I2(GND_net), 
            .I3(n32042), .O(n9714[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_20_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3489[3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3489[4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3489[5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3489[6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3489[7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3489[8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3489[9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3489[10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3489[11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3489[12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3489[13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3489[14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3489[15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3489[16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3489[17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3489[18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3489[19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3489[20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3489[21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3489[22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3489[23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i1  (.Q(\PID_CONTROLLER.integral [1]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i2  (.Q(\PID_CONTROLLER.integral [2]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i3  (.Q(\PID_CONTROLLER.integral [3]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i4  (.Q(\PID_CONTROLLER.integral [4]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i5  (.Q(\PID_CONTROLLER.integral [5]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i6  (.Q(\PID_CONTROLLER.integral [6]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i7  (.Q(\PID_CONTROLLER.integral [7]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i8  (.Q(\PID_CONTROLLER.integral [8]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i9  (.Q(\PID_CONTROLLER.integral [9]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i10  (.Q(\PID_CONTROLLER.integral [10]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i11  (.Q(\PID_CONTROLLER.integral [11]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i12  (.Q(\PID_CONTROLLER.integral [12]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i13  (.Q(\PID_CONTROLLER.integral [13]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i14  (.Q(\PID_CONTROLLER.integral [14]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i15  (.Q(\PID_CONTROLLER.integral [15]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i16  (.Q(\PID_CONTROLLER.integral [16]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i17  (.Q(\PID_CONTROLLER.integral [17]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i18  (.Q(\PID_CONTROLLER.integral [18]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i19  (.Q(\PID_CONTROLLER.integral [19]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i20  (.Q(\PID_CONTROLLER.integral [20]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i21  (.Q(\PID_CONTROLLER.integral [21]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i22  (.Q(\PID_CONTROLLER.integral [22]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i23  (.Q(\PID_CONTROLLER.integral [23]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3513 [23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_5151_20 (.CI(n32042), .I0(n9738[17]), .I1(GND_net), .CO(n32043));
    SB_LUT4 add_5151_19_lut (.I0(GND_net), .I1(n9738[16]), .I2(GND_net), 
            .I3(n32041), .O(n9714[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_19 (.CI(n32041), .I0(n9738[16]), .I1(GND_net), .CO(n32042));
    SB_LUT4 add_5151_18_lut (.I0(GND_net), .I1(n9738[15]), .I2(GND_net), 
            .I3(n32040), .O(n9714[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_18 (.CI(n32040), .I0(n9738[15]), .I1(GND_net), .CO(n32041));
    SB_LUT4 add_5151_17_lut (.I0(GND_net), .I1(n9738[14]), .I2(GND_net), 
            .I3(n32039), .O(n9714[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_17 (.CI(n32039), .I0(n9738[14]), .I1(GND_net), .CO(n32040));
    SB_LUT4 add_5151_16_lut (.I0(GND_net), .I1(n9738[13]), .I2(n1099_adj_4628), 
            .I3(n32038), .O(n9714[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_16 (.CI(n32038), .I0(n9738[13]), .I1(n1099_adj_4628), 
            .CO(n32039));
    SB_LUT4 add_5151_15_lut (.I0(GND_net), .I1(n9738[12]), .I2(n1026_adj_4629), 
            .I3(n32037), .O(n9714[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_15 (.CI(n32037), .I0(n9738[12]), .I1(n1026_adj_4629), 
            .CO(n32038));
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19129_2_lut (.I0(n28[2]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[2]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19129_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_4631));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5151_14_lut (.I0(GND_net), .I1(n9738[11]), .I2(n953_adj_4632), 
            .I3(n32036), .O(n9714[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_14 (.CI(n32036), .I0(n9738[11]), .I1(n953_adj_4632), 
            .CO(n32037));
    SB_LUT4 add_5151_13_lut (.I0(GND_net), .I1(n9738[10]), .I2(n880_adj_4633), 
            .I3(n32035), .O(n9714[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_13 (.CI(n32035), .I0(n9738[10]), .I1(n880_adj_4633), 
            .CO(n32036));
    SB_LUT4 add_5151_12_lut (.I0(GND_net), .I1(n9738[9]), .I2(n807_adj_4634), 
            .I3(n32034), .O(n9714[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1[21]), .I3(n30920), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5151_12 (.CI(n32034), .I0(n9738[9]), .I1(n807_adj_4634), 
            .CO(n32035));
    SB_LUT4 add_5151_11_lut (.I0(GND_net), .I1(n9738[8]), .I2(n734_adj_4636), 
            .I3(n32033), .O(n9714[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_11 (.CI(n32033), .I0(n9738[8]), .I1(n734_adj_4636), 
            .CO(n32034));
    SB_LUT4 add_5313_2_lut (.I0(GND_net), .I1(n32_adj_4637), .I2(n101_adj_4638), 
            .I3(GND_net), .O(n12717[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5313_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_23 (.CI(n30920), .I0(GND_net), .I1(n1[21]), 
            .CO(n30921));
    SB_LUT4 add_5151_10_lut (.I0(GND_net), .I1(n9738[7]), .I2(n661_adj_4639), 
            .I3(n32032), .O(n9714[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_723_9 (.CI(n30800), .I0(\PID_CONTROLLER.integral [7]), 
            .I1(n3141[7]), .CO(n30801));
    SB_CARRY add_5151_10 (.CI(n32032), .I0(n9738[7]), .I1(n661_adj_4639), 
            .CO(n32033));
    SB_LUT4 add_5151_9_lut (.I0(GND_net), .I1(n9738[6]), .I2(n588_adj_4640), 
            .I3(n32031), .O(n9714[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_9 (.CI(n32031), .I0(n9738[6]), .I1(n588_adj_4640), 
            .CO(n32032));
    SB_LUT4 add_5151_8_lut (.I0(GND_net), .I1(n9738[5]), .I2(n515_adj_4641), 
            .I3(n32030), .O(n9714[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_8 (.CI(n32030), .I0(n9738[5]), .I1(n515_adj_4641), 
            .CO(n32031));
    SB_LUT4 add_5151_7_lut (.I0(GND_net), .I1(n9738[4]), .I2(n442_adj_4642), 
            .I3(n32029), .O(n9714[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_7 (.CI(n32029), .I0(n9738[4]), .I1(n442_adj_4642), 
            .CO(n32030));
    SB_LUT4 add_5151_6_lut (.I0(GND_net), .I1(n9738[3]), .I2(n369_adj_4643), 
            .I3(n32028), .O(n9714[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_6 (.CI(n32028), .I0(n9738[3]), .I1(n369_adj_4643), 
            .CO(n32029));
    SB_LUT4 add_5151_5_lut (.I0(GND_net), .I1(n9738[2]), .I2(n296_adj_4644), 
            .I3(n32027), .O(n9714[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_5 (.CI(n32027), .I0(n9738[2]), .I1(n296_adj_4644), 
            .CO(n32028));
    SB_LUT4 add_5151_4_lut (.I0(GND_net), .I1(n9738[1]), .I2(n223_adj_4645), 
            .I3(n32026), .O(n9714[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_4 (.CI(n32026), .I0(n9738[1]), .I1(n223_adj_4645), 
            .CO(n32027));
    SB_LUT4 add_723_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n3141[6]), .I3(n30799), .O(\PID_CONTROLLER.integral_23__N_3513 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5151_3_lut (.I0(GND_net), .I1(n9738[0]), .I2(n150_adj_4646), 
            .I3(n32025), .O(n9714[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_5_lut (.I0(GND_net), .I1(n106[3]), .I2(n155[3]), .I3(n30719), 
            .O(duty_23__N_3613[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_3 (.CI(n32025), .I0(n9738[0]), .I1(n150_adj_4646), 
            .CO(n32026));
    SB_LUT4 add_5151_2_lut (.I0(GND_net), .I1(n8_adj_4647), .I2(n77_adj_4648), 
            .I3(GND_net), .O(n9714[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5151_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5151_2 (.CI(GND_net), .I0(n8_adj_4647), .I1(n77_adj_4648), 
            .CO(n32025));
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1[20]), .I3(n30919), .O(n41_adj_4422)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_723_8 (.CI(n30799), .I0(\PID_CONTROLLER.integral [6]), 
            .I1(n3141[6]), .CO(n30800));
    SB_LUT4 add_723_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n3141[5]), .I3(n30798), .O(\PID_CONTROLLER.integral_23__N_3513 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_723_7 (.CI(n30798), .I0(\PID_CONTROLLER.integral [5]), 
            .I1(n3141[5]), .CO(n30799));
    SB_CARRY add_5313_2 (.CI(GND_net), .I0(n32_adj_4637), .I1(n101_adj_4638), 
            .CO(n30987));
    SB_CARRY unary_minus_5_add_3_22 (.CI(n30919), .I0(GND_net), .I1(n1[20]), 
            .CO(n30920));
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1[19]), .I3(n30918), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n30918), .I0(GND_net), .I1(n1[19]), 
            .CO(n30919));
    SB_LUT4 add_5326_14_lut (.I0(GND_net), .I1(n13080[11]), .I2(n980_adj_4651), 
            .I3(n30986), .O(n12912[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1[18]), .I3(n30917), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615_adj_4653));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_10_add_1225_11 (.CI(n31508), .I0(n9589[8]), .I1(n731_adj_4655), 
            .CO(n31509));
    SB_LUT4 add_723_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n3141[4]), .I3(n30797), .O(\PID_CONTROLLER.integral_23__N_3513 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5326_13_lut (.I0(GND_net), .I1(n13080[10]), .I2(n907_adj_4656), 
            .I3(n30985), .O(n12912[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n30917), .I0(GND_net), .I1(n1[18]), 
            .CO(n30918));
    SB_LUT4 mult_10_add_1225_11_lut (.I0(GND_net), .I1(n9589[8]), .I2(n731_adj_4655), 
            .I3(n31508), .O(n106[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_5 (.CI(n30719), .I0(n106[3]), .I1(n155[3]), .CO(n30720));
    SB_CARRY add_5326_13 (.CI(n30985), .I0(n13080[10]), .I1(n907_adj_4656), 
            .CO(n30986));
    SB_LUT4 add_5326_12_lut (.I0(GND_net), .I1(n13080[9]), .I2(n834_adj_4657), 
            .I3(n30984), .O(n12912[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688_adj_4658));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_10_add_1225_12 (.CI(n31509), .I0(n9589[9]), .I1(n804_adj_4660), 
            .CO(n31510));
    SB_LUT4 mult_10_add_1225_12_lut (.I0(GND_net), .I1(n9589[9]), .I2(n804_adj_4660), 
            .I3(n31509), .O(n106[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_13 (.CI(n31510), .I0(n9589[10]), .I1(n877_adj_4661), 
            .CO(n31511));
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1[17]), .I3(n30916), .O(n35_adj_4405)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_723_6 (.CI(n30797), .I0(\PID_CONTROLLER.integral [4]), 
            .I1(n3141[4]), .CO(n30798));
    SB_LUT4 mult_10_add_1225_13_lut (.I0(GND_net), .I1(n9589[10]), .I2(n877_adj_4661), 
            .I3(n31510), .O(n106[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_4_lut (.I0(GND_net), .I1(n106[2]), .I2(n155[2]), .I3(n30718), 
            .O(duty_23__N_3613[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_12 (.CI(n30984), .I0(n13080[9]), .I1(n834_adj_4657), 
            .CO(n30985));
    SB_LUT4 add_5349_12_lut (.I0(GND_net), .I1(n13343[9]), .I2(n840_adj_4663), 
            .I3(n32002), .O(n13223[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5349_11_lut (.I0(GND_net), .I1(n13343[8]), .I2(n767_adj_4664), 
            .I3(n32001), .O(n13223[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5349_11 (.CI(n32001), .I0(n13343[8]), .I1(n767_adj_4664), 
            .CO(n32002));
    SB_CARRY mult_10_add_1225_14 (.CI(n31511), .I0(n9589[11]), .I1(n950), 
            .CO(n31512));
    SB_LUT4 add_5349_10_lut (.I0(GND_net), .I1(n13343[7]), .I2(n694_adj_4665), 
            .I3(n32000), .O(n13223[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5349_10 (.CI(n32000), .I0(n13343[7]), .I1(n694_adj_4665), 
            .CO(n32001));
    SB_LUT4 add_5349_9_lut (.I0(GND_net), .I1(n13343[6]), .I2(n621_adj_4666), 
            .I3(n31999), .O(n13223[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5349_9 (.CI(n31999), .I0(n13343[6]), .I1(n621_adj_4666), 
            .CO(n32000));
    SB_LUT4 add_5349_8_lut (.I0(GND_net), .I1(n13343[5]), .I2(n548_adj_4667), 
            .I3(n31998), .O(n13223[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5349_8 (.CI(n31998), .I0(n13343[5]), .I1(n548_adj_4667), 
            .CO(n31999));
    SB_LUT4 add_5349_7_lut (.I0(GND_net), .I1(n13343[4]), .I2(n475_adj_4668), 
            .I3(n31997), .O(n13223[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5349_7 (.CI(n31997), .I0(n13343[4]), .I1(n475_adj_4668), 
            .CO(n31998));
    SB_CARRY unary_minus_5_add_3_19 (.CI(n30916), .I0(GND_net), .I1(n1[17]), 
            .CO(n30917));
    SB_LUT4 add_5349_6_lut (.I0(GND_net), .I1(n13343[3]), .I2(n402_adj_4669), 
            .I3(n31996), .O(n13223[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1[16]), .I3(n30915), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5349_6 (.CI(n31996), .I0(n13343[3]), .I1(n402_adj_4669), 
            .CO(n31997));
    SB_LUT4 add_5349_5_lut (.I0(GND_net), .I1(n13343[2]), .I2(n329_adj_4671), 
            .I3(n31995), .O(n13223[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5349_5 (.CI(n31995), .I0(n13343[2]), .I1(n329_adj_4671), 
            .CO(n31996));
    SB_LUT4 add_723_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n3141[3]), .I3(n30796), .O(\PID_CONTROLLER.integral_23__N_3513 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5349_4_lut (.I0(GND_net), .I1(n13343[1]), .I2(n256_adj_4672), 
            .I3(n31994), .O(n13223[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5349_4 (.CI(n31994), .I0(n13343[1]), .I1(n256_adj_4672), 
            .CO(n31995));
    SB_LUT4 add_5349_3_lut (.I0(GND_net), .I1(n13343[0]), .I2(n183_adj_4673), 
            .I3(n31993), .O(n13223[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5349_3 (.CI(n31993), .I0(n13343[0]), .I1(n183_adj_4673), 
            .CO(n31994));
    SB_LUT4 add_5349_2_lut (.I0(GND_net), .I1(n41_adj_4674), .I2(n110_adj_4675), 
            .I3(GND_net), .O(n13223[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5349_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5349_2 (.CI(GND_net), .I0(n41_adj_4674), .I1(n110_adj_4675), 
            .CO(n31993));
    SB_LUT4 add_5326_11_lut (.I0(GND_net), .I1(n13080[8]), .I2(n761_adj_4676), 
            .I3(n30983), .O(n12912[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n30915), .I0(GND_net), .I1(n1[16]), 
            .CO(n30916));
    SB_CARRY add_5326_11 (.CI(n30983), .I0(n13080[8]), .I1(n761_adj_4676), 
            .CO(n30984));
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1[15]), .I3(n30914), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5326_10_lut (.I0(GND_net), .I1(n13080[7]), .I2(n688_adj_4658), 
            .I3(n30982), .O(n12912[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_17 (.CI(n30914), .I0(GND_net), .I1(n1[15]), 
            .CO(n30915));
    SB_CARRY add_723_5 (.CI(n30796), .I0(\PID_CONTROLLER.integral [3]), 
            .I1(n3141[3]), .CO(n30797));
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1[14]), .I3(n30913), .O(n29_adj_4404)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5326_10 (.CI(n30982), .I0(n13080[7]), .I1(n688_adj_4658), 
            .CO(n30983));
    SB_LUT4 add_5326_9_lut (.I0(GND_net), .I1(n13080[6]), .I2(n615_adj_4653), 
            .I3(n30981), .O(n12912[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_9 (.CI(n30981), .I0(n13080[6]), .I1(n615_adj_4653), 
            .CO(n30982));
    SB_CARRY unary_minus_5_add_3_16 (.CI(n30913), .I0(GND_net), .I1(n1[14]), 
            .CO(n30914));
    SB_CARRY add_12_4 (.CI(n30718), .I0(n106[2]), .I1(n155[2]), .CO(n30719));
    SB_LUT4 add_5326_8_lut (.I0(GND_net), .I1(n13080[5]), .I2(n542_adj_4631), 
            .I3(n30980), .O(n12912[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_8 (.CI(n30980), .I0(n13080[5]), .I1(n542_adj_4631), 
            .CO(n30981));
    SB_LUT4 add_723_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n3141[2]), .I3(n30795), .O(\PID_CONTROLLER.integral_23__N_3513 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_723_4 (.CI(n30795), .I0(\PID_CONTROLLER.integral [2]), 
            .I1(n3141[2]), .CO(n30796));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1[13]), .I3(n30912), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761_adj_4676));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110_adj_4675));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(n28[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4674));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183_adj_4673));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4672));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19130_2_lut (.I0(n28[3]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[3]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_4671));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_4669));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4668));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_4667));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_4666));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5326_7_lut (.I0(GND_net), .I1(n13080[4]), .I2(n469_adj_4566), 
            .I3(n30979), .O(n12912[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_4665));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_4664));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(n28[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_4663));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n30912), .I0(GND_net), .I1(n1[13]), 
            .CO(n30913));
    SB_LUT4 add_12_3_lut (.I0(GND_net), .I1(n106[1]), .I2(n155[1]), .I3(n30717), 
            .O(duty_23__N_3613[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1[12]), .I3(n30911), .O(n25_adj_4402)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_723_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n3141[1]), .I3(n30794), .O(\PID_CONTROLLER.integral_23__N_3513 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_7 (.CI(n30979), .I0(n13080[4]), .I1(n469_adj_4566), 
            .CO(n30980));
    SB_CARRY add_723_3 (.CI(n30794), .I0(\PID_CONTROLLER.integral [1]), 
            .I1(n3141[1]), .CO(n30795));
    SB_CARRY add_12_3 (.CI(n30717), .I0(n106[1]), .I1(n155[1]), .CO(n30718));
    SB_LUT4 add_12_2_lut (.I0(GND_net), .I1(n106[0]), .I2(n155[0]), .I3(GND_net), 
            .O(duty_23__N_3613[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n30911), .I0(GND_net), .I1(n1[12]), 
            .CO(n30912));
    SB_LUT4 add_5326_6_lut (.I0(GND_net), .I1(n13080[3]), .I2(n396_adj_4451), 
            .I3(n30978), .O(n12912[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1[11]), .I3(n30910), .O(n23_adj_4403)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877_adj_4661));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_723_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n3141[0]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3513 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_723_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n30910), .I0(GND_net), .I1(n1[11]), 
            .CO(n30911));
    SB_CARRY add_5326_6 (.CI(n30978), .I0(n13080[3]), .I1(n396_adj_4451), 
            .CO(n30979));
    SB_CARRY add_723_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n3141[0]), .CO(n30794));
    SB_LUT4 add_5326_5_lut (.I0(GND_net), .I1(n13080[2]), .I2(n323_adj_4444), 
            .I3(n30977), .O(n12912[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_5 (.CI(n30977), .I0(n13080[2]), .I1(n323_adj_4444), 
            .CO(n30978));
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1[10]), .I3(n30909), .O(n21_adj_4396)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804_adj_4660));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_2 (.CI(GND_net), .I0(n106[0]), .I1(n155[0]), .CO(n30717));
    SB_LUT4 add_5389_7_lut (.I0(GND_net), .I1(n37173), .I2(n490_adj_4429), 
            .I3(n30845), .O(n13633[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5389_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5326_4_lut (.I0(GND_net), .I1(n13080[1]), .I2(n250_adj_4426), 
            .I3(n30976), .O(n12912[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_4 (.CI(n30976), .I0(n13080[1]), .I1(n250_adj_4426), 
            .CO(n30977));
    SB_LUT4 add_5326_3_lut (.I0(GND_net), .I1(n13080[0]), .I2(n177_adj_4425), 
            .I3(n30975), .O(n12912[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5389_6_lut (.I0(GND_net), .I1(n13668[3]), .I2(n417_adj_4419), 
            .I3(n30844), .O(n13633[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5389_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_3 (.CI(n30975), .I0(n13080[0]), .I1(n177_adj_4425), 
            .CO(n30976));
    SB_CARRY add_5389_6 (.CI(n30844), .I0(n13668[3]), .I1(n417_adj_4419), 
            .CO(n30845));
    SB_CARRY unary_minus_5_add_3_12 (.CI(n30909), .I0(GND_net), .I1(n1[10]), 
            .CO(n30910));
    SB_LUT4 add_5389_5_lut (.I0(GND_net), .I1(n13668[2]), .I2(n344_adj_4415), 
            .I3(n30843), .O(n13633[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5389_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1[9]), .I3(n30908), .O(n19_adj_4397)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i29353_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3613[21]), 
            .I2(PWMLimit[9]), .I3(duty_23__N_3613[9]), .O(n39381));
    defparam i29353_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_5389_5 (.CI(n30843), .I0(n13668[2]), .I1(n344_adj_4415), 
            .CO(n30844));
    SB_LUT4 add_5389_4_lut (.I0(GND_net), .I1(n13668[1]), .I2(n271_adj_4376), 
            .I3(n30842), .O(n13633[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5389_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29364_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3613[16]), 
            .I2(PWMLimit[7]), .I3(duty_23__N_3613[7]), .O(n39392));
    defparam i29364_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i29317_2_lut_4_lut (.I0(duty_23__N_3613[21]), .I1(n257[21]), 
            .I2(duty_23__N_3613[9]), .I3(n257[9]), .O(n39345));
    defparam i29317_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834_adj_4657));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907_adj_4656));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5368_10_lut (.I0(GND_net), .I1(n13522[7]), .I2(n700_adj_4374), 
            .I3(n31088), .O(n13442[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5368_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19131_2_lut (.I0(n28[4]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[4]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19131_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731_adj_4655));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5368_9_lut (.I0(GND_net), .I1(n13522[6]), .I2(n627_adj_4373), 
            .I3(n31087), .O(n13442[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5368_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29327_2_lut_4_lut (.I0(duty_23__N_3613[16]), .I1(n257[16]), 
            .I2(duty_23__N_3613[7]), .I3(n257[7]), .O(n39355));
    defparam i29327_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_5368_9 (.CI(n31087), .I0(n13522[6]), .I1(n627_adj_4373), 
            .CO(n31088));
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980_adj_4651));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5368_8_lut (.I0(GND_net), .I1(n13522[5]), .I2(n554_adj_4372), 
            .I3(n31086), .O(n13442[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5368_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5368_8 (.CI(n31086), .I0(n13522[5]), .I1(n554_adj_4372), 
            .CO(n31087));
    SB_LUT4 add_5368_7_lut (.I0(GND_net), .I1(n13522[4]), .I2(n481), .I3(n31085), 
            .O(n13442[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5368_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5368_7 (.CI(n31085), .I0(n13522[4]), .I1(n481), .CO(n31086));
    SB_LUT4 add_5368_6_lut (.I0(GND_net), .I1(n13522[3]), .I2(n408), .I3(n31084), 
            .O(n13442[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5368_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5368_6 (.CI(n31084), .I0(n13522[3]), .I1(n408), .CO(n31085));
    SB_LUT4 add_5368_5_lut (.I0(GND_net), .I1(n13522[2]), .I2(n335), .I3(n31083), 
            .O(n13442[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5368_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5368_5 (.CI(n31083), .I0(n13522[2]), .I1(n335), .CO(n31084));
    SB_LUT4 add_5368_4_lut (.I0(GND_net), .I1(n13522[1]), .I2(n262), .I3(n31082), 
            .O(n13442[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5368_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5368_4 (.CI(n31082), .I0(n13522[1]), .I1(n262), .CO(n31083));
    SB_LUT4 add_5368_3_lut (.I0(GND_net), .I1(n13522[0]), .I2(n189), .I3(n31081), 
            .O(n13442[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5368_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5368_3 (.CI(n31081), .I0(n13522[0]), .I1(n189), .CO(n31082));
    SB_LUT4 add_5368_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n13442[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5368_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5368_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n31081));
    SB_LUT4 add_5269_18_lut (.I0(GND_net), .I1(n12255[15]), .I2(GND_net), 
            .I3(n31080), .O(n11968[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29389_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3613[3]), 
            .I2(duty_23__N_3613[2]), .I3(PWMLimit[2]), .O(n39417));   // verilog/motorControl.v(36[10:25])
    defparam i29389_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_5269_17_lut (.I0(GND_net), .I1(n12255[14]), .I2(GND_net), 
            .I3(n31079), .O(n11968[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_831_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3613[3]), 
            .I2(duty_23__N_3613[2]), .I3(GND_net), .O(n6_adj_4508));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_831_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_CARRY add_5269_17 (.CI(n31079), .I0(n12255[14]), .I1(GND_net), 
            .CO(n31080));
    SB_LUT4 add_5269_16_lut (.I0(GND_net), .I1(n12255[13]), .I2(n1114), 
            .I3(n31078), .O(n11968[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_16 (.CI(n31078), .I0(n12255[13]), .I1(n1114), .CO(n31079));
    SB_LUT4 add_5326_2_lut (.I0(GND_net), .I1(n35_adj_4321), .I2(n104_adj_4319), 
            .I3(GND_net), .O(n12912[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5326_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5269_15_lut (.I0(GND_net), .I1(n12255[12]), .I2(n1041), 
            .I3(n31077), .O(n11968[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_15 (.CI(n31077), .I0(n12255[12]), .I1(n1041), .CO(n31078));
    SB_LUT4 add_5269_14_lut (.I0(GND_net), .I1(n12255[11]), .I2(n968), 
            .I3(n31076), .O(n11968[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_14 (.CI(n31076), .I0(n12255[11]), .I1(n968), .CO(n31077));
    SB_CARRY unary_minus_5_add_3_11 (.CI(n30908), .I0(GND_net), .I1(n1[9]), 
            .CO(n30909));
    SB_LUT4 add_5269_13_lut (.I0(GND_net), .I1(n12255[10]), .I2(n895), 
            .I3(n31075), .O(n11968[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_13 (.CI(n31075), .I0(n12255[10]), .I1(n895), .CO(n31076));
    SB_CARRY add_5389_4 (.CI(n30842), .I0(n13668[1]), .I1(n271_adj_4376), 
            .CO(n30843));
    SB_LUT4 add_5269_12_lut (.I0(GND_net), .I1(n12255[9]), .I2(n822), 
            .I3(n31074), .O(n11968[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19132_2_lut (.I0(n28[5]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[5]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19132_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5269_12 (.CI(n31074), .I0(n12255[9]), .I1(n822), .CO(n31075));
    SB_LUT4 add_5269_11_lut (.I0(GND_net), .I1(n12255[8]), .I2(n749), 
            .I3(n31073), .O(n11968[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_11 (.CI(n31073), .I0(n12255[8]), .I1(n749), .CO(n31074));
    SB_LUT4 add_5269_10_lut (.I0(GND_net), .I1(n12255[7]), .I2(n676), 
            .I3(n31072), .O(n11968[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_10 (.CI(n31072), .I0(n12255[7]), .I1(n676), .CO(n31073));
    SB_LUT4 add_5269_9_lut (.I0(GND_net), .I1(n12255[6]), .I2(n603), .I3(n31071), 
            .O(n11968[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_9 (.CI(n31071), .I0(n12255[6]), .I1(n603), .CO(n31072));
    SB_LUT4 add_5269_8_lut (.I0(GND_net), .I1(n12255[5]), .I2(n530), .I3(n31070), 
            .O(n11968[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29351_3_lut_4_lut (.I0(duty_23__N_3613[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty_23__N_3613[2]), .O(n39379));   // verilog/motorControl.v(38[19:35])
    defparam i29351_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_CARRY add_5269_8 (.CI(n31070), .I0(n12255[5]), .I1(n530), .CO(n31071));
    SB_LUT4 add_5389_3_lut (.I0(GND_net), .I1(n13668[0]), .I2(n198), .I3(n30841), 
            .O(n13633[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5389_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5269_7_lut (.I0(GND_net), .I1(n12255[4]), .I2(n457), .I3(n31069), 
            .O(n11968[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_7 (.CI(n31069), .I0(n12255[4]), .I1(n457), .CO(n31070));
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty_23__N_3613[3]), .I1(n257[3]), 
            .I2(n257[2]), .I3(GND_net), .O(n6_adj_4480));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 add_5269_6_lut (.I0(GND_net), .I1(n12255[3]), .I2(n384), .I3(n31068), 
            .O(n11968[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_6 (.CI(n31068), .I0(n12255[3]), .I1(n384), .CO(n31069));
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1[8]), .I3(n30907), .O(n17_adj_4398)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5269_5_lut (.I0(GND_net), .I1(n12255[2]), .I2(n311), .I3(n31067), 
            .O(n11968[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5269_5 (.CI(n31067), .I0(n12255[2]), .I1(n311), .CO(n31068));
    SB_LUT4 add_5269_4_lut (.I0(GND_net), .I1(n12255[1]), .I2(n238), .I3(n31066), 
            .O(n11968[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n30907), .I0(GND_net), .I1(n1[8]), 
            .CO(n30908));
    SB_CARRY add_5269_4 (.CI(n31066), .I0(n12255[1]), .I1(n238), .CO(n31067));
    SB_LUT4 add_5269_3_lut (.I0(GND_net), .I1(n12255[0]), .I2(n165), .I3(n31065), 
            .O(n11968[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5326_2 (.CI(GND_net), .I0(n35_adj_4321), .I1(n104_adj_4319), 
            .CO(n30975));
    SB_CARRY add_5269_3 (.CI(n31065), .I0(n12255[0]), .I1(n165), .CO(n31066));
    SB_LUT4 add_5269_2_lut (.I0(GND_net), .I1(n23), .I2(n92), .I3(GND_net), 
            .O(n11968[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5269_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5269_2 (.CI(GND_net), .I0(n23), .I1(n92), .CO(n31065));
    SB_CARRY add_5389_3 (.CI(n30841), .I0(n13668[0]), .I1(n198), .CO(n30842));
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_4648));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4647));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1[7]), .I3(n30906), .O(n15_adj_4394)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5285_17_lut (.I0(GND_net), .I1(n12509[14]), .I2(GND_net), 
            .I3(n31064), .O(n12255[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_4646));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5285_16_lut (.I0(GND_net), .I1(n12509[13]), .I2(n1117_adj_4311), 
            .I3(n31063), .O(n12255[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5389_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n13633[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5389_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5285_16 (.CI(n31063), .I0(n12509[13]), .I1(n1117_adj_4311), 
            .CO(n31064));
    SB_LUT4 add_5285_15_lut (.I0(GND_net), .I1(n12509[12]), .I2(n1044_adj_4310), 
            .I3(n31062), .O(n12255[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5285_15 (.CI(n31062), .I0(n12509[12]), .I1(n1044_adj_4310), 
            .CO(n31063));
    SB_LUT4 add_5285_14_lut (.I0(GND_net), .I1(n12509[11]), .I2(n971_adj_4309), 
            .I3(n31061), .O(n12255[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5389_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n30841));
    SB_LUT4 i19133_2_lut (.I0(n28[6]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[6]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19133_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_4645));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_4644));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_4643));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4677));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5285_14 (.CI(n31061), .I0(n12509[11]), .I1(n971_adj_4309), 
            .CO(n31062));
    SB_LUT4 add_5285_13_lut (.I0(GND_net), .I1(n12509[10]), .I2(n898_adj_4308), 
            .I3(n31060), .O(n12255[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5285_13 (.CI(n31060), .I0(n12509[10]), .I1(n898_adj_4308), 
            .CO(n31061));
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_4678));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_4679));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5285_12_lut (.I0(GND_net), .I1(n12509[9]), .I2(n825_adj_4306), 
            .I3(n31059), .O(n12255[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n30906), .I0(GND_net), .I1(n1[7]), 
            .CO(n30907));
    SB_CARRY add_5285_12 (.CI(n31059), .I0(n12509[9]), .I1(n825_adj_4306), 
            .CO(n31060));
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_4680));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_4681));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5285_11_lut (.I0(GND_net), .I1(n12509[8]), .I2(n752_adj_4305), 
            .I3(n31058), .O(n12255[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_4642));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5285_11 (.CI(n31058), .I0(n12509[8]), .I1(n752_adj_4305), 
            .CO(n31059));
    SB_LUT4 add_5285_10_lut (.I0(GND_net), .I1(n12509[7]), .I2(n679_adj_4297), 
            .I3(n31057), .O(n12255[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5285_10 (.CI(n31057), .I0(n12509[7]), .I1(n679_adj_4297), 
            .CO(n31058));
    SB_LUT4 add_5285_9_lut (.I0(GND_net), .I1(n12509[6]), .I2(n606), .I3(n31056), 
            .O(n12255[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_4682));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_4641));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588_adj_4640));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5285_9 (.CI(n31056), .I0(n12509[6]), .I1(n606), .CO(n31057));
    SB_LUT4 add_5285_8_lut (.I0(GND_net), .I1(n12509[5]), .I2(n533), .I3(n31055), 
            .O(n12255[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_4683));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661_adj_4639));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101_adj_4638));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5285_8 (.CI(n31055), .I0(n12509[5]), .I1(n533), .CO(n31056));
    SB_LUT4 add_5285_7_lut (.I0(GND_net), .I1(n12509[4]), .I2(n460_adj_4684), 
            .I3(n31054), .O(n12255[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(n28[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32_adj_4637));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_4636));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5285_7 (.CI(n31054), .I0(n12509[4]), .I1(n460_adj_4684), 
            .CO(n31055));
    SB_LUT4 add_5285_6_lut (.I0(GND_net), .I1(n12509[3]), .I2(n387_adj_4685), 
            .I3(n31053), .O(n12255[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807_adj_4634));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880_adj_4633));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953_adj_4632));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5285_6 (.CI(n31053), .I0(n12509[3]), .I1(n387_adj_4685), 
            .CO(n31054));
    SB_LUT4 add_5285_5_lut (.I0(GND_net), .I1(n12509[2]), .I2(n314_adj_4686), 
            .I3(n31052), .O(n12255[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5285_5 (.CI(n31052), .I0(n12509[2]), .I1(n314_adj_4686), 
            .CO(n31053));
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026_adj_4629));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099_adj_4628));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i24_3_lut (.I0(duty_23__N_3613[23]), .I1(n257[23]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(duty_23__N_3588[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i23_3_lut (.I0(duty_23__N_3613[22]), .I1(n257[22]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i23_3_lut (.I0(duty_23__N_3588[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5285_4_lut (.I0(GND_net), .I1(n12509[1]), .I2(n241_adj_4687), 
            .I3(n31051), .O(n12255[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5285_4 (.CI(n31051), .I0(n12509[1]), .I1(n241_adj_4687), 
            .CO(n31052));
    SB_LUT4 add_5285_3_lut (.I0(GND_net), .I1(n12509[0]), .I2(n168_adj_4688), 
            .I3(n31050), .O(n12255[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5285_3 (.CI(n31050), .I0(n12509[0]), .I1(n168_adj_4688), 
            .CO(n31051));
    SB_LUT4 add_5285_2_lut (.I0(GND_net), .I1(n26_adj_4689), .I2(n95_adj_4690), 
            .I3(GND_net), .O(n12255[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5285_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i22_3_lut (.I0(duty_23__N_3613[21]), .I1(n257[21]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5285_2 (.CI(GND_net), .I0(n26_adj_4689), .I1(n95_adj_4690), 
            .CO(n31050));
    SB_LUT4 add_5376_9_lut (.I0(GND_net), .I1(n13585[6]), .I2(n630_adj_4691), 
            .I3(n31049), .O(n13522[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5376_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5376_8_lut (.I0(GND_net), .I1(n13585[5]), .I2(n557_adj_4692), 
            .I3(n31048), .O(n13522[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5376_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5376_8 (.CI(n31048), .I0(n13585[5]), .I1(n557_adj_4692), 
            .CO(n31049));
    SB_LUT4 add_5376_7_lut (.I0(GND_net), .I1(n13585[4]), .I2(n484_adj_4693), 
            .I3(n31047), .O(n13522[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5376_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5376_7 (.CI(n31047), .I0(n13585[4]), .I1(n484_adj_4693), 
            .CO(n31048));
    SB_LUT4 add_5376_6_lut (.I0(GND_net), .I1(n13585[3]), .I2(n411_adj_4694), 
            .I3(n31046), .O(n13522[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5376_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5376_6 (.CI(n31046), .I0(n13585[3]), .I1(n411_adj_4694), 
            .CO(n31047));
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1[6]), .I3(n30905), .O(n13_adj_4395)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_LUT4 duty_23__I_0_i22_3_lut (.I0(duty_23__N_3588[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5376_5_lut (.I0(GND_net), .I1(n13585[2]), .I2(n338_adj_4696), 
            .I3(n31045), .O(n13522[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5376_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i21_3_lut (.I0(duty_23__N_3613[20]), .I1(n257[20]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5376_5 (.CI(n31045), .I0(n13585[2]), .I1(n338_adj_4696), 
            .CO(n31046));
    SB_LUT4 add_5376_4_lut (.I0(GND_net), .I1(n13585[1]), .I2(n265_adj_4697), 
            .I3(n31044), .O(n13522[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5376_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5376_4 (.CI(n31044), .I0(n13585[1]), .I1(n265_adj_4697), 
            .CO(n31045));
    SB_LUT4 add_5376_3_lut (.I0(GND_net), .I1(n13585[0]), .I2(n192_adj_4698), 
            .I3(n31043), .O(n13522[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5376_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5376_3 (.CI(n31043), .I0(n13585[0]), .I1(n192_adj_4698), 
            .CO(n31044));
    SB_LUT4 duty_23__I_0_i21_3_lut (.I0(duty_23__N_3588[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5376_2_lut (.I0(GND_net), .I1(n50_adj_4699), .I2(n119_adj_4700), 
            .I3(GND_net), .O(n13522[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5376_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5376_2 (.CI(GND_net), .I0(n50_adj_4699), .I1(n119_adj_4700), 
            .CO(n31043));
    SB_LUT4 mux_17_i20_3_lut (.I0(duty_23__N_3613[19]), .I1(n257[19]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_4701));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i20_3_lut (.I0(duty_23__N_3588[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_4702));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i19_3_lut (.I0(duty_23__N_3613[18]), .I1(n257[18]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n30905), .I0(GND_net), .I1(n1[6]), 
            .CO(n30906));
    SB_LUT4 add_5300_16_lut (.I0(GND_net), .I1(n12717[13]), .I2(n1120_adj_4702), 
            .I3(n31042), .O(n12509[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5300_15_lut (.I0(GND_net), .I1(n12717[12]), .I2(n1047_adj_4701), 
            .I3(n31041), .O(n12509[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5300_15 (.CI(n31041), .I0(n12717[12]), .I1(n1047_adj_4701), 
            .CO(n31042));
    SB_LUT4 duty_23__I_0_i19_3_lut (.I0(duty_23__N_3588[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i18_3_lut (.I0(duty_23__N_3613[17]), .I1(n257[17]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119_adj_4700));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5300_14_lut (.I0(GND_net), .I1(n12717[11]), .I2(n974_adj_4683), 
            .I3(n31040), .O(n12509[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(n28[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50_adj_4699));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5300_14 (.CI(n31040), .I0(n12717[11]), .I1(n974_adj_4683), 
            .CO(n31041));
    SB_LUT4 add_5300_13_lut (.I0(GND_net), .I1(n12717[10]), .I2(n901_adj_4682), 
            .I3(n31039), .O(n12509[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5300_13 (.CI(n31039), .I0(n12717[10]), .I1(n901_adj_4682), 
            .CO(n31040));
    SB_LUT4 add_5300_12_lut (.I0(GND_net), .I1(n12717[9]), .I2(n828_adj_4681), 
            .I3(n31038), .O(n12509[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5300_12 (.CI(n31038), .I0(n12717[9]), .I1(n828_adj_4681), 
            .CO(n31039));
    SB_LUT4 add_5300_11_lut (.I0(GND_net), .I1(n12717[8]), .I2(n755_adj_4680), 
            .I3(n31037), .O(n12509[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5300_11 (.CI(n31037), .I0(n12717[8]), .I1(n755_adj_4680), 
            .CO(n31038));
    SB_LUT4 add_5300_10_lut (.I0(GND_net), .I1(n12717[7]), .I2(n682_adj_4679), 
            .I3(n31036), .O(n12509[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5300_10 (.CI(n31036), .I0(n12717[7]), .I1(n682_adj_4679), 
            .CO(n31037));
    SB_LUT4 add_5300_9_lut (.I0(GND_net), .I1(n12717[6]), .I2(n609_adj_4678), 
            .I3(n31035), .O(n12509[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5300_9 (.CI(n31035), .I0(n12717[6]), .I1(n609_adj_4678), 
            .CO(n31036));
    SB_LUT4 add_5300_8_lut (.I0(GND_net), .I1(n12717[5]), .I2(n536_adj_4677), 
            .I3(n31034), .O(n12509[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192_adj_4698));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5300_8 (.CI(n31034), .I0(n12717[5]), .I1(n536_adj_4677), 
            .CO(n31035));
    SB_LUT4 add_5300_7_lut (.I0(GND_net), .I1(n12717[4]), .I2(n463), .I3(n31033), 
            .O(n12509[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5300_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i18_3_lut (.I0(duty_23__N_3588[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i17_3_lut (.I0(duty_23__N_3613[16]), .I1(n257[16]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i17_3_lut (.I0(duty_23__N_3588[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265_adj_4697));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i16_3_lut (.I0(duty_23__N_3613[15]), .I1(n257[15]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i16_3_lut (.I0(duty_23__N_3588[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i15_3_lut (.I0(duty_23__N_3613[14]), .I1(n257[14]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i15_3_lut (.I0(duty_23__N_3588[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i14_3_lut (.I0(duty_23__N_3613[13]), .I1(n257[13]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i14_3_lut (.I0(duty_23__N_3588[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i13_3_lut (.I0(duty_23__N_3613[12]), .I1(n257[12]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338_adj_4696));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i13_3_lut (.I0(duty_23__N_3588[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i12_3_lut (.I0(duty_23__N_3613[11]), .I1(n257[11]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i12_3_lut (.I0(duty_23__N_3588[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411_adj_4694));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i11_3_lut (.I0(duty_23__N_3613[10]), .I1(n257[10]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i11_3_lut (.I0(duty_23__N_3588[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484_adj_4693));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i10_3_lut (.I0(duty_23__N_3613[9]), .I1(n257[9]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i10_3_lut (.I0(duty_23__N_3588[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557_adj_4692));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i9_3_lut (.I0(duty_23__N_3613[8]), .I1(n257[8]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i9_3_lut (.I0(duty_23__N_3588[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i8_3_lut (.I0(duty_23__N_3613[7]), .I1(n257[7]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i8_3_lut (.I0(duty_23__N_3588[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i7_3_lut (.I0(duty_23__N_3613[6]), .I1(n257[6]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i7_3_lut (.I0(duty_23__N_3588[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i6_3_lut (.I0(duty_23__N_3613[5]), .I1(n257[5]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i6_3_lut (.I0(duty_23__N_3588[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i5_3_lut (.I0(duty_23__N_3613[4]), .I1(n257[4]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i5_3_lut (.I0(duty_23__N_3588[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i4_3_lut (.I0(duty_23__N_3613[3]), .I1(n257[3]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(n28[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630_adj_4691));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i4_3_lut (.I0(duty_23__N_3588[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_4690));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_4627));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(n28[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4689));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4626));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22112_3_lut_4_lut (.I0(\Kp[3] ), .I1(n28[18]), .I2(n4_adj_4703), 
            .I3(n13692[1]), .O(n6_adj_4420));   // verilog/motorControl.v(34[16:22])
    defparam i22112_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_4625));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_4624));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168_adj_4688));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1520 (.I0(\Kp[3] ), .I1(n28[18]), .I2(n13692[1]), 
            .I3(n4_adj_4703), .O(n13668[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1520.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_1521 (.I0(\Kp[2] ), .I1(n28[18]), .I2(n13692[0]), 
            .I3(n30468), .O(n13668[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1521.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4687));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_4623));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_4622));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_4621));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22104_3_lut_4_lut (.I0(\Kp[2] ), .I1(n28[18]), .I2(n30468), 
            .I3(n13692[0]), .O(n4_adj_4703));   // verilog/motorControl.v(34[16:22])
    defparam i22104_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_4620));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22091_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[19]), .I2(n28[18]), 
            .I3(\Kp[1] ), .O(n13668[0]));   // verilog/motorControl.v(34[16:22])
    defparam i22091_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585_adj_4619));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658_adj_4618));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19134_2_lut (.I0(n28[7]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[7]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22093_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[19]), .I2(n28[18]), 
            .I3(\Kp[1] ), .O(n30468));   // verilog/motorControl.v(34[16:22])
    defparam i22093_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950_adj_4617));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023_adj_4616));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096_adj_4615));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174_adj_4614));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_4613));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4612));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22055_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[20]), .I2(n28[19]), 
            .I3(\Kp[1] ), .O(n30427));   // verilog/motorControl.v(34[16:22])
    defparam i22055_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i22053_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[20]), .I2(n28[19]), 
            .I3(\Kp[1] ), .O(n13692[0]));   // verilog/motorControl.v(34[16:22])
    defparam i22053_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i19135_2_lut (.I0(n28[8]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[8]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19135_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_4611));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_4610));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247_adj_4609));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_4608));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_4607));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_4606));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_4605));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591_adj_4604));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664_adj_4603));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_4602));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1522 (.I0(\Kp[2] ), .I1(n28[19]), .I2(n13707[0]), 
            .I3(n30427), .O(n13692[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1522.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810_adj_4601));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883_adj_4600));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956_adj_4599));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22066_3_lut_4_lut (.I0(\Kp[2] ), .I1(n28[19]), .I2(n30427), 
            .I3(n13707[0]), .O(n4_adj_4428));   // verilog/motorControl.v(34[16:22])
    defparam i22066_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i22017_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[21]), .I2(n28[20]), 
            .I3(\Kp[1] ), .O(n30386));   // verilog/motorControl.v(34[16:22])
    defparam i22017_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i22015_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n28[21]), .I2(n28[20]), 
            .I3(\Kp[1] ), .O(n13707[0]));   // verilog/motorControl.v(34[16:22])
    defparam i22015_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_4598));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102_adj_4597));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83_adj_4596));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4595));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_4594));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_4593));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_4592));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320_adj_4591));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_4589));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22028_3_lut_4_lut (.I0(\Kp[2] ), .I1(n28[20]), .I2(n30386), 
            .I3(n13712[0]), .O(n4_adj_4439));   // verilog/motorControl.v(34[16:22])
    defparam i22028_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314_adj_4686));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1523 (.I0(\Kp[2] ), .I1(n28[20]), .I2(n13712[0]), 
            .I3(n30386), .O(n13707[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1523.LUT_INIT = 16'h8778;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_4587));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_4586));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594_adj_4585));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_17_i3_3_lut (.I0(duty_23__N_3613[2]), .I1(n257[2]), .I2(n256), 
            .I3(GND_net), .O(duty_23__N_3588[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i3_3_lut (.I0(duty_23__N_3588[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3612), .I3(GND_net), .O(duty_23__N_3489[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667_adj_4584));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_4583));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813_adj_4582));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_4581));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_4580));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_4579));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_4578));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_4577));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4576));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_4575));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_4574));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_4573));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[0]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19136_2_lut (.I0(n28[9]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[9]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19136_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[1]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393_adj_4569));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466_adj_4568));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[2]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19137_2_lut (.I0(n28[10]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[10]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19137_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4413));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387_adj_4685));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4565));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[3]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_4563));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19138_2_lut (.I0(n28[11]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[11]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22158_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [18]), 
            .I2(n4), .I3(n9993[1]), .O(n6_adj_4371));   // verilog/motorControl.v(34[25:36])
    defparam i22158_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_4562));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1524 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [18]), 
            .I2(n9993[1]), .I3(n4), .O(n9986[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1524.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_1525 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [19]), 
            .I2(n9999[0]), .I3(n30561), .O(n9993[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1525.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597_adj_4561));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22189_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [19]), 
            .I2(n30561), .I3(n9999[0]), .O(n4_adj_4375));   // verilog/motorControl.v(34[25:36])
    defparam i22189_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670_adj_4560));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[4]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743_adj_4558));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816_adj_4557));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889_adj_4556));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962_adj_4555));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035_adj_4554));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22176_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [20]), 
            .I2(\PID_CONTROLLER.integral_23__N_3513 [19]), .I3(\Ki[1] ), 
            .O(n9993[0]));   // verilog/motorControl.v(34[25:36])
    defparam i22176_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108_adj_4553));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22178_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [20]), 
            .I2(\PID_CONTROLLER.integral_23__N_3513 [19]), .I3(\Ki[1] ), 
            .O(n30561));   // verilog/motorControl.v(34[25:36])
    defparam i22178_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_4552));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4551));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4550));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4549));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4548));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_4546));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19139_2_lut (.I0(n28[12]), .I1(\PID_CONTROLLER.integral_23__N_3561 ), 
            .I2(GND_net), .I3(GND_net), .O(n3141[12]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i19139_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_4545));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_4544));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600_adj_4543));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673_adj_4542));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746_adj_4541));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819_adj_4540));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892_adj_4539));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539_adj_4538));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965_adj_4537));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038_adj_4536));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111_adj_4535));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_4534));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4533));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_4532));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_4531));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_4530));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_4529));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_4528));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_4527));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603_adj_4526));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676_adj_4525));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22220_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [20]), 
            .I2(n30595), .I3(n10004[0]), .O(n4_adj_4383));   // verilog/motorControl.v(34[25:36])
    defparam i22220_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_4524));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(n28[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4704[5]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut_adj_1526 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [20]), 
            .I2(n10004[0]), .I3(n30595), .O(n9999[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1526.LUT_INIT = 16'h8778;
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822_adj_4522));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895_adj_4521));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968_adj_4520));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(n28[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612_adj_4519));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041_adj_4518));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114_adj_4517));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4516));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(n28[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460_adj_4684));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22207_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3513 [20]), .I3(\Ki[1] ), 
            .O(n9999[0]));   // verilog/motorControl.v(34[25:36])
    defparam i22207_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_4515));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22209_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3513 [20]), .I3(\Ki[1] ), 
            .O(n30595));   // verilog/motorControl.v(34[25:36])
    defparam i22209_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3513 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_4514));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=51, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=37 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (GND_net, CLK_c, n3460, \state[1] , \state[1]_adj_12 , 
            \state[2] , n7, read, \state[0] , n15, \state[3] , n6, 
            n35272, n36440, n35591, n27098, n35254, VCC_net, n22318, 
            rw, n35362, data_ready, n4760, \saved_addr[0] , \state[0]_adj_13 , 
            n3957, n27086, n4, n4_adj_14, n10, n10_adj_15, \state_7__N_3881[3] , 
            n10_adj_16, scl_enable_N_3958, scl_enable, sda_enable, \state_7__N_3865[0] , 
            n5180, n15_adj_17, n8, n987, n20731, n20726, n39285, 
            n22330, \data[0] , n22321, n22300, \data[1] , n22299, 
            \data[2] , n22298, \data[3] , n22297, \data[4] , n22296, 
            \data[5] , n22295, \data[6] , n22294, \data[7] ) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    output [0:0]n3460;
    output \state[1] ;
    output \state[1]_adj_12 ;
    output \state[2] ;
    output n7;
    input read;
    output \state[0] ;
    input n15;
    output \state[3] ;
    output n6;
    input n35272;
    input n36440;
    output n35591;
    output n27098;
    input n35254;
    input VCC_net;
    input n22318;
    output rw;
    input n35362;
    output data_ready;
    output n4760;
    output \saved_addr[0] ;
    output \state[0]_adj_13 ;
    input n3957;
    output n27086;
    output n4;
    output n4_adj_14;
    output n10;
    input n10_adj_15;
    output \state_7__N_3881[3] ;
    output n10_adj_16;
    input scl_enable_N_3958;
    output scl_enable;
    output sda_enable;
    output \state_7__N_3865[0] ;
    input n5180;
    output n15_adj_17;
    input n8;
    output [0:0]n987;
    output n20731;
    output n20726;
    output n39285;
    input n22330;
    output \data[0] ;
    input n22321;
    input n22300;
    output \data[1] ;
    input n22299;
    output \data[2] ;
    input n22298;
    output \data[3] ;
    input n22297;
    output \data[4] ;
    input n22296;
    output \data[5] ;
    input n22295;
    output \data[6] ;
    input n22294;
    output \data[7] ;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [15:0]delay_counter_15__N_3767;
    wire [15:0]delay_counter;   // verilog/eeprom.v(23[12:25])
    wire [15:0]n3177;
    
    wire n30783, n30784, n22002, n22163, n30782, n30781, enable, 
        n30780, n30779, n20600, n28, n26, n27, n25, n30793, 
        n30792, n30791, n30790, n30789, n30788, n30787, n30786, 
        n30785;
    
    SB_LUT4 add_727_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n3177[14]), 
            .I3(n30783), .O(delay_counter_15__N_3767[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_727_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_727_7 (.CI(n30783), .I0(delay_counter[5]), .I1(n3177[14]), 
            .CO(n30784));
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n22002), 
            .D(delay_counter_15__N_3767[15]), .R(n22163));   // verilog/eeprom.v(25[8] 57[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n22002), 
            .D(delay_counter_15__N_3767[14]), .R(n22163));   // verilog/eeprom.v(25[8] 57[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n22002), 
            .D(delay_counter_15__N_3767[13]), .R(n22163));   // verilog/eeprom.v(25[8] 57[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n22002), 
            .D(delay_counter_15__N_3767[12]), .R(n22163));   // verilog/eeprom.v(25[8] 57[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n22002), 
            .D(delay_counter_15__N_3767[11]), .R(n22163));   // verilog/eeprom.v(25[8] 57[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n22002), 
            .D(delay_counter_15__N_3767[10]), .S(n22163));   // verilog/eeprom.v(25[8] 57[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n22002), 
            .D(delay_counter_15__N_3767[9]), .S(n22163));   // verilog/eeprom.v(25[8] 57[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n22002), 
            .D(delay_counter_15__N_3767[8]), .S(n22163));   // verilog/eeprom.v(25[8] 57[4])
    SB_LUT4 add_727_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(n3177[14]), 
            .I3(n30782), .O(delay_counter_15__N_3767[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_727_6_lut.LUT_INIT = 16'hC33C;
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n22002), 
            .D(delay_counter_15__N_3767[7]), .S(n22163));   // verilog/eeprom.v(25[8] 57[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n22002), 
            .D(delay_counter_15__N_3767[6]), .S(n22163));   // verilog/eeprom.v(25[8] 57[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n22002), 
            .D(delay_counter_15__N_3767[5]), .R(n22163));   // verilog/eeprom.v(25[8] 57[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n22002), 
            .D(delay_counter_15__N_3767[4]), .S(n22163));   // verilog/eeprom.v(25[8] 57[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n22002), 
            .D(delay_counter_15__N_3767[3]), .R(n22163));   // verilog/eeprom.v(25[8] 57[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n22002), 
            .D(delay_counter_15__N_3767[2]), .R(n22163));   // verilog/eeprom.v(25[8] 57[4])
    SB_CARRY add_727_6 (.CI(n30782), .I0(delay_counter[4]), .I1(n3177[14]), 
            .CO(n30783));
    SB_LUT4 add_727_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n3177[14]), 
            .I3(n30781), .O(delay_counter_15__N_3767[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_727_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR enable_39 (.Q(enable), .C(CLK_c), .D(n3460[0]), .R(\state[1] ));   // verilog/eeprom.v(25[8] 57[4])
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n22002), 
            .D(delay_counter_15__N_3767[1]), .R(n22163));   // verilog/eeprom.v(25[8] 57[4])
    SB_CARRY add_727_5 (.CI(n30781), .I0(delay_counter[3]), .I1(n3177[14]), 
            .CO(n30782));
    SB_LUT4 add_727_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n3177[14]), 
            .I3(n30780), .O(delay_counter_15__N_3767[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_727_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_727_4 (.CI(n30780), .I0(delay_counter[2]), .I1(n3177[14]), 
            .CO(n30781));
    SB_LUT4 add_727_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n3177[14]), 
            .I3(n30779), .O(delay_counter_15__N_3767[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_727_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_727_3 (.CI(n30779), .I0(delay_counter[1]), .I1(n3177[14]), 
            .CO(n30780));
    SB_LUT4 add_727_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n3177[14]), 
            .I3(GND_net), .O(delay_counter_15__N_3767[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_727_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_727_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n3177[14]), 
            .CO(n30779));
    SB_LUT4 i2_2_lut (.I0(\state[1]_adj_12 ), .I1(\state[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n7));   // verilog/eeprom.v(41[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mux_902_Mux_0_i1_4_lut (.I0(read), .I1(n20600), .I2(\state[0] ), 
            .I3(n15), .O(n3460[0]));   // verilog/eeprom.v(28[3] 56[10])
    defparam mux_902_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_LUT4 i13773_2_lut (.I0(n22002), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n22163));   // verilog/eeprom.v(25[8] 57[4])
    defparam i13773_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut (.I0(read), .I1(\state[1] ), .I2(\state[0] ), .I3(GND_net), 
            .O(n22002));
    defparam i1_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 i2_2_lut_adj_1510 (.I0(\state[3] ), .I1(n20600), .I2(GND_net), 
            .I3(GND_net), .O(n6));   // verilog/eeprom.v(41[12:28])
    defparam i2_2_lut_adj_1510.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut (.I0(delay_counter[6]), .I1(delay_counter[10]), .I2(delay_counter[12]), 
            .I3(delay_counter[8]), .O(n28));   // verilog/eeprom.v(41[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[11]), .I1(delay_counter[2]), .I2(delay_counter[7]), 
            .I3(delay_counter[5]), .O(n26));   // verilog/eeprom.v(41[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n22002), 
            .D(delay_counter_15__N_3767[0]), .R(n22163));   // verilog/eeprom.v(25[8] 57[4])
    SB_DFF state__i1 (.Q(\state[1] ), .C(CLK_c), .D(n35272));   // verilog/eeprom.v(25[8] 57[4])
    SB_LUT4 i1_4_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(n36440), 
            .I3(n15), .O(n35591));   // verilog/eeprom.v(50[5:9])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hfcf8;
    SB_LUT4 i19403_2_lut_3_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(n15), 
            .I3(GND_net), .O(n27098));   // verilog/eeprom.v(50[5:9])
    defparam i19403_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_DFFE state__i0 (.Q(\state[0] ), .C(CLK_c), .E(VCC_net), .D(n35254));   // verilog/eeprom.v(25[8] 57[4])
    SB_LUT4 i11_4_lut (.I0(delay_counter[15]), .I1(delay_counter[3]), .I2(delay_counter[14]), 
            .I3(delay_counter[1]), .O(n27));   // verilog/eeprom.v(41[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[9]), .I2(delay_counter[13]), 
            .I3(delay_counter[0]), .O(n25));   // verilog/eeprom.v(41[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n20600));   // verilog/eeprom.v(41[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i30125_2_lut (.I0(n20600), .I1(n15), .I2(GND_net), .I3(GND_net), 
            .O(n3177[14]));   // verilog/eeprom.v(45[18] 47[12])
    defparam i30125_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 add_727_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n3177[14]), 
            .I3(n30793), .O(delay_counter_15__N_3767[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_727_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_727_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n3177[14]), 
            .I3(n30792), .O(delay_counter_15__N_3767[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_727_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_727_16 (.CI(n30792), .I0(delay_counter[14]), .I1(n3177[14]), 
            .CO(n30793));
    SB_LUT4 add_727_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n3177[14]), 
            .I3(n30791), .O(delay_counter_15__N_3767[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_727_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_727_15 (.CI(n30791), .I0(delay_counter[13]), .I1(n3177[14]), 
            .CO(n30792));
    SB_LUT4 add_727_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n3177[14]), 
            .I3(n30790), .O(delay_counter_15__N_3767[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_727_14_lut.LUT_INIT = 16'hC33C;
    SB_DFF rw_43 (.Q(rw), .C(CLK_c), .D(n22318));   // verilog/eeprom.v(25[8] 57[4])
    SB_DFF data_ready_42 (.Q(data_ready), .C(CLK_c), .D(n35362));   // verilog/eeprom.v(25[8] 57[4])
    SB_CARRY add_727_14 (.CI(n30790), .I0(delay_counter[12]), .I1(n3177[14]), 
            .CO(n30791));
    SB_LUT4 add_727_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n3177[14]), 
            .I3(n30789), .O(delay_counter_15__N_3767[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_727_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_727_13 (.CI(n30789), .I0(delay_counter[11]), .I1(n3177[14]), 
            .CO(n30790));
    SB_LUT4 add_727_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(n3177[14]), 
            .I3(n30788), .O(delay_counter_15__N_3767[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_727_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_727_12 (.CI(n30788), .I0(delay_counter[10]), .I1(n3177[14]), 
            .CO(n30789));
    SB_LUT4 add_727_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(n3177[14]), 
            .I3(n30787), .O(delay_counter_15__N_3767[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_727_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_727_11 (.CI(n30787), .I0(delay_counter[9]), .I1(n3177[14]), 
            .CO(n30788));
    SB_LUT4 add_727_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(n3177[14]), 
            .I3(n30786), .O(delay_counter_15__N_3767[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_727_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_727_10 (.CI(n30786), .I0(delay_counter[8]), .I1(n3177[14]), 
            .CO(n30787));
    SB_LUT4 add_727_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(n3177[14]), 
            .I3(n30785), .O(delay_counter_15__N_3767[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_727_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_727_9 (.CI(n30785), .I0(delay_counter[7]), .I1(n3177[14]), 
            .CO(n30786));
    SB_LUT4 add_727_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(n3177[14]), 
            .I3(n30784), .O(delay_counter_15__N_3767[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_727_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_727_8 (.CI(n30784), .I0(delay_counter[6]), .I1(n3177[14]), 
            .CO(n30785));
    i2c_controller i2c (.n4760(n4760), .\state[3] (\state[3] ), .\state[2] (\state[2] ), 
            .\state[1] (\state[1]_adj_12 ), .\saved_addr[0] (\saved_addr[0] ), 
            .GND_net(GND_net), .\state[0] (\state[0]_adj_13 ), .n3957(n3957), 
            .n27086(n27086), .n4(n4), .n4_adj_8(n4_adj_14), .n10(n10), 
            .n10_adj_9(n10_adj_15), .\state_7__N_3881[3] (\state_7__N_3881[3] ), 
            .enable(enable), .n10_adj_10(n10_adj_16), .CLK_c(CLK_c), .scl_enable_N_3958(scl_enable_N_3958), 
            .scl_enable(scl_enable), .sda_enable(sda_enable), .\state_7__N_3865[0] (\state_7__N_3865[0] ), 
            .n5180(n5180), .n15(n15_adj_17), .n8(n8), .VCC_net(VCC_net), 
            .n987({n987}), .n20731(n20731), .n20726(n20726), .n15_adj_11(n15), 
            .n39285(n39285), .n22330(n22330), .\data[0] (\data[0] ), .n22321(n22321), 
            .n22300(n22300), .\data[1] (\data[1] ), .n22299(n22299), .\data[2] (\data[2] ), 
            .n22298(n22298), .\data[3] (\data[3] ), .n22297(n22297), .\data[4] (\data[4] ), 
            .n22296(n22296), .\data[5] (\data[5] ), .n22295(n22295), .\data[6] (\data[6] ), 
            .n22294(n22294), .\data[7] (\data[7] )) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(59[16] 72[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (n4760, \state[3] , \state[2] , \state[1] , \saved_addr[0] , 
            GND_net, \state[0] , n3957, n27086, n4, n4_adj_8, n10, 
            n10_adj_9, \state_7__N_3881[3] , enable, n10_adj_10, CLK_c, 
            scl_enable_N_3958, scl_enable, sda_enable, \state_7__N_3865[0] , 
            n5180, n15, n8, VCC_net, n987, n20731, n20726, n15_adj_11, 
            n39285, n22330, \data[0] , n22321, n22300, \data[1] , 
            n22299, \data[2] , n22298, \data[3] , n22297, \data[4] , 
            n22296, \data[5] , n22295, \data[6] , n22294, \data[7] ) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    output n4760;
    output \state[3] ;
    output \state[2] ;
    output \state[1] ;
    output \saved_addr[0] ;
    input GND_net;
    output \state[0] ;
    input n3957;
    output n27086;
    output n4;
    output n4_adj_8;
    output n10;
    input n10_adj_9;
    output \state_7__N_3881[3] ;
    input enable;
    output n10_adj_10;
    input CLK_c;
    input scl_enable_N_3958;
    output scl_enable;
    output sda_enable;
    output \state_7__N_3865[0] ;
    input n5180;
    output n15;
    input n8;
    input VCC_net;
    output [0:0]n987;
    output n20731;
    output n20726;
    input n15_adj_11;
    output n39285;
    input n22330;
    output \data[0] ;
    input n22321;
    input n22300;
    output \data[1] ;
    input n22299;
    output \data[2] ;
    input n22298;
    output \data[3] ;
    input n22297;
    output \data[4] ;
    input n22296;
    output \data[5] ;
    input n22295;
    output \data[6] ;
    input n22294;
    output \data[7] ;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(40[6:13])
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [7:0]n988;
    
    wire n22043;
    wire [7:0]counter;   // verilog/i2c_controller.v(35[12:19])
    
    wire n22208, n35408, n37171, n27237, n27550, n5, n27852, n39269, 
        n39205;
    wire [0:0]n3958;
    
    wire counter2_7__N_3852, n14136, n4_c, n33, n37, n22154, n34, 
        n5057, n13981;
    wire [7:0]counter2;   // verilog/i2c_controller.v(36[12:20])
    
    wire n6, i2c_clk_N_3957, n21849, n4753, n11, n27154, n39290, 
        n7, n21937, n22149, sda_out, n12, n36448;
    wire [4:0]n25;
    
    wire n11_adj_4271, n11_adj_4272, n9, n11_adj_4273, n31104, n31103, 
        n31102, n31101, n31100, n31099, n31098, n31698, n31697, 
        n31696, n31695;
    
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n22043), .D(n988[7]), 
            .R(n22208));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n22043), .D(n988[6]), 
            .R(n22208));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n22043), .D(n988[5]), 
            .R(n22208));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n22043), .D(n988[4]), 
            .R(n22208));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n22043), .D(n988[3]), 
            .R(n22208));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n22043), .D(n988[2]), 
            .S(n22208));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n22043), .D(n988[1]), 
            .S(n22208));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n4760), .D(n35408), 
            .S(n37171));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n4760), .D(n27237), 
            .S(n27550));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n4760), .D(n5), 
            .S(n27852));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_LUT4 i29540_2_lut (.I0(counter[1]), .I1(\saved_addr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n39269));   // verilog/i2c_controller.v(180[28:35])
    defparam i29540_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i29531_4_lut (.I0(n39269), .I1(\state[1] ), .I2(counter[0]), 
            .I3(counter[2]), .O(n39205));   // verilog/i2c_controller.v(163[4] 196[11])
    defparam i29531_4_lut.LUT_INIT = 16'hc008;
    SB_LUT4 mux_1055_i1_4_lut (.I0(n39205), .I1(\state[0] ), .I2(n3957), 
            .I3(\state[2] ), .O(n3958[0]));   // verilog/i2c_controller.v(163[4] 196[11])
    defparam mux_1055_i1_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 i30150_2_lut (.I0(i2c_clk), .I1(counter2_7__N_3852), .I2(GND_net), 
            .I3(GND_net), .O(n14136));   // verilog/i2c_controller.v(68[8:33])
    defparam i30150_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i18695_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n27086));
    defparam i18695_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut (.I0(\state[2] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n4_c));   // verilog/i2c_controller.v(163[4] 196[11])
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_3_lut (.I0(\state[1] ), .I1(n33), .I2(n37), .I3(GND_net), 
            .O(n22154));
    defparam i1_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i30152_4_lut (.I0(n3957), .I1(n34), .I2(n4_c), .I3(n37), 
            .O(n5057));
    defparam i30152_4_lut.LUT_INIT = 16'haf8c;
    SB_LUT4 i30182_2_lut (.I0(\state[0] ), .I1(n3957), .I2(GND_net), .I3(GND_net), 
            .O(n13981));   // verilog/i2c_controller.v(163[4] 196[11])
    defparam i30182_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 equal_148_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(138[6:23])
    defparam equal_148_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_150_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_8));   // verilog/i2c_controller.v(138[6:23])
    defparam equal_150_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_1503 (.I0(counter2[0]), .I1(counter2[4]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i1_2_lut_adj_1503.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[2]), .I2(counter2[1]), 
            .I3(n6), .O(counter2_7__N_3852));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_1504 (.I0(i2c_clk), .I1(counter2_7__N_3852), .I2(GND_net), 
            .I3(GND_net), .O(i2c_clk_N_3957));
    defparam i1_2_lut_adj_1504.LUT_INIT = 16'h6666;
    SB_LUT4 state_7__I_0_144_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(137[5:14])
    defparam state_7__I_0_144_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i30102_4_lut (.I0(n21849), .I1(n4753), .I2(n11), .I3(n27154), 
            .O(n4760));
    defparam i30102_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i29498_4_lut (.I0(n10_adj_9), .I1(n10), .I2(\state_7__N_3881[3] ), 
            .I3(enable), .O(n39290));   // verilog/i2c_controller.v(90[4] 154[11])
    defparam i29498_4_lut.LUT_INIT = 16'h7073;
    SB_LUT4 i1_4_lut (.I0(\state[1] ), .I1(n7), .I2(n39290), .I3(\state[0] ), 
            .O(n35408));   // verilog/i2c_controller.v(90[4] 154[11])
    defparam i1_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_10));   // verilog/i2c_controller.v(107[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_DFF i2c_clk_122 (.Q(i2c_clk), .C(CLK_c), .D(i2c_clk_N_3957));   // verilog/i2c_controller.v(57[9] 69[5])
    SB_DFFN i2c_scl_enable_124 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_3958));   // verilog/i2c_controller.v(74[12] 80[6])
    SB_DFFNESS write_enable_132 (.Q(sda_enable), .C(i2c_clk), .E(n5057), 
            .D(n13981), .S(n22154));   // verilog/i2c_controller.v(162[12] 197[6])
    SB_DFFESS enable_slow_121 (.Q(\state_7__N_3865[0] ), .C(CLK_c), .E(n21937), 
            .D(n14136), .S(enable));   // verilog/i2c_controller.v(57[9] 69[5])
    SB_DFFNE sda_out_133 (.Q(sda_out), .C(i2c_clk), .E(n22149), .D(n3958[0]));   // verilog/i2c_controller.v(162[12] 197[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n22043), .D(n988[0]), 
            .S(n22208));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(107[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10_adj_10), 
            .O(n4753));   // verilog/i2c_controller.v(107[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n4753), .I1(n36448), .I2(n5180), .I3(n37), 
            .O(n22043));
    defparam i17_4_lut.LUT_INIT = 16'h3a30;
    SB_DFFSR counter2_1516_1517__i1 (.Q(counter2[0]), .C(CLK_c), .D(n25[0]), 
            .R(counter2_7__N_3852));   // verilog/i2c_controller.v(68[20:32])
    SB_LUT4 i1_4_lut_adj_1505 (.I0(n11_adj_4271), .I1(n11_adj_4272), .I2(\state_7__N_3881[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(90[4] 154[11])
    defparam i1_4_lut_adj_1505.LUT_INIT = 16'h5755;
    SB_LUT4 i18762_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n27154));
    defparam i18762_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_adj_1506 (.I0(\state[3] ), .I1(\state[2] ), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i1_2_lut_adj_1506.LUT_INIT = 16'h2222;
    SB_LUT4 state_7__I_0_144_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(137[5:14])
    defparam state_7__I_0_144_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 state_7__I_0_140_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4272));
    defparam state_7__I_0_140_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 equal_92_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n15));   // verilog/i2c_controller.v(75[27:43])
    defparam equal_92_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 state_7__I_0_145_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4271));   // verilog/i2c_controller.v(75[27:43])
    defparam state_7__I_0_145_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i30258_2_lut_3_lut (.I0(sda_out), .I1(sda_enable), .I2(n11_adj_4272), 
            .I3(GND_net), .O(n27237));
    defparam i30258_2_lut_3_lut.LUT_INIT = 16'h0707;
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_LUT4 i18690_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(n987[0]));   // verilog/i2c_controller.v(44[19:55])
    defparam i18690_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1765_2_lut (.I0(sda_out), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(\state_7__N_3881[3] ));   // verilog/i2c_controller.v(45[9:16])
    defparam i1765_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut (.I0(n9), .I1(n10), .I2(counter[0]), .I3(GND_net), 
            .O(n20731));   // verilog/i2c_controller.v(137[5:14])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_1507 (.I0(n9), .I1(n10), .I2(counter[0]), 
            .I3(GND_net), .O(n20726));   // verilog/i2c_controller.v(137[5:14])
    defparam i1_2_lut_3_lut_adj_1507.LUT_INIT = 16'hfefe;
    SB_LUT4 i30301_3_lut_4_lut (.I0(n9), .I1(n10), .I2(n11_adj_4273), 
            .I3(n4760), .O(n27550));   // verilog/i2c_controller.v(137[5:14])
    defparam i30301_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_LUT4 sub_95_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n31104), .O(n988[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_95_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29501_3_lut_4_lut (.I0(n11), .I1(n11_adj_4273), .I2(n15_adj_11), 
            .I3(\state_7__N_3865[0] ), .O(n39285));
    defparam i29501_3_lut_4_lut.LUT_INIT = 16'h8088;
    SB_LUT4 sub_95_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n31103), .O(n988[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_95_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i30299_3_lut_4_lut (.I0(n11), .I1(n11_adj_4273), .I2(n15), 
            .I3(n4760), .O(n27852));
    defparam i30299_3_lut_4_lut.LUT_INIT = 16'h7f00;
    SB_CARRY sub_95_add_2_8 (.CI(n31103), .I0(counter[6]), .I1(VCC_net), 
            .CO(n31104));
    SB_LUT4 sub_95_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n31102), .O(n988[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_95_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_95_add_2_7 (.CI(n31102), .I0(counter[5]), .I1(VCC_net), 
            .CO(n31103));
    SB_LUT4 sub_95_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n31101), .O(n988[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_95_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_95_add_2_6 (.CI(n31101), .I0(counter[4]), .I1(VCC_net), 
            .CO(n31102));
    SB_LUT4 sub_95_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n31100), .O(n988[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_95_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_95_add_2_5 (.CI(n31100), .I0(counter[3]), .I1(VCC_net), 
            .CO(n31101));
    SB_LUT4 sub_95_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n31099), .O(n988[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_95_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_95_add_2_4 (.CI(n31099), .I0(counter[2]), .I1(VCC_net), 
            .CO(n31100));
    SB_LUT4 sub_95_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n31098), .O(n988[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_95_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_95_add_2_3 (.CI(n31098), .I0(counter[1]), .I1(VCC_net), 
            .CO(n31099));
    SB_LUT4 sub_95_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n988[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_95_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_95_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n31098));
    SB_DFF data_out__i1 (.Q(\data[0] ), .C(i2c_clk), .D(n22330));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n22321));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFF data_out__i2 (.Q(\data[1] ), .C(i2c_clk), .D(n22300));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFF data_out__i3 (.Q(\data[2] ), .C(i2c_clk), .D(n22299));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFF data_out__i4 (.Q(\data[3] ), .C(i2c_clk), .D(n22298));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFF data_out__i5 (.Q(\data[4] ), .C(i2c_clk), .D(n22297));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFF data_out__i6 (.Q(\data[5] ), .C(i2c_clk), .D(n22296));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFF data_out__i7 (.Q(\data[6] ), .C(i2c_clk), .D(n22295));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFF data_out__i8 (.Q(\data[7] ), .C(i2c_clk), .D(n22294));   // verilog/i2c_controller.v(89[8] 155[6])
    SB_DFFSR counter2_1516_1517__i2 (.Q(counter2[1]), .C(CLK_c), .D(n25[1]), 
            .R(counter2_7__N_3852));   // verilog/i2c_controller.v(68[20:32])
    SB_DFFSR counter2_1516_1517__i3 (.Q(counter2[2]), .C(CLK_c), .D(n25[2]), 
            .R(counter2_7__N_3852));   // verilog/i2c_controller.v(68[20:32])
    SB_DFFSR counter2_1516_1517__i4 (.Q(counter2[3]), .C(CLK_c), .D(n25[3]), 
            .R(counter2_7__N_3852));   // verilog/i2c_controller.v(68[20:32])
    SB_DFFSR counter2_1516_1517__i5 (.Q(counter2[4]), .C(CLK_c), .D(n25[4]), 
            .R(counter2_7__N_3852));   // verilog/i2c_controller.v(68[20:32])
    SB_LUT4 counter2_1516_1517_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n31698), .O(n25[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1516_1517_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_1516_1517_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n31697), .O(n25[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1516_1517_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1516_1517_add_4_5 (.CI(n31697), .I0(GND_net), .I1(counter2[3]), 
            .CO(n31698));
    SB_LUT4 counter2_1516_1517_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n31696), .O(n25[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1516_1517_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1516_1517_add_4_4 (.CI(n31696), .I0(GND_net), .I1(counter2[2]), 
            .CO(n31697));
    SB_LUT4 counter2_1516_1517_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n31695), .O(n25[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1516_1517_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i26387_2_lut_4_lut (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(n36448), .O(n22208));   // verilog/i2c_controller.v(89[8] 155[6])
    defparam i26387_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n11_adj_4273));   // verilog/i2c_controller.v(75[27:43])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_CARRY counter2_1516_1517_add_4_3 (.CI(n31695), .I0(GND_net), .I1(counter2[1]), 
            .CO(n31696));
    SB_LUT4 counter2_1516_1517_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n25[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1516_1517_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1516_1517_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n31695));
    SB_LUT4 i26433_2_lut_3_lut (.I0(sda_out), .I1(sda_enable), .I2(n15), 
            .I3(GND_net), .O(n36448));
    defparam i26433_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_4_lut_4_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n37));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h0554;
    SB_LUT4 i30304_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[1] ), 
            .I3(n4760), .O(n37171));
    defparam i30304_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 i1_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n21849));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[1] ), .I1(\state[3] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n34));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h1104;
    SB_LUT4 i56_3_lut_3_lut (.I0(\state[3] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n33));
    defparam i56_3_lut_3_lut.LUT_INIT = 16'h5252;
    SB_LUT4 i1_2_lut_3_lut_adj_1508 (.I0(enable), .I1(i2c_clk), .I2(counter2_7__N_3852), 
            .I3(GND_net), .O(n21937));
    defparam i1_2_lut_3_lut_adj_1508.LUT_INIT = 16'heaea;
    SB_LUT4 i1_4_lut_4_lut_adj_1509 (.I0(\state[0] ), .I1(\state[3] ), .I2(\state[1] ), 
            .I3(\state[2] ), .O(n22149));
    defparam i1_4_lut_4_lut_adj_1509.LUT_INIT = 16'h0316;
    SB_LUT4 state_7__I_0_139_i11_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11));   // verilog/i2c_controller.v(106[5:12])
    defparam state_7__I_0_139_i11_2_lut_4_lut.LUT_INIT = 16'hfffb;
    
endmodule
//
// Verilog Description of module coms
//

module coms (GND_net, n22423, \data_in_frame[14] , clk32MHz, n22422, 
            \data_in_frame[10] , n22421, \data_in_frame[5] , n22420, 
            n22419, n22418, \data_in_frame[15] , n22417, n22416, n22415, 
            n22414, n36883, \data_in_frame[1] , n22413, ID, \data_in_frame[11] , 
            \data_in_frame[12] , \data_in_frame[8] , \data_in_frame[13] , 
            \data_in_frame[9] , rx_data, n22412, \data_in_frame[2] , 
            rx_data_ready, \data_in_frame[21] , n22411, setpoint, \data_in_frame[7] , 
            \data_in_frame[3] , \data_in_frame[6] , \data_in_frame[4] , 
            \data_out_frame[25] , \data_out_frame[19] , \data_out_frame[23] , 
            \data_out_frame[24] , \data_out_frame[15] , \data_out_frame[17] , 
            \data_out_frame[20] , \data_out_frame[18] , n18082, \data_out_frame[16] , 
            \data_out_frame[13] , \data_out_frame[14] , \data_out_frame[12] , 
            \data_out_frame[8] , \data_out_frame[7] , \data_out_frame[5] , 
            \data_out_frame[9] , \data_out_frame[11] , \data_out_frame[10] , 
            \data_out_frame[4] , \data_out_frame[6] , \data_in[2] , \data_in[1] , 
            \data_in[3] , \data_in[0] , tx_active, n35579, n35562, 
            \state[0] , \state[1] , \state[2] , \state[3] , n15, n35561, 
            n35586, n10, n22370, n22369, n22368, n22367, n22366, 
            n22365, n22364, n22363, n22362, control_mode, n22361, 
            n22360, n22359, n22358, n22357, n22356, n22355, PWMLimit, 
            n22354, n22353, n22352, n22351, n22350, n22349, n22348, 
            n22347, n22346, n22345, DE_c, n22344, n22343, n22342, 
            n22341, n22340, LED_c, n35575, n35585, n35568, n22840, 
            IntegralLimit, n22839, n22838, n22837, n22836, n22835, 
            n22834, n22833, n22832, n22831, n22830, n22829, n22828, 
            n22827, n22826, n22825, n22824, n22823, n22822, n22821, 
            n22820, n22819, n22818, n22783, n22782, n22781, n22780, 
            n22779, n22778, n22777, n22776, n22775, n22774, n22773, 
            n22772, n22771, n22770, n22769, n22768, n22767, n22766, 
            n22765, n22764, n22763, n22762, n22761, n22760, n22759, 
            n22758, n22757, n22756, n22755, n22754, n22753, n22752, 
            \Kp[1] , n22751, \Kp[2] , n22750, \Kp[3] , n22749, \Kp[4] , 
            n22748, \Kp[5] , n22747, \Kp[6] , n22746, \Kp[7] , n22745, 
            \Kp[8] , n22744, \Kp[9] , n22743, \Kp[10] , n22742, 
            \Kp[11] , n22741, \Kp[12] , n22740, \Kp[13] , n22739, 
            \Kp[14] , n22738, \Kp[15] , n22737, \Ki[1] , n22736, 
            \Ki[2] , n22735, \Ki[3] , n22734, \Ki[4] , n22733, \Ki[5] , 
            n22732, \Ki[6] , n22731, \Ki[7] , n22730, \Ki[8] , n22729, 
            \Ki[9] , n22728, \Ki[10] , n22727, \Ki[11] , n22726, 
            \Ki[12] , n22725, \Ki[13] , n22724, \Ki[14] , n22721, 
            \Ki[15] , n22720, n22719, n22718, n22717, n22716, n22715, 
            n22714, n22713, n22712, n22711, n22710, n22709, n22708, 
            n22707, n22706, n22705, n22704, n22703, n22702, n22701, 
            n22700, n22699, n22698, n22697, n22696, n22695, n22694, 
            n22693, n22692, n22691, n22690, n22689, n22688, n22687, 
            n22686, n22685, n22684, n22683, n22682, n22681, n22680, 
            n22679, n22678, n22677, n22676, n22675, n22674, n22673, 
            n22672, n22671, n22670, n22669, n22668, n22667, n22666, 
            n22665, n22664, n22663, n22662, n22661, n22660, n22659, 
            n22658, n22657, n22656, n21865, n22339, n22338, n22337, 
            n22336, n22335, n22334, n22333, n22315, n22314, n22312, 
            neopxl_color, n22311, \Ki[0] , n22310, \Kp[0] , n22309, 
            n22655, n22654, n22653, n22652, n22651, n22650, n22649, 
            n22648, n22647, n22646, n22645, n22644, n22643, n22642, 
            n22641, n22640, n22639, n22638, n22637, n22636, n22635, 
            n22634, n22633, n22632, n22631, n22630, n22629, n22628, 
            n22627, n22626, n22625, n22624, n22623, n22622, n22621, 
            n22620, n22619, n22618, n22617, n22616, n22615, n22614, 
            n22613, n22612, n22611, n22610, n22609, n22608, n22607, 
            n22606, n22605, n22604, n22603, n22602, n22601, n22600, 
            n22599, n22598, n22597, n22596, n22595, n22594, n22593, 
            n22592, n22591, n22590, n22589, n22588, n22587, n22586, 
            n22585, n22584, n22583, n22582, n22581, n22580, n22579, 
            n22578, n22577, n22576, n22575, n22574, n22573, n22572, 
            n22571, n22570, n22569, n22568, n22567, n22566, n22565, 
            n22564, n22563, n22292, n22562, n3957, n15_adj_3, scl_enable_N_3958, 
            n22561, n22560, n22559, n22558, n22557, n22556, n22555, 
            n22554, n22553, n22552, n22551, n22550, n22549, n22548, 
            n22547, n22546, n22545, n22544, n22543, n22542, n22541, 
            n22540, n22539, n22538, n22498, n22497, n22496, n22495, 
            n22494, n22493, n22492, n22491, n22490, n22489, n22488, 
            n22487, n22486, n22485, n22484, n22483, n22482, n22481, 
            n22480, n22479, n22478, n22477, n22476, n22475, n5180, 
            n22434, n22433, n22432, n22431, n22430, n22429, n22428, 
            n22427, n22426, n22425, n22424, n21920, n22195, r_SM_Main, 
            \r_SM_Main_2__N_3454[1] , tx_o, n13920, VCC_net, \r_Bit_Index[0] , 
            n4, n22817, n22319, n41168, tx_enable, n22012, n22193, 
            n26980, n4_adj_4, n4_adj_5, \r_Bit_Index[0]_adj_6 , n20781, 
            r_Rx_Data, RX_N_10, n20776, n4_adj_7, n22843, n22847, 
            n22308, n22307, n22306, n22305, n22304, n22303, n22302) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input n22423;
    output [7:0]\data_in_frame[14] ;
    input clk32MHz;
    input n22422;
    output [7:0]\data_in_frame[10] ;
    input n22421;
    output [7:0]\data_in_frame[5] ;
    input n22420;
    input n22419;
    input n22418;
    output [7:0]\data_in_frame[15] ;
    input n22417;
    input n22416;
    input n22415;
    input n22414;
    output n36883;
    output [7:0]\data_in_frame[1] ;
    input n22413;
    input [7:0]ID;
    output [7:0]\data_in_frame[11] ;
    output [7:0]\data_in_frame[12] ;
    output [7:0]\data_in_frame[8] ;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_in_frame[9] ;
    output [7:0]rx_data;
    input n22412;
    output [7:0]\data_in_frame[2] ;
    output rx_data_ready;
    output [7:0]\data_in_frame[21] ;
    input n22411;
    output [23:0]setpoint;
    output [7:0]\data_in_frame[7] ;
    output [7:0]\data_in_frame[3] ;
    output [7:0]\data_in_frame[6] ;
    output [7:0]\data_in_frame[4] ;
    output [7:0]\data_out_frame[25] ;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[24] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[20] ;
    output [7:0]\data_out_frame[18] ;
    output n18082;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[13] ;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[4] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_in[2] ;
    output [7:0]\data_in[1] ;
    output [7:0]\data_in[3] ;
    output [7:0]\data_in[0] ;
    output tx_active;
    output n35579;
    output n35562;
    input \state[0] ;
    input \state[1] ;
    input \state[2] ;
    input \state[3] ;
    output n15;
    output n35561;
    output n35586;
    output n10;
    input n22370;
    input n22369;
    input n22368;
    input n22367;
    input n22366;
    input n22365;
    input n22364;
    input n22363;
    input n22362;
    output [7:0]control_mode;
    input n22361;
    input n22360;
    input n22359;
    input n22358;
    input n22357;
    input n22356;
    input n22355;
    output [23:0]PWMLimit;
    input n22354;
    input n22353;
    input n22352;
    input n22351;
    input n22350;
    input n22349;
    input n22348;
    input n22347;
    input n22346;
    input n22345;
    output DE_c;
    input n22344;
    input n22343;
    input n22342;
    input n22341;
    input n22340;
    output LED_c;
    output n35575;
    output n35585;
    output n35568;
    input n22840;
    output [23:0]IntegralLimit;
    input n22839;
    input n22838;
    input n22837;
    input n22836;
    input n22835;
    input n22834;
    input n22833;
    input n22832;
    input n22831;
    input n22830;
    input n22829;
    input n22828;
    input n22827;
    input n22826;
    input n22825;
    input n22824;
    input n22823;
    input n22822;
    input n22821;
    input n22820;
    input n22819;
    input n22818;
    input n22783;
    input n22782;
    input n22781;
    input n22780;
    input n22779;
    input n22778;
    input n22777;
    input n22776;
    input n22775;
    input n22774;
    input n22773;
    input n22772;
    input n22771;
    input n22770;
    input n22769;
    input n22768;
    input n22767;
    input n22766;
    input n22765;
    input n22764;
    input n22763;
    input n22762;
    input n22761;
    input n22760;
    input n22759;
    input n22758;
    input n22757;
    input n22756;
    input n22755;
    input n22754;
    input n22753;
    input n22752;
    output \Kp[1] ;
    input n22751;
    output \Kp[2] ;
    input n22750;
    output \Kp[3] ;
    input n22749;
    output \Kp[4] ;
    input n22748;
    output \Kp[5] ;
    input n22747;
    output \Kp[6] ;
    input n22746;
    output \Kp[7] ;
    input n22745;
    output \Kp[8] ;
    input n22744;
    output \Kp[9] ;
    input n22743;
    output \Kp[10] ;
    input n22742;
    output \Kp[11] ;
    input n22741;
    output \Kp[12] ;
    input n22740;
    output \Kp[13] ;
    input n22739;
    output \Kp[14] ;
    input n22738;
    output \Kp[15] ;
    input n22737;
    output \Ki[1] ;
    input n22736;
    output \Ki[2] ;
    input n22735;
    output \Ki[3] ;
    input n22734;
    output \Ki[4] ;
    input n22733;
    output \Ki[5] ;
    input n22732;
    output \Ki[6] ;
    input n22731;
    output \Ki[7] ;
    input n22730;
    output \Ki[8] ;
    input n22729;
    output \Ki[9] ;
    input n22728;
    output \Ki[10] ;
    input n22727;
    output \Ki[11] ;
    input n22726;
    output \Ki[12] ;
    input n22725;
    output \Ki[13] ;
    input n22724;
    output \Ki[14] ;
    input n22721;
    output \Ki[15] ;
    input n22720;
    input n22719;
    input n22718;
    input n22717;
    input n22716;
    input n22715;
    input n22714;
    input n22713;
    input n22712;
    input n22711;
    input n22710;
    input n22709;
    input n22708;
    input n22707;
    input n22706;
    input n22705;
    input n22704;
    input n22703;
    input n22702;
    input n22701;
    input n22700;
    input n22699;
    input n22698;
    input n22697;
    input n22696;
    input n22695;
    input n22694;
    input n22693;
    input n22692;
    input n22691;
    input n22690;
    input n22689;
    input n22688;
    input n22687;
    input n22686;
    input n22685;
    input n22684;
    input n22683;
    input n22682;
    input n22681;
    input n22680;
    input n22679;
    input n22678;
    input n22677;
    input n22676;
    input n22675;
    input n22674;
    input n22673;
    input n22672;
    input n22671;
    input n22670;
    input n22669;
    input n22668;
    input n22667;
    input n22666;
    input n22665;
    input n22664;
    input n22663;
    input n22662;
    input n22661;
    input n22660;
    input n22659;
    input n22658;
    input n22657;
    input n22656;
    output n21865;
    input n22339;
    input n22338;
    input n22337;
    input n22336;
    input n22335;
    input n22334;
    input n22333;
    input n22315;
    input n22314;
    input n22312;
    output [23:0]neopxl_color;
    input n22311;
    output \Ki[0] ;
    input n22310;
    output \Kp[0] ;
    input n22309;
    input n22655;
    input n22654;
    input n22653;
    input n22652;
    input n22651;
    input n22650;
    input n22649;
    input n22648;
    input n22647;
    input n22646;
    input n22645;
    input n22644;
    input n22643;
    input n22642;
    input n22641;
    input n22640;
    input n22639;
    input n22638;
    input n22637;
    input n22636;
    input n22635;
    input n22634;
    input n22633;
    input n22632;
    input n22631;
    input n22630;
    input n22629;
    input n22628;
    input n22627;
    input n22626;
    input n22625;
    input n22624;
    input n22623;
    input n22622;
    input n22621;
    input n22620;
    input n22619;
    input n22618;
    input n22617;
    input n22616;
    input n22615;
    input n22614;
    input n22613;
    input n22612;
    input n22611;
    input n22610;
    input n22609;
    input n22608;
    input n22607;
    input n22606;
    input n22605;
    input n22604;
    input n22603;
    input n22602;
    input n22601;
    input n22600;
    input n22599;
    input n22598;
    input n22597;
    input n22596;
    input n22595;
    input n22594;
    input n22593;
    input n22592;
    input n22591;
    input n22590;
    input n22589;
    input n22588;
    input n22587;
    input n22586;
    input n22585;
    input n22584;
    input n22583;
    input n22582;
    input n22581;
    input n22580;
    input n22579;
    input n22578;
    input n22577;
    input n22576;
    input n22575;
    input n22574;
    input n22573;
    input n22572;
    input n22571;
    input n22570;
    input n22569;
    input n22568;
    input n22567;
    input n22566;
    input n22565;
    input n22564;
    input n22563;
    input n22292;
    input n22562;
    output n3957;
    input n15_adj_3;
    output scl_enable_N_3958;
    input n22561;
    input n22560;
    input n22559;
    input n22558;
    input n22557;
    input n22556;
    input n22555;
    input n22554;
    input n22553;
    input n22552;
    input n22551;
    input n22550;
    input n22549;
    input n22548;
    input n22547;
    input n22546;
    input n22545;
    input n22544;
    input n22543;
    input n22542;
    input n22541;
    input n22540;
    input n22539;
    input n22538;
    input n22498;
    input n22497;
    input n22496;
    input n22495;
    input n22494;
    input n22493;
    input n22492;
    input n22491;
    input n22490;
    input n22489;
    input n22488;
    input n22487;
    input n22486;
    input n22485;
    input n22484;
    input n22483;
    input n22482;
    input n22481;
    input n22480;
    input n22479;
    input n22478;
    input n22477;
    input n22476;
    input n22475;
    output n5180;
    input n22434;
    input n22433;
    input n22432;
    input n22431;
    input n22430;
    input n22429;
    input n22428;
    input n22427;
    input n22426;
    input n22425;
    input n22424;
    output n21920;
    output n22195;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3454[1] ;
    output tx_o;
    output n13920;
    input VCC_net;
    output \r_Bit_Index[0] ;
    output n4;
    input n22817;
    input n22319;
    input n41168;
    output tx_enable;
    output n22012;
    output n22193;
    output n26980;
    output n4_adj_4;
    output n4_adj_5;
    output \r_Bit_Index[0]_adj_6 ;
    output n20781;
    output r_Rx_Data;
    input RX_N_10;
    output n20776;
    output n4_adj_7;
    input n22843;
    input n22847;
    input n22308;
    input n22307;
    input n22306;
    input n22305;
    input n22304;
    input n22303;
    input n22302;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    
    wire n11, n35060, n35102, n35098, n35096, n35094, n35092, 
        n35020, n35090, n35088, n35116, n20619;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(115[11:12])
    
    wire n3303, n17948, n18028, n11_adj_3975, n35086, n27759, n35084, 
        n35240, n3, n30684, n30685, n35082, n36265, n36102, n35738, 
        n10_c, n36850, n17985, n1, n20715, n4452, n4_c, n6, 
        n20617, n32519, n36527, n35062;
    wire [7:0]n8825;
    
    wire n21904;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(102[12:33])
    
    wire n22179, n19152, n21454, n31, n18279, n20795, n27040, 
        n4915, Kp_23__N_829;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(96[12:25])
    
    wire n19969, n21045, n27024, n35569, n12, n10_adj_3976, n11_adj_3977, 
        n9, n36060, n32997;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(96[12:25])
    
    wire n36244, n10_adj_3978, n7, n36127, n34001, n36002, n36235, 
        n35644, n21174, n36041, n10_adj_3979;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(96[12:25])
    
    wire n37804;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(96[12:25])
    
    wire n35920, n33952, n10_adj_3980;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(96[12:25])
    
    wire n21149, n35675, n6_adj_3981, n37779, n35834, n36290, n36161, 
        n36253, n10_adj_3982, n36158, n37455, n33843, n10_adj_3983, 
        n6_adj_3984, Kp_23__N_702, n37949, n21212, n36293, n11_adj_3985, 
        n21223, n36315, n35906, n6_adj_3986;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(96[12:25])
    
    wire n36185, n35954, n36189, n37310, n35774, n33879, n33837, 
        n4_adj_3987, n6_adj_3988, n36139, n36308, n30, n35866, n34, 
        n36250, n35900, n32, n6_adj_3989, n38075, n36, n32886, 
        n20891, n31_adj_3990, n18, n35671, n36314, n36262, n21, 
        n35886, n36219, n14, n35893, n36063, n13, n14_adj_3991, 
        Kp_23__N_834, n37847, n15_c, n24, n37930, n19, n20, n36200, 
        n36037, n4_adj_3992, n20951, n12_adj_3993, n36275, n32987, 
        n32855, n32664, Kp_23__N_1151, n20881, n18_adj_3994, n30_adj_3995, 
        n21620, n28, n36081, n35849, n21296, n29, n36084, n36311, 
        n35996, n27, n10_adj_3996, n33890, n14_adj_3997, n21290, 
        n36831, n6_adj_3998, n33950, n35914, n8, n22403, Kp_23__N_1377, 
        Kp_23__N_1162, n35923, n22404, n10_adj_3999, n3_adj_4000, 
        n2, n35154, n22405;
    wire [0:0]n3412;
    wire [2:0]r_SM_Main_2__N_3457;
    
    wire n36486, n12_adj_4001, n21722, n2841, n3_adj_4002, n3_adj_4003, 
        n3_adj_4004, n3_adj_4005, n36005, n21171, n14_adj_4006, n10_adj_4007, 
        n35635, n22406, n8_adj_4008, n3_adj_4009, n22407, n22408, 
        n22409, n5, n3_adj_4010, n3_adj_4011, n3_adj_4012, n3_adj_4013, 
        n3_adj_4014, n3_adj_4015, \FRAME_MATCHER.rx_data_ready_prev , 
        n35046, n35160, n3_adj_4016, n3_adj_4017, n36672, n3_adj_4018, 
        tx_transmit_N_3354, n3_adj_4019, n3_adj_4020, n3_adj_4021, n20900, 
        n3_adj_4022, n3_adj_4023, n3_adj_4024, n21085, n35748, n22410, 
        n3_adj_4025, n3_adj_4026, n3_adj_4027, n3_adj_4028, n3_adj_4029, 
        n3_adj_4030, n4916, n21925, n3_adj_4031, n3_adj_4032, n3_adj_4033, 
        n8_adj_4034, n22395, n22396, n3_adj_4035, n36130, n35709, 
        n14_adj_4036, n10_adj_4037, n36099, n15_adj_4038, n14_adj_4039, 
        n36136, n21815, n12_adj_4040, n35993, n14_adj_4041, n13_adj_4042, 
        n21568, n38298, n36188, n37330, n12_adj_4043, n36215, n10_adj_4044, 
        n22397, n33841, n37418, n63, n63_adj_4045;
    wire [31:0]n92;
    
    wire n33849, n35957, n20844, n8_adj_4046, n35724;
    wire [31:0]\FRAME_MATCHER.state_31__N_2501 ;
    
    wire n7_adj_4047, n20794, n6_adj_4048, n20793, n13961, n8_adj_4049, 
        n35, n35589, n41164, n5_adj_4050, n12_adj_4051, n21479, 
        n33683, n35587, n34_adj_4052, n35789, n20979, n20704, n42, 
        n6_adj_4053, n8_adj_4054, n36078, n36420, n41163, n21060, 
        n6_adj_4055, n30710, n8_adj_4056, n6_adj_4057, n21127, n36069, 
        n35696, n21100, n22398, n2_adj_4058, n30709, n6_adj_4059, 
        n22399, n6_adj_4060, n35114, n33933, Kp_23__N_1147, n11_adj_4061, 
        n35764, n22400, n36075, n33636, n6_adj_4062, n36772, n21048, 
        n35805, n20847, n10_adj_4063, n22401, n10_adj_4064, n16, 
        n36142, n12_adj_4065, n20961, n35624, n35967, n36121, n10_adj_4066, 
        n22402, n21181, n21797, n38098, n8_adj_4067, n24_adj_4068, 
        Kp_23__N_777, n37091, n35687, n22, Kp_23__N_934, n35798, 
        n4_adj_4069, n23, n35730, n21690, n35699, n10_adj_4070, 
        n12_adj_4071, n21436, n35702, n10_adj_4072, n2_adj_4073, n30708, 
        n21_adj_4074, n2_adj_4075, n30707, n35184, n30683, n35647, 
        n2_adj_4076, n30706, n34638, n30705, n6_adj_4077, n37542, 
        n35248, n30682, n3_adj_4078, n33870, n36933, n35889, n10_adj_4079, 
        n32851, n36178, n6_adj_4080, n37877, n33963, n6_adj_4081, 
        n36611, n33893, n32954, n33954, n36986, n35246, n30681, 
        n35945, n21586, n32951, n6_adj_4082, n38149, n35929, n35618, 
        n36278, n35975, n33872, n36066, n33921, n10_adj_4083, n18_adj_4084, 
        n36899, n33007, n36317, n36151, n36268, n12_adj_4085, n35926, 
        n35690, n36247, n36248, n33815, n34646, n30704, n34650, 
        n30703, n7_adj_4086, n33928, n37228, n8_adj_4087, n22387, 
        n32920, n21611, n36090, n6_adj_4088, n37246, n26, n30_adj_4089, 
        n17, n31_adj_4090, n22388, n35118, n35158, n35156, n27009, 
        n35200, n34990, n35186, n35152, n35150, n35148, n35146, 
        n35144, n35142, n35140, n35138, n35100, n35136, n35134, 
        n35132, n35104, n35130, n35106, n27007, n27755, n35128, 
        n35108, n27005, n27753, n35126, n35110, n7_adj_4091, n8_adj_4092, 
        n35124, n35058, n7_adj_4093, n8_adj_4094, n35122, n35112, 
        n35120, n35056, n35048, n35036, n32949, n21278, n35881, 
        n21451, n35904, n21961;
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    
    wire n35897, n36087, n35840, n36272, n35878, n22389, n36207, 
        n35912, n35909, n32_adj_4095, n22_adj_4096, n35716, n36_adj_4097, 
        n35948, n34_adj_4098, n32964, n35_adj_4099, n22390, n22391, 
        n35972, n32876, n33, n22392, Kp_23__N_943, n20771;
    wire [31:0]\FRAME_MATCHER.state_31__N_2565 ;
    
    wire n17814, n36210, n37142, n28068, n27756, n13_adj_4100, n11_adj_4101, 
        n27954, n35863;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(97[12:26])
    
    wire n36761, n36204, n32865, n35871, n36148, n6_adj_4102, n36801, 
        n37037, n35917, n36164, n22393, n34660, n30702, n22394, 
        n8_adj_4103, n6_adj_4104, Kp_23__N_940, n35727, n10_adj_4105, 
        n35684, n35713, n35663, n35802, n35768, n6_adj_4106, n35757, 
        n33327, n32945, n10_adj_4107, n35244, n30680, n35862, n35935, 
        n36115, n10_adj_4108, n36944, n34668, n30701, n35242, n30679, 
        n37644, n2208, n32934, n32942, n161, n35983, n35600, n36014, 
        n34672, n30700, n32867, n36259, n19038, n33064, n10_adj_4109, 
        n34684, n34700, n6_adj_4110, n34722, n34746, n34766, n34790, 
        n34816, n34842, n34866, n34890, n34920, n34940, n34962, 
        n34988, n35022, n33979, n33991, n36008, n33961, n30699, 
        n37273, n35987, n30698, n6_adj_4111, n36011, n32863, n2206, 
        n33986, n6_adj_4112, n20475, n33015, n6_adj_4113, n33939, 
        n36209, n35932, n6_adj_4114, n35777, n10_adj_4115, n36051, 
        n20861, n12_adj_4116, n35656, n35820, n1519, n21789, n35837, 
        n36133, n10_adj_4117, n38156, n21015, n36146, n35980, n36222, 
        n21647, n12_adj_4118, n27129, n28_adj_4119, n26_adj_4120, 
        n27_adj_4121, n36167, n25, n10_adj_4122, n9_adj_4123, n36256, 
        n35615, n36034, n12_adj_4124, n36109, n4_adj_4125, n20703, 
        n35771, n14_adj_4126, n21032, n1168, n15_adj_4127, n4_adj_4128, 
        n35745, n35612, n36228, n14_adj_4129, n9_adj_4130, n21812, 
        n33493, n36212, n14_adj_4131, n20792, n36406, n10_adj_4132, 
        n10_adj_4133, n36027, n36238, n35638, n10_adj_4134, n14_adj_4135, 
        n36105, n36044, n20824, n20_adj_4136, n36302, n32930, n19_adj_4137, 
        n35650, n21026, n21_adj_4138, n6_adj_4139, n21227, n36124, 
        n35629, n36096, n20804, n36030, n33839, n26_adj_4140, n24_adj_4141, 
        n36174, n25_adj_4142, n30697, n23_adj_4143, n37842, n35827, 
        n44, n35681, n43, n49, n35785, n48, n36296, n46, n22386, 
        n22385, n35795, n36112, n47, n45, n54, n53, n40, n38, 
        n39, n22384, n35659, n37, n35_adj_4144, n36057, n36072, 
        n10_adj_4145, n46_adj_4146, n33886, n41, n36_adj_4147, n21333, 
        n36197, n6_adj_4148, n33813, n34025, n4_adj_4149, n16_adj_4150, 
        n22383, n22382, n22381, n36093, n12_adj_4151, n21249, n22_adj_4152, 
        n36194, n36231, n12_adj_4153, n36017, n36024, n21420, n21216, 
        n6_adj_4154, n20789, n35539, n35533, n39281, n38292, n44_adj_4155, 
        n42_adj_4156, n43_adj_4157, n41_adj_4158, n40_adj_4159, n39_adj_4160, 
        n50, n45_adj_4161, n30696, n20713, n20768, n18_adj_4162, 
        n20_adj_4163, n15_adj_4164, n20620, n10_adj_4165, n14_adj_4166, 
        n20762, n10_adj_4167, n38341, n9_adj_4168, n20710, n16_adj_4169, 
        n17_adj_4170, n37965, n12_adj_4171, n37935, n16_adj_4172, 
        n17_adj_4173, n63_adj_4174, n26_adj_4175, n10_adj_4176, n31_adj_4177, 
        n22_adj_4178, n35990, n36225, n30695, n4_adj_4179, n4_adj_4180, 
        n36412, n28158, n8_adj_4181, n35844, n15_adj_4182, n22379, 
        n30694, n35754, n30693, n18_adj_4183, n35780, n18_adj_4184, 
        n27000, n20_adj_4185, n36241, n16_adj_4186, n37915, n30_adj_4187, 
        n35678, n28_adj_4188, n36020, n29_adj_4189, n27_adj_4190, 
        n22380, n36191, n21522, n36305, n6_adj_4191, n35964, n16_adj_4192, 
        n35961, n17_adj_4193, n36287, n10_adj_4194, n20912, n40897, 
        n39278, n40924, n14_adj_4195, n7_adj_4196;
    wire [7:0]tx_data;   // verilog/coms.v(105[13:20])
    
    wire n38348, n38349, n40918, n38358, n38357, n14_adj_4197, n40912, 
        n40915, n40906, n40909, n40900, n40903, n39279, n39280, 
        n40894, n6_adj_4198, n17_adj_4199, n16_adj_4200, n40888, n40891, 
        n40882, n40885, n40876, n40879, n40864, n40867, n40858, 
        n40861, n40852, n40855, n40846, n40849, n10_adj_4201, n40828, 
        n40831, n40816, n40819, n40810, n10_adj_4202, n40813, n40804, 
        n40807, n40798, n40801, n40792, n40795, n40786, n36054, 
        n24_adj_4203, n20_adj_4204, n30692, n40789, n40663, n39274, 
        n40780, n14_adj_4205, n7_adj_4206, n40669, n39263, n40774, 
        n7_adj_4207, n40675, n39260, n40768, n35792, n14_adj_4208, 
        n7_adj_4209, n40681, n39257, n40762, n14_adj_4210, n7_adj_4211, 
        n40687, n39254, n40756, n14_adj_4212, n10_adj_4213, n14_adj_4214, 
        n7_adj_4215, n40693, n39251, n40750, n14_adj_4216, n7_adj_4217, 
        n6_adj_4218, n21240, Kp_23__N_937, n35751, n35578, n6_adj_4219, 
        n35560, n30691, n10_adj_4221, n8_adj_4222, n22499, n22500, 
        n22501, n22502, n22503, n22504, n22505, n22506, n38425, 
        n38423, n7_adj_4223, n6_adj_4224, Kp_23__N_810, n35811, n38419, 
        n38417, n26_adj_4225, n27_adj_4226, n30_adj_4227, n23_adj_4228, 
        n22_adj_4229, n31_adj_4230, n38325, n38413, n38411, n30690, 
        n38407, n38405, n38401, n38399, n4_adj_4231, n6_adj_4232, 
        n38386, n38384, n30689, n38389, n38387, n38395, n38393, 
        n30687, n30688, n22467, n22468, n22469, n22138, n40711, 
        n39248, n40744, n22470, n22471, n7_adj_4234, n23_adj_4235, 
        n22472, n12_adj_4236, n22378, n14_adj_4237, n22128, n22473, 
        n22377, n4917, n22376, n20723, n22474, n37904, n22459, 
        n22460, n5_adj_4238, n6_adj_4239, n35502, n22461, n22462, 
        n22463, n22464, n22465, n10_adj_4240, n22466, n22451, n22452, 
        n22453, n22454, n35814, n14_adj_4241, n22455, n22456, n22457, 
        n22375, n22374, n22373, n22372, n22371, n40738, n37539, 
        n22458, n4902, n36508, n22443, n38079, n4918, n4939, n4938, 
        n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, 
        n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, 
        n4935, n4936, n4937, n26_adj_4242, n22444, n20700, n27_adj_4243, 
        n22445, n22446, n22447, n22448, n22449, n22450, n18_adj_4244, 
        n29_adj_4245, n22435, n22436, n22437, n22438, n38300, n22439, 
        n30686, n22440, n22441, n22442, n40741, n40732, n40735, 
        n36155, n20629, n1_adj_4246, n21440, n22523, n30716, n30715, 
        n22524, n30714, n22313, n22525, n22526, n30713, n22527, 
        n22528, n30712, n22529, n16_adj_4247, n17_adj_4248, n39277, 
        n22530, n39276, n22515, n22516, n16_adj_4250, n17_adj_4251, 
        n30711, n39265, n39264, n22517, n16_adj_4252, n17_adj_4253, 
        n39262, n39261, n16_adj_4254, n17_adj_4255, n39259, n39258, 
        n16_adj_4256, n17_adj_4257, n39256, n39255, n16_adj_4258, 
        n17_adj_4259, n39253, n39252, n16_adj_4260, n17_adj_4261, 
        n22537, n22536, n22535, n22534, n22533, n22518, n22532, 
        n22519, n22531, n22522, n22521, n22520, n22514, n22513, 
        n22512, n39250, n22511, n22510, n22509, n39249, n22508, 
        n22507, n40708, n33831, n40696, n40699, n40690, n40684, 
        n40678, n40672, n40666, n40660, n40648, n40651, n35858, 
        n38412, n38406, n40645, n38400, n40642, n38394, n38385;
    
    SB_LUT4 i1_2_lut (.I0(\FRAME_MATCHER.state [15]), .I1(n11), .I2(GND_net), 
            .I3(GND_net), .O(n35060));
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_843 (.I0(\FRAME_MATCHER.state [16]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35102));
    defparam i1_2_lut_adj_843.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_844 (.I0(\FRAME_MATCHER.state [18]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35098));
    defparam i1_2_lut_adj_844.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_845 (.I0(\FRAME_MATCHER.state [19]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35096));
    defparam i1_2_lut_adj_845.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_846 (.I0(\FRAME_MATCHER.state [20]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35094));
    defparam i1_2_lut_adj_846.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_847 (.I0(\FRAME_MATCHER.state [21]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35092));
    defparam i1_2_lut_adj_847.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n22423));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_848 (.I0(\FRAME_MATCHER.state [22]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35020));
    defparam i1_2_lut_adj_848.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_849 (.I0(\FRAME_MATCHER.state [23]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35090));
    defparam i1_2_lut_adj_849.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_850 (.I0(\FRAME_MATCHER.state [24]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35088));
    defparam i1_2_lut_adj_850.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_851 (.I0(\FRAME_MATCHER.state [25]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35116));
    defparam i1_2_lut_adj_851.LUT_INIT = 16'h8888;
    SB_LUT4 i18768_2_lut (.I0(n20619), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(GND_net), .O(n3303));   // verilog/coms.v(227[9:54])
    defparam i18768_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i30082_3_lut (.I0(n17948), .I1(n18028), .I2(\FRAME_MATCHER.state [2]), 
            .I3(GND_net), .O(n11_adj_3975));
    defparam i30082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_852 (.I0(\FRAME_MATCHER.state [27]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35086));
    defparam i1_2_lut_adj_852.LUT_INIT = 16'h8888;
    SB_LUT4 i19358_2_lut (.I0(\FRAME_MATCHER.state [28]), .I1(n11), .I2(GND_net), 
            .I3(GND_net), .O(n27759));
    defparam i19358_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_853 (.I0(\FRAME_MATCHER.state [29]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35084));
    defparam i1_2_lut_adj_853.LUT_INIT = 16'h8888;
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n35240), .S(n3));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_8 (.CI(n30684), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n30685));
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n22422));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_854 (.I0(\FRAME_MATCHER.state [30]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35082));
    defparam i1_2_lut_adj_854.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut (.I0(\data_in_frame[10] [2]), .I1(n36265), .I2(n36102), 
            .I3(n35738), .O(n10_c));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_855 (.I0(n36850), .I1(n17985), .I2(GND_net), 
            .I3(GND_net), .O(n1));
    defparam i1_2_lut_adj_855.LUT_INIT = 16'h4444;
    SB_LUT4 i18770_2_lut (.I0(n20715), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(GND_net), .O(n4452));   // verilog/coms.v(259[9:58])
    defparam i18770_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i3_3_lut (.I0(n4_c), .I1(n6), .I2(n20617), .I3(GND_net), 
            .O(n32519));
    defparam i3_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i26504_4_lut (.I0(\FRAME_MATCHER.i [31]), .I1(n32519), .I2(n20619), 
            .I3(\FRAME_MATCHER.state [2]), .O(n36527));
    defparam i26504_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i1_2_lut_adj_856 (.I0(\FRAME_MATCHER.state [31]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35062));
    defparam i1_2_lut_adj_856.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n22421));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk32MHz), 
            .E(n21904), .D(n8825[7]), .R(n22179));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk32MHz), 
            .E(n21904), .D(n8825[6]), .R(n22179));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk32MHz), 
            .E(n21904), .D(n8825[5]), .R(n22179));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk32MHz), 
            .E(n21904), .D(n8825[4]), .R(n22179));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk32MHz), 
            .E(n21904), .D(n8825[3]), .R(n22179));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk32MHz), 
            .E(n21904), .D(n8825[2]), .R(n22179));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk32MHz), 
            .E(n21904), .D(n8825[1]), .R(n22179));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_857 (.I0(n19152), .I1(\data_in_frame[5] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n21454));
    defparam i1_2_lut_adj_857.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n22420));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n22419));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n22418));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n22417));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n22416));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n22415));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n22414));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(n31), .I1(n18279), .I2(n20795), .I3(n27040), 
            .O(n36883));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1315_2_lut_3_lut (.I0(n31), .I1(n18279), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n4915));
    defparam i1315_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i2_3_lut (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_829), .I2(\data_in_frame[0] [5]), 
            .I3(GND_net), .O(n19969));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_858 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[1] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n21045));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_858.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n22413));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut (.I0(n27024), .I1(\FRAME_MATCHER.i [5]), .I2(\FRAME_MATCHER.i [4]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n35569));   // verilog/coms.v(154[7:23])
    defparam i3_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i4_4_lut_adj_859 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [6]), 
            .I2(ID[4]), .I3(ID[6]), .O(n12));   // verilog/coms.v(238[12:32])
    defparam i4_4_lut_adj_859.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_4_lut (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(ID[1]), .I3(ID[2]), .O(n10_adj_3976));   // verilog/coms.v(238[12:32])
    defparam i2_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i3_4_lut_adj_860 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(ID[7]), .I3(ID[5]), .O(n11_adj_3977));   // verilog/coms.v(238[12:32])
    defparam i3_4_lut_adj_860.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [3]), 
            .I2(ID[0]), .I3(ID[3]), .O(n9));   // verilog/coms.v(238[12:32])
    defparam i1_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i7_4_lut (.I0(n9), .I1(n11_adj_3977), .I2(n10_adj_3976), .I3(n12), 
            .O(n18279));   // verilog/coms.v(238[12:32])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_861 (.I0(n36060), .I1(n32997), .I2(\data_in_frame[19] [0]), 
            .I3(n36244), .O(n10_adj_3978));
    defparam i4_4_lut_adj_861.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_862 (.I0(n7), .I1(\data_in_frame[11] [4]), .I2(n36127), 
            .I3(n34001), .O(n36002));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_862.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_863 (.I0(n36235), .I1(n35644), .I2(n21174), .I3(n36041), 
            .O(n10_adj_3979));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_863.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_864 (.I0(\data_in_frame[16] [4]), .I1(n37804), 
            .I2(\data_in_frame[18] [5]), .I3(GND_net), .O(n35920));
    defparam i2_3_lut_adj_864.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_865 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[16] [6]), 
            .I2(\data_in_frame[12] [3]), .I3(n33952), .O(n10_adj_3980));
    defparam i4_4_lut_adj_865.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_866 (.I0(\data_in_frame[17] [0]), .I1(n21149), 
            .I2(n35675), .I3(n6_adj_3981), .O(n37779));
    defparam i4_4_lut_adj_866.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_867 (.I0(\data_in_frame[8] [1]), .I1(n35834), .I2(\data_in_frame[10] [3]), 
            .I3(GND_net), .O(n21174));
    defparam i2_3_lut_adj_867.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_868 (.I0(\data_in_frame[14] [3]), .I1(n36290), 
            .I2(n36161), .I3(n36253), .O(n10_adj_3982));
    defparam i4_4_lut_adj_868.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_869 (.I0(n36158), .I1(\data_in_frame[12] [4]), 
            .I2(n37804), .I3(n21174), .O(n32997));
    defparam i3_4_lut_adj_869.LUT_INIT = 16'h9669;
    SB_LUT4 i3_3_lut_adj_870 (.I0(\data_in_frame[16] [0]), .I1(n37455), 
            .I2(n33843), .I3(GND_net), .O(n10_adj_3983));   // verilog/coms.v(70[16:27])
    defparam i3_3_lut_adj_870.LUT_INIT = 16'h9696;
    SB_LUT4 i2_4_lut_adj_871 (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[19] [2]), 
            .I2(\data_in_frame[19] [5]), .I3(\data_in_frame[19] [1]), .O(n6_adj_3984));   // verilog/coms.v(268[9:85])
    defparam i2_4_lut_adj_871.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_872 (.I0(\data_in_frame[19] [3]), .I1(n6_adj_3984), 
            .I2(\data_in_frame[19] [7]), .I3(\data_in_frame[19] [6]), .O(Kp_23__N_702));   // verilog/coms.v(268[9:85])
    defparam i3_4_lut_adj_872.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_873 (.I0(n37949), .I1(n37779), .I2(GND_net), 
            .I3(GND_net), .O(n21212));   // verilog/coms.v(268[9:85])
    defparam i1_2_lut_adj_873.LUT_INIT = 16'h6666;
    SB_LUT4 i4_3_lut (.I0(n36293), .I1(n21212), .I2(Kp_23__N_702), .I3(GND_net), 
            .O(n11_adj_3985));
    defparam i4_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut (.I0(n11_adj_3985), .I1(n21223), .I2(n10_adj_3983), 
            .I3(n36315), .O(n35906));
    defparam i6_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_874 (.I0(\data_in_frame[18] [7]), .I1(n32997), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3986));
    defparam i1_2_lut_adj_874.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_875 (.I0(\data_in_frame[20] [5]), .I1(n36185), 
            .I2(n35954), .I3(n36189), .O(n37310));
    defparam i3_4_lut_adj_875.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_876 (.I0(\data_in_frame[14] [5]), .I1(n37779), 
            .I2(n35774), .I3(n6_adj_3986), .O(n33879));
    defparam i4_4_lut_adj_876.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_877 (.I0(n33837), .I1(\data_in_frame[14] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_3987));
    defparam i1_2_lut_adj_877.LUT_INIT = 16'h9999;
    SB_LUT4 i2_4_lut_adj_878 (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[16] [4]), 
            .I2(\data_in_frame[18] [7]), .I3(n4_adj_3987), .O(n36244));   // verilog/coms.v(78[16:27])
    defparam i2_4_lut_adj_878.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_879 (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3988));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_879.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_880 (.I0(\data_in_frame[12] [7]), .I1(\data_in_frame[15] [1]), 
            .I2(\data_in_frame[13] [1]), .I3(n6_adj_3988), .O(n36041));   // verilog/coms.v(71[16:27])
    defparam i4_4_lut_adj_880.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_881 (.I0(\data_in_frame[16] [6]), .I1(\data_in_frame[16] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n35774));
    defparam i1_2_lut_adj_881.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_882 (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[14] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n36139));
    defparam i1_2_lut_adj_882.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_883 (.I0(\data_in_frame[11] [7]), .I1(\data_in_frame[9] [5]), 
            .I2(\data_in_frame[10] [1]), .I3(GND_net), .O(n36161));
    defparam i2_3_lut_adj_883.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut (.I0(n36308), .I1(\data_in_frame[11] [0]), .I2(\data_in_frame[9] [7]), 
            .I3(n36161), .O(n30));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut (.I0(n35866), .I1(n30), .I2(\data_in_frame[10] [3]), 
            .I3(\data_in_frame[10] [4]), .O(n34));
    defparam i15_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i13_4_lut (.I0(n36250), .I1(\data_in_frame[10] [6]), .I2(n35900), 
            .I3(\data_in_frame[11] [5]), .O(n32));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut (.I0(\data_in_frame[9] [3]), .I1(n34), .I2(n6_adj_3989), 
            .I3(n38075), .O(n36));
    defparam i17_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut (.I0(n32886), .I1(\data_in_frame[11] [3]), .I2(\data_in_frame[10] [2]), 
            .I3(n20891), .O(n31_adj_3990));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut (.I0(n31_adj_3990), .I1(\data_in_frame[12] [0]), .I2(n36), 
            .I3(n32), .O(n18));
    defparam i5_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_884 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35671));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_884.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut (.I0(n36314), .I1(\data_in_frame[14] [3]), .I2(n36262), 
            .I3(\data_in_frame[14] [0]), .O(n21));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_885 (.I0(n35886), .I1(n36219), .I2(n36185), .I3(n36139), 
            .O(n14));
    defparam i6_4_lut_adj_885.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_886 (.I0(n35774), .I1(n35893), .I2(n36063), .I3(n36041), 
            .O(n13));
    defparam i5_4_lut_adj_886.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_887 (.I0(\data_in_frame[14] [1]), .I1(\data_in_frame[15] [3]), 
            .I2(n13), .I3(n14), .O(n14_adj_3991));
    defparam i5_4_lut_adj_887.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_888 (.I0(\data_in_frame[1] [3]), .I1(n35671), .I2(Kp_23__N_834), 
            .I3(n21045), .O(Kp_23__N_829));   // verilog/coms.v(70[16:69])
    defparam i3_4_lut_adj_888.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_889 (.I0(\data_in_frame[12] [1]), .I1(n37847), 
            .I2(\data_in_frame[14] [6]), .I3(\data_in_frame[17] [0]), .O(n15_c));
    defparam i6_4_lut_adj_889.LUT_INIT = 16'h9669;
    SB_LUT4 i11_4_lut_adj_890 (.I0(n21), .I1(\data_in_frame[18] [5]), .I2(n18), 
            .I3(\data_in_frame[14] [2]), .O(n24));
    defparam i11_4_lut_adj_890.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_891 (.I0(n15_c), .I1(\data_in_frame[13] [3]), .I2(n14_adj_3991), 
            .I3(\data_in_frame[11] [4]), .O(n37930));
    defparam i8_4_lut_adj_891.LUT_INIT = 16'h6996;
    SB_LUT4 i6_2_lut (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[17] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n19));
    defparam i6_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i28_4_lut (.I0(n19), .I1(n37930), .I2(n24), .I3(n20), .O(n36315));
    defparam i28_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_892 (.I0(\data_in_frame[8] [0]), .I1(n36200), .I2(n36037), 
            .I3(n4_adj_3992), .O(n36290));   // verilog/coms.v(75[16:27])
    defparam i3_4_lut_adj_892.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_893 (.I0(n36290), .I1(\data_in_frame[10] [1]), 
            .I2(\data_in_frame[9] [7]), .I3(GND_net), .O(n35893));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_893.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_894 (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n20951));
    defparam i1_2_lut_adj_894.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_895 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n21149));
    defparam i1_2_lut_adj_895.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_896 (.I0(\data_in_frame[12] [6]), .I1(n36158), 
            .I2(\data_in_frame[17] [1]), .I3(n21149), .O(n12_adj_3993));
    defparam i5_4_lut_adj_896.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_897 (.I0(n20951), .I1(n12_adj_3993), .I2(n36275), 
            .I3(\data_in_frame[14] [7]), .O(n37847));
    defparam i6_4_lut_adj_897.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_898 (.I0(n32987), .I1(n32855), .I2(\data_in_frame[12] [1]), 
            .I3(GND_net), .O(n36253));
    defparam i2_3_lut_adj_898.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_899 (.I0(n32664), .I1(\data_in_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n32886));
    defparam i1_2_lut_adj_899.LUT_INIT = 16'h6666;
    SB_LUT4 i13_4_lut_adj_900 (.I0(Kp_23__N_1151), .I1(\data_in_frame[11] [6]), 
            .I2(n20881), .I3(n18_adj_3994), .O(n30_adj_3995));
    defparam i13_4_lut_adj_900.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_901 (.I0(n21620), .I1(n32886), .I2(\data_in_frame[9] [6]), 
            .I3(n36253), .O(n28));
    defparam i11_4_lut_adj_901.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_902 (.I0(n36081), .I1(n19152), .I2(n35849), 
            .I3(n21296), .O(n29));
    defparam i12_4_lut_adj_902.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut (.I0(n36084), .I1(n36311), .I2(\data_in_frame[9] [0]), 
            .I3(n35996), .O(n27));
    defparam i10_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut (.I0(n27), .I1(n29), .I2(n28), .I3(n30_adj_3995), 
            .O(n33837));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut (.I0(n36127), .I1(\data_in_frame[13] [6]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_3996));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_903 (.I0(n36262), .I1(n33890), .I2(\data_in_frame[16] [2]), 
            .I3(\data_in_frame[11] [5]), .O(n14_adj_3997));
    defparam i6_4_lut_adj_903.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_904 (.I0(\data_in_frame[16] [1]), .I1(n14_adj_3997), 
            .I2(n10_adj_3996), .I3(n21290), .O(n36831));
    defparam i7_4_lut_adj_904.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_905 (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[14] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3998));
    defparam i1_2_lut_adj_905.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_906 (.I0(n33950), .I1(n33837), .I2(n35914), .I3(n6_adj_3998), 
            .O(n36314));
    defparam i4_4_lut_adj_906.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_907 (.I0(\data_in_frame[16] [2]), .I1(n36314), 
            .I2(GND_net), .I3(GND_net), .O(n35954));
    defparam i1_2_lut_adj_907.LUT_INIT = 16'h6666;
    SB_LUT4 i14000_3_lut_4_lut (.I0(n8), .I1(n35569), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n22403));
    defparam i14000_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_908 (.I0(\data_in_frame[18] [3]), .I1(n36831), 
            .I2(\data_in_frame[16] [3]), .I3(GND_net), .O(n36185));
    defparam i2_3_lut_adj_908.LUT_INIT = 16'h6969;
    SB_LUT4 i1_3_lut (.I0(\data_in_frame[11] [2]), .I1(\data_in_frame[9] [1]), 
            .I2(\data_in_frame[9] [0]), .I3(GND_net), .O(n6_adj_3989));   // verilog/coms.v(72[16:41])
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_909 (.I0(Kp_23__N_1377), .I1(Kp_23__N_1151), .I2(Kp_23__N_1162), 
            .I3(n6_adj_3989), .O(n35923));   // verilog/coms.v(72[16:41])
    defparam i4_4_lut_adj_909.LUT_INIT = 16'h6996;
    SB_LUT4 i14001_3_lut_4_lut (.I0(n8), .I1(n35569), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n22404));
    defparam i14001_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_910 (.I0(\data_in_frame[18] [1]), .I1(n35923), 
            .I2(\data_in_frame[18] [2]), .I3(GND_net), .O(n35886));
    defparam i2_3_lut_adj_910.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_911 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[13] [4]), 
            .I2(\data_in_frame[16] [1]), .I3(\data_in_frame[11] [6]), .O(n10_adj_3999));
    defparam i4_4_lut_adj_911.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [27]), 
            .I3(GND_net), .O(n35154));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i14002_3_lut_4_lut (.I0(n8), .I1(n35569), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n22405));
    defparam i14002_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_912 (.I0(\data_in_frame[14] [6]), .I1(n33952), 
            .I2(GND_net), .I3(GND_net), .O(n35675));
    defparam i1_2_lut_adj_912.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_913 (.I0(\data_in_frame[12] [6]), .I1(\data_in_frame[12] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n36235));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_913.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_914 (.I0(\data_in_frame[13] [0]), .I1(\data_in_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n36063));
    defparam i1_2_lut_adj_914.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n22412));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSR tx_transmit_3871 (.Q(r_SM_Main_2__N_3457[0]), .C(clk32MHz), 
            .D(n3412[0]), .R(n36486));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_4_lut_adj_915 (.I0(n36063), .I1(n36235), .I2(\data_in_frame[15] [1]), 
            .I3(n35675), .O(n12_adj_4001));
    defparam i5_4_lut_adj_915.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_916 (.I0(\data_in_frame[12] [4]), .I1(n12_adj_4001), 
            .I2(n36275), .I3(n21722), .O(n37949));
    defparam i6_4_lut_adj_916.LUT_INIT = 16'h6996;
    SB_LUT4 select_400_Select_1_i3_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4002));
    defparam select_400_Select_1_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_2_i3_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4003));
    defparam select_400_Select_2_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_3_i3_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4004));
    defparam select_400_Select_3_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_4_i3_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4005));
    defparam select_400_Select_4_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_917 (.I0(n36005), .I1(\data_in_frame[12] [6]), 
            .I2(n21171), .I3(\data_in_frame[15] [2]), .O(n14_adj_4006));
    defparam i6_4_lut_adj_917.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_918 (.I0(\data_in_frame[17] [4]), .I1(n14_adj_4006), 
            .I2(n10_adj_4007), .I3(n35635), .O(n37455));
    defparam i7_4_lut_adj_918.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_919 (.I0(n37455), .I1(n37949), .I2(GND_net), 
            .I3(GND_net), .O(n21223));   // verilog/coms.v(268[9:85])
    defparam i1_2_lut_adj_919.LUT_INIT = 16'h6666;
    SB_LUT4 i14003_3_lut_4_lut (.I0(n8), .I1(n35569), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n22406));
    defparam i14003_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_adj_920 (.I0(n37847), .I1(\data_in_frame[19] [3]), 
            .I2(\data_in_frame[19] [4]), .I3(GND_net), .O(n8_adj_4008));
    defparam i3_3_lut_adj_920.LUT_INIT = 16'h6969;
    SB_LUT4 select_400_Select_5_i3_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4009));
    defparam select_400_Select_5_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14004_3_lut_4_lut (.I0(n8), .I1(n35569), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n22407));
    defparam i14004_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14005_3_lut_4_lut (.I0(n8), .I1(n35569), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n22408));
    defparam i14005_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14006_3_lut_4_lut (.I0(n8), .I1(n35569), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n22409));
    defparam i14006_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_921 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n5));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_adj_921.LUT_INIT = 16'h9696;
    SB_LUT4 select_400_Select_6_i3_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4010));
    defparam select_400_Select_6_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_7_i3_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4011));
    defparam select_400_Select_7_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_8_i3_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4012));
    defparam select_400_Select_8_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_9_i3_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4013));
    defparam select_400_Select_9_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_10_i3_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4014));
    defparam select_400_Select_10_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_11_i3_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4015));
    defparam select_400_Select_11_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3872  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state [0]), .C(clk32MHz), 
            .D(n35046), .S(n35160));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_400_Select_12_i3_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4016));
    defparam select_400_Select_12_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_13_i3_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4017));
    defparam select_400_Select_13_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_922 (.I0(n33879), .I1(n35906), .I2(\data_in_frame[21] [1]), 
            .I3(GND_net), .O(n36672));
    defparam i2_3_lut_adj_922.LUT_INIT = 16'h9696;
    SB_LUT4 select_400_Select_14_i3_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4018));
    defparam select_400_Select_14_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3971_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3354), .I3(GND_net), .O(n8825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 select_400_Select_15_i3_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4019));
    defparam select_400_Select_15_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_16_i3_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4020));
    defparam select_400_Select_16_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_17_i3_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4021));
    defparam select_400_Select_17_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_4_lut_adj_923 (.I0(n20900), .I1(\data_in_frame[1] [3]), .I2(n36102), 
            .I3(n4_adj_3992), .O(n35834));   // verilog/coms.v(75[16:27])
    defparam i3_4_lut_adj_923.LUT_INIT = 16'h6996;
    SB_LUT4 select_400_Select_18_i3_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4022));
    defparam select_400_Select_18_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_19_i3_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4023));
    defparam select_400_Select_19_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_20_i3_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4024));
    defparam select_400_Select_20_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_924 (.I0(n21085), .I1(\data_in_frame[9] [2]), .I2(GND_net), 
            .I3(GND_net), .O(n35748));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_924.LUT_INIT = 16'h6666;
    SB_LUT4 i14007_3_lut_4_lut (.I0(n8), .I1(n35569), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n22410));
    defparam i14007_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n22411));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_400_Select_21_i3_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4025));
    defparam select_400_Select_21_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_22_i3_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4026));
    defparam select_400_Select_22_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_23_i3_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4027));
    defparam select_400_Select_23_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_24_i3_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4028));
    defparam select_400_Select_24_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_25_i3_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4029));
    defparam select_400_Select_25_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_26_i3_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4030));
    defparam select_400_Select_26_i3_2_lut.LUT_INIT = 16'h8888;
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .E(n21925), .D(n4916));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_400_Select_27_i3_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4031));
    defparam select_400_Select_27_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_28_i3_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4032));
    defparam select_400_Select_28_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_400_Select_29_i3_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4033));
    defparam select_400_Select_29_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13992_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35569), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n22395));
    defparam i13992_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13993_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35569), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n22396));
    defparam i13993_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n22410));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 select_400_Select_30_i3_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4035));
    defparam select_400_Select_30_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_925 (.I0(n35834), .I1(n36130), .I2(n36308), .I3(n35709), 
            .O(n14_adj_4036));
    defparam i6_4_lut_adj_925.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_926 (.I0(n36265), .I1(n14_adj_4036), .I2(n10_adj_4037), 
            .I3(\data_in_frame[9] [6]), .O(n38075));
    defparam i7_4_lut_adj_926.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_927 (.I0(\data_in_frame[7] [7]), .I1(n38075), .I2(n35748), 
            .I3(n36099), .O(n15_adj_4038));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_927.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut_adj_928 (.I0(n15_adj_4038), .I1(\data_in_frame[8] [3]), 
            .I2(n14_adj_4039), .I3(\data_in_frame[8] [2]), .O(n36311));   // verilog/coms.v(74[16:43])
    defparam i8_4_lut_adj_928.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_929 (.I0(n36136), .I1(n21815), .I2(\data_in_frame[11] [7]), 
            .I3(n21454), .O(n12_adj_4040));
    defparam i5_4_lut_adj_929.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_930 (.I0(\data_in_frame[14] [1]), .I1(n12_adj_4040), 
            .I2(n36311), .I3(\data_in_frame[13] [7]), .O(n35914));
    defparam i6_4_lut_adj_930.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_931 (.I0(n35993), .I1(n36315), .I2(\data_in_frame[16] [3]), 
            .I3(\data_in_frame[20] [7]), .O(n14_adj_4041));
    defparam i6_4_lut_adj_931.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_932 (.I0(Kp_23__N_702), .I1(n35920), .I2(n21290), 
            .I3(\data_in_frame[19] [0]), .O(n13_adj_4042));
    defparam i5_4_lut_adj_932.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1377));   // verilog/coms.v(70[16:27])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i28271_4_lut (.I0(\data_in_frame[21] [5]), .I1(n36672), .I2(n8_adj_4008), 
            .I3(n21568), .O(n38298));
    defparam i28271_4_lut.LUT_INIT = 16'h8448;
    SB_LUT4 i3_4_lut_adj_933 (.I0(\data_in_frame[20] [6]), .I1(n36188), 
            .I2(n35954), .I3(n35920), .O(n37330));
    defparam i3_4_lut_adj_933.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_934 (.I0(\data_in_frame[19] [7]), .I1(n10_adj_3983), 
            .I2(\data_in_frame[15] [7]), .I3(\data_in_frame[19] [6]), .O(n12_adj_4043));   // verilog/coms.v(70[16:27])
    defparam i5_4_lut_adj_934.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_935 (.I0(n36002), .I1(\data_in_frame[20] [2]), 
            .I2(\data_in_frame[15] [6]), .I3(n36215), .O(n10_adj_4044));
    defparam i4_4_lut_adj_935.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n22409));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13994_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35569), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n22397));
    defparam i13994_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_936 (.I0(\data_in_frame[20] [0]), .I1(n12_adj_4043), 
            .I2(n36002), .I3(n33841), .O(n37418));   // verilog/coms.v(70[16:27])
    defparam i6_4_lut_adj_936.LUT_INIT = 16'h9669;
    SB_LUT4 i18809_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n63), .I2(n63_adj_4045), 
            .I3(GND_net), .O(n92[2]));   // verilog/coms.v(139[4] 141[7])
    defparam i18809_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 i1_2_lut_adj_937 (.I0(\data_in_frame[11] [4]), .I1(\data_in_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35900));
    defparam i1_2_lut_adj_937.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_938 (.I0(\data_in_frame[14] [0]), .I1(n33849), 
            .I2(GND_net), .I3(GND_net), .O(n35957));
    defparam i1_2_lut_adj_938.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_939 (.I0(n20844), .I1(n35957), .I2(n35900), .I3(Kp_23__N_1377), 
            .O(n36188));
    defparam i3_4_lut_adj_939.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_940 (.I0(n33950), .I1(n35914), .I2(GND_net), 
            .I3(GND_net), .O(n21290));
    defparam i1_2_lut_adj_940.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_941 (.I0(n33879), .I1(n37779), .I2(\data_in_frame[19] [2]), 
            .I3(\data_in_frame[19] [1]), .O(n8_adj_4046));
    defparam i3_4_lut_adj_941.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_942 (.I0(n21296), .I1(Kp_23__N_829), .I2(GND_net), 
            .I3(GND_net), .O(n35724));   // verilog/coms.v(71[16:69])
    defparam i1_2_lut_adj_942.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_943 (.I0(\FRAME_MATCHER.state_31__N_2501 [2]), .I1(n7_adj_4047), 
            .I2(n20794), .I3(n3303), .O(n6_adj_4048));
    defparam i1_4_lut_adj_943.LUT_INIT = 16'hcfce;
    SB_LUT4 i3_4_lut_adj_944 (.I0(n20793), .I1(n6_adj_4048), .I2(n13961), 
            .I3(n92[2]), .O(n8_adj_4049));
    defparam i3_4_lut_adj_944.LUT_INIT = 16'hdccc;
    SB_LUT4 i4_4_lut_adj_945 (.I0(\FRAME_MATCHER.state_31__N_2501 [2]), .I1(n8_adj_4049), 
            .I2(n35), .I3(n35589), .O(n41164));
    defparam i4_4_lut_adj_945.LUT_INIT = 16'hefcf;
    SB_LUT4 i5_4_lut_adj_946 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[13] [3]), 
            .I2(n5_adj_4050), .I3(\data_in_frame[9] [1]), .O(n12_adj_4051));   // verilog/coms.v(75[16:43])
    defparam i5_4_lut_adj_946.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_947 (.I0(Kp_23__N_1162), .I1(n12_adj_4051), .I2(n35635), 
            .I3(n21479), .O(n33683));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_947.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_948 (.I0(\data_in_frame[15] [4]), .I1(n33683), 
            .I2(GND_net), .I3(GND_net), .O(n34001));
    defparam i1_2_lut_adj_948.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n22408));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_adj_949 (.I0(n20794), .I1(n3303), .I2(n35587), .I3(GND_net), 
            .O(n34_adj_4052));
    defparam i1_3_lut_adj_949.LUT_INIT = 16'h5454;
    SB_LUT4 i3_4_lut_adj_950 (.I0(\data_in_frame[10] [6]), .I1(n35789), 
            .I2(\data_in_frame[10] [5]), .I3(n20979), .O(n21722));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_950.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_951 (.I0(n35587), .I1(n4452), .I2(n35589), .I3(n20704), 
            .O(n42));
    defparam i1_4_lut_adj_951.LUT_INIT = 16'ha0a2;
    SB_LUT4 i2_4_lut_adj_952 (.I0(n34_adj_4052), .I1(n20793), .I2(n92[1]), 
            .I3(n13961), .O(n6_adj_4053));
    defparam i2_4_lut_adj_952.LUT_INIT = 16'hbabb;
    SB_LUT4 i1_4_lut_adj_953 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[11] [1]), 
            .I2(n8_adj_4054), .I3(n36078), .O(n36005));
    defparam i1_4_lut_adj_953.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_954 (.I0(\FRAME_MATCHER.state [3]), .I1(n6_adj_4053), 
            .I2(n42), .I3(n36420), .O(n41163));
    defparam i3_4_lut_adj_954.LUT_INIT = 16'hfcfe;
    SB_LUT4 i1_2_lut_adj_955 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n21060));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_955.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_956 (.I0(\data_in_frame[7] [4]), .I1(\data_in_frame[5] [3]), 
            .I2(\data_in_frame[5] [2]), .I3(GND_net), .O(n36081));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_956.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_957 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n35996));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_957.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_958 (.I0(\data_in_frame[9] [5]), .I1(n20891), .I2(n35996), 
            .I3(n6_adj_4055), .O(n35866));   // verilog/coms.v(85[17:63])
    defparam i4_4_lut_adj_958.LUT_INIT = 16'h6996;
    SB_CARRY add_3971_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3354), 
            .CO(n30710));
    SB_LUT4 i1_2_lut_adj_959 (.I0(n21085), .I1(n8_adj_4056), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1162));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_959.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_960 (.I0(n35724), .I1(\data_in_frame[3] [0]), .I2(n5), 
            .I3(n6_adj_4057), .O(n21127));   // verilog/coms.v(77[16:27])
    defparam i4_4_lut_adj_960.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_961 (.I0(\data_in_frame[8] [7]), .I1(n36069), .I2(n35696), 
            .I3(\data_in_frame[8] [6]), .O(Kp_23__N_1151));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_961.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_962 (.I0(\data_in_frame[9] [0]), .I1(Kp_23__N_1151), 
            .I2(GND_net), .I3(GND_net), .O(n21815));
    defparam i1_2_lut_adj_962.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_963 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n20891));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_963.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_964 (.I0(n21085), .I1(n21100), .I2(GND_net), 
            .I3(GND_net), .O(n35709));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_adj_964.LUT_INIT = 16'h6666;
    SB_LUT4 i13995_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35569), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n22398));
    defparam i13995_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_33_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [31]), 
            .I2(GND_net), .I3(n30709), .O(n2_adj_4058)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13996_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35569), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n22399));
    defparam i13996_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_965 (.I0(\data_in_frame[18] [0]), .I1(n21479), 
            .I2(n6_adj_4060), .I3(n35709), .O(n36215));
    defparam i1_4_lut_adj_965.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_966 (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[15] [7]), 
            .I2(n36215), .I3(GND_net), .O(n36293));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_966.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_8_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n30684), .O(n35114)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_967 (.I0(n21127), .I1(\data_in_frame[10] [7]), 
            .I2(n32855), .I3(GND_net), .O(n33933));
    defparam i2_3_lut_adj_967.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_9__7__I_0_2_lut (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1147));   // verilog/coms.v(85[17:28])
    defparam data_in_frame_9__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_968 (.I0(n11_adj_4061), .I1(\data_in_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n35764));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_968.LUT_INIT = 16'h6666;
    SB_LUT4 i13997_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35569), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n22400));
    defparam i13997_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_969 (.I0(\data_in_frame[11] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n36075));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_adj_969.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_970 (.I0(n33636), .I1(\data_in_frame[6] [0]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4062));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_970.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_971 (.I0(\data_in_frame[19] [3]), .I1(n21212), 
            .I2(\data_in_frame[21] [4]), .I3(\data_in_frame[19] [2]), .O(n36772));   // verilog/coms.v(268[9:85])
    defparam i3_4_lut_adj_971.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_972 (.I0(n33843), .I1(n36293), .I2(\data_in_frame[16] [0]), 
            .I3(GND_net), .O(n35993));
    defparam i2_3_lut_adj_972.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_973 (.I0(\data_in_frame[6] [2]), .I1(n21048), .I2(n35805), 
            .I3(n6_adj_4062), .O(n35849));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_973.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_974 (.I0(n36075), .I1(n20847), .I2(\data_in_frame[13] [3]), 
            .I3(n36250), .O(n10_adj_4063));
    defparam i4_4_lut_adj_974.LUT_INIT = 16'h6996;
    SB_LUT4 i13998_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35569), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n22401));
    defparam i13998_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_975 (.I0(n35866), .I1(n35764), .I2(n10_adj_4063), 
            .I3(n33849), .O(n10_adj_4064));
    defparam i1_4_lut_adj_975.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_976 (.I0(n21085), .I1(\data_in_frame[17] [7]), 
            .I2(\data_in_frame[15] [7]), .I3(n10_adj_4064), .O(n16));
    defparam i7_4_lut_adj_976.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_977 (.I0(n36142), .I1(n16), .I2(n12_adj_4065), 
            .I3(n21060), .O(n33841));
    defparam i8_4_lut_adj_977.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_978 (.I0(\data_in_frame[13] [1]), .I1(n36219), 
            .I2(n36005), .I3(n21722), .O(n20961));
    defparam i3_4_lut_adj_978.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_979 (.I0(\data_in_frame[7] [5]), .I1(n21296), .I2(n35624), 
            .I3(GND_net), .O(n36037));   // verilog/coms.v(70[16:69])
    defparam i2_3_lut_adj_979.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_980 (.I0(n35967), .I1(\data_in_frame[5] [7]), .I2(\data_in_frame[8] [2]), 
            .I3(n36121), .O(n10_adj_4066));   // verilog/coms.v(76[16:43])
    defparam i4_4_lut_adj_980.LUT_INIT = 16'h6996;
    SB_LUT4 i13999_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35569), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n22402));
    defparam i13999_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_981 (.I0(\data_in_frame[5] [6]), .I1(n21181), .I2(GND_net), 
            .I3(GND_net), .O(n35967));
    defparam i1_2_lut_adj_981.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_982 (.I0(\data_in_frame[1] [4]), .I1(n36037), .I2(\data_in_frame[1] [3]), 
            .I3(GND_net), .O(n32855));   // verilog/coms.v(70[16:69])
    defparam i2_3_lut_adj_982.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_983 (.I0(n21797), .I1(n35849), .I2(GND_net), 
            .I3(GND_net), .O(n36136));
    defparam i1_2_lut_adj_983.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut_adj_984 (.I0(n38098), .I1(\data_in_frame[20] [1]), 
            .I2(n8_adj_4067), .I3(\data_in_frame[19] [7]), .O(n24_adj_4068));
    defparam i8_4_lut_adj_984.LUT_INIT = 16'hbeeb;
    SB_LUT4 i1_2_lut_adj_985 (.I0(\data_in_frame[6] [1]), .I1(Kp_23__N_777), 
            .I2(GND_net), .I3(GND_net), .O(n36121));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_985.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_986 (.I0(n37091), .I1(\data_in_frame[21] [2]), 
            .I2(n35687), .I3(\data_in_frame[19] [1]), .O(n22));
    defparam i6_4_lut_adj_986.LUT_INIT = 16'hebbe;
    SB_LUT4 i2_3_lut_adj_987 (.I0(\data_in_frame[8] [4]), .I1(\data_in_frame[6] [3]), 
            .I2(Kp_23__N_934), .I3(GND_net), .O(n36099));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_987.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_988 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[7] [1]), 
            .I2(\data_in_frame[5] [0]), .I3(GND_net), .O(n36084));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_988.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_adj_989 (.I0(n35798), .I1(n4_adj_4069), .I2(GND_net), 
            .I3(GND_net), .O(n20979));   // verilog/coms.v(73[16:42])
    defparam i2_2_lut_adj_989.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_990 (.I0(\data_in_frame[21] [3]), .I1(n36772), 
            .I2(n8_adj_4046), .I3(n37847), .O(n23));
    defparam i7_4_lut_adj_990.LUT_INIT = 16'hdeed;
    SB_LUT4 i2_3_lut_adj_991 (.I0(n35730), .I1(n36084), .I2(n21797), .I3(GND_net), 
            .O(n21100));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_991.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_992 (.I0(n21690), .I1(n19969), .I2(n21620), .I3(n35699), 
            .O(n10_adj_4070));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_992.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_993 (.I0(n35798), .I1(n36099), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4050));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_993.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_994 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n21690));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_994.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_995 (.I0(n21690), .I1(\data_in_frame[2] [6]), .I2(\data_in_frame[4] [7]), 
            .I3(GND_net), .O(n35730));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_995.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_996 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[3] [1]), 
            .I2(n35730), .I3(n35724), .O(n12_adj_4071));   // verilog/coms.v(85[17:70])
    defparam i5_4_lut_adj_996.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_997 (.I0(\data_in_frame[5] [2]), .I1(n12_adj_4071), 
            .I2(\data_in_frame[5] [1]), .I3(\data_in_frame[7] [3]), .O(n32987));   // verilog/coms.v(85[17:70])
    defparam i6_4_lut_adj_997.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_998 (.I0(n20881), .I1(n21436), .I2(\data_in_frame[7] [0]), 
            .I3(n35702), .O(n10_adj_4072));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_998.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_999 (.I0(n21181), .I1(n21045), .I2(\data_in_frame[0] [7]), 
            .I3(\data_in_frame[3] [3]), .O(n19152));
    defparam i3_4_lut_adj_999.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_32_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [30]), 
            .I2(GND_net), .I3(n30708), .O(n2_adj_4073)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i5_4_lut_adj_1000 (.I0(n37418), .I1(n33841), .I2(n10_adj_4044), 
            .I3(\data_in_frame[18] [1]), .O(n21_adj_4074));
    defparam i5_4_lut_adj_1000.LUT_INIT = 16'hebbe;
    SB_CARRY add_43_32 (.CI(n30708), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n30709));
    SB_LUT4 add_43_31_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [29]), 
            .I2(GND_net), .I3(n30707), .O(n2_adj_4075)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_31 (.CI(n30707), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n30708));
    SB_LUT4 add_43_7_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n30683), .O(n35184)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1001 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n35647));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1001.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_30_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [28]), 
            .I2(GND_net), .I3(n30706), .O(n2_adj_4076)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_30 (.CI(n30706), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n30707));
    SB_LUT4 add_43_29_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(n30705), .O(n34638)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_7 (.CI(n30683), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n30684));
    SB_LUT4 i1_2_lut_adj_1002 (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[19] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4077));
    defparam i1_2_lut_adj_1002.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1003 (.I0(\data_in_frame[21] [7]), .I1(n20961), 
            .I2(n21568), .I3(n6_adj_4077), .O(n37542));
    defparam i4_4_lut_adj_1003.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_6_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n30682), .O(n35248)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_6 (.CI(n30682), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n30683));
    SB_LUT4 select_400_Select_31_i3_2_lut (.I0(\FRAME_MATCHER.i [31]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4078));
    defparam select_400_Select_31_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut_adj_1004 (.I0(\data_out_frame[25] [7]), .I1(n33870), 
            .I2(n36933), .I3(n35889), .O(n10_adj_4079));
    defparam i4_4_lut_adj_1004.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1005 (.I0(n32851), .I1(\data_out_frame[25] [7]), 
            .I2(n36178), .I3(n6_adj_4080), .O(n37877));
    defparam i4_4_lut_adj_1005.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1006 (.I0(\data_out_frame[19] [2]), .I1(n33963), 
            .I2(\data_out_frame[23] [6]), .I3(GND_net), .O(n36933));
    defparam i2_3_lut_adj_1006.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1007 (.I0(n36933), .I1(\data_out_frame[24] [1]), 
            .I2(\data_out_frame[24] [0]), .I3(n6_adj_4081), .O(n36611));
    defparam i4_4_lut_adj_1007.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1008 (.I0(n33893), .I1(n32954), .I2(\data_out_frame[19] [7]), 
            .I3(n33954), .O(n36986));
    defparam i3_4_lut_adj_1008.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_5_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n30681), .O(n35246)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_1009 (.I0(n33870), .I1(n36986), .I2(\data_out_frame[23] [7]), 
            .I3(GND_net), .O(n35945));
    defparam i2_3_lut_adj_1009.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1010 (.I0(n35945), .I1(n21586), .I2(n32951), 
            .I3(n6_adj_4082), .O(n38149));
    defparam i4_4_lut_adj_1010.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1011 (.I0(\data_out_frame[19] [4]), .I1(\data_out_frame[15] [0]), 
            .I2(n35929), .I3(n35618), .O(n33870));
    defparam i3_4_lut_adj_1011.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1012 (.I0(n35929), .I1(n36278), .I2(n35975), 
            .I3(GND_net), .O(n33893));
    defparam i2_3_lut_adj_1012.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1013 (.I0(n32951), .I1(n33893), .I2(n33870), 
            .I3(GND_net), .O(n33872));
    defparam i2_3_lut_adj_1013.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1014 (.I0(n36066), .I1(n33921), .I2(n33872), 
            .I3(GND_net), .O(n32851));
    defparam i2_3_lut_adj_1014.LUT_INIT = 16'h6969;
    SB_LUT4 i2_4_lut_adj_1015 (.I0(n36831), .I1(n37310), .I2(n10_adj_4083), 
            .I3(n35923), .O(n18_adj_4084));
    defparam i2_4_lut_adj_1015.LUT_INIT = 16'hedde;
    SB_LUT4 i2_3_lut_adj_1016 (.I0(\data_out_frame[24] [3]), .I1(\data_out_frame[24] [2]), 
            .I2(n32851), .I3(GND_net), .O(n36899));
    defparam i2_3_lut_adj_1016.LUT_INIT = 16'h6969;
    SB_LUT4 i5_4_lut_adj_1017 (.I0(n33007), .I1(n36317), .I2(n36151), 
            .I3(n36268), .O(n12_adj_4085));
    defparam i5_4_lut_adj_1017.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1018 (.I0(n35926), .I1(n12_adj_4085), .I2(n36278), 
            .I3(n35690), .O(n36066));
    defparam i6_4_lut_adj_1018.LUT_INIT = 16'h6996;
    SB_CARRY add_43_29 (.CI(n30705), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n30706));
    SB_LUT4 i1_2_lut_adj_1019 (.I0(n36066), .I1(n36247), .I2(GND_net), 
            .I3(GND_net), .O(n36248));
    defparam i1_2_lut_adj_1019.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1020 (.I0(\data_out_frame[17] [4]), .I1(\data_out_frame[15] [2]), 
            .I2(\data_out_frame[15] [3]), .I3(n33815), .O(n35975));
    defparam i3_4_lut_adj_1020.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_28_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [26]), 
            .I2(GND_net), .I3(n30704), .O(n34646)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_28 (.CI(n30704), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n30705));
    SB_LUT4 add_43_27_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [25]), 
            .I2(GND_net), .I3(n30703), .O(n34650)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1021 (.I0(\data_out_frame[20] [2]), .I1(n32951), 
            .I2(GND_net), .I3(GND_net), .O(n33921));
    defparam i1_2_lut_adj_1021.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1022 (.I0(n7_adj_4086), .I1(n33928), .I2(n33921), 
            .I3(n36178), .O(n37228));
    defparam i4_4_lut_adj_1022.LUT_INIT = 16'h9669;
    SB_LUT4 i13984_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35569), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n22387));
    defparam i13984_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1023 (.I0(n32920), .I1(n21611), .I2(n36090), 
            .I3(n6_adj_4088), .O(n37246));
    defparam i4_4_lut_adj_1023.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_1024 (.I0(n37330), .I1(n38298), .I2(n13_adj_4042), 
            .I3(n14_adj_4041), .O(n26));
    defparam i10_4_lut_adj_1024.LUT_INIT = 16'hfbbf;
    SB_LUT4 i14_4_lut (.I0(n21_adj_4074), .I1(n23), .I2(n22), .I3(n24_adj_4068), 
            .O(n30_adj_4089));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1025 (.I0(n35687), .I1(n37542), .I2(n35906), 
            .I3(\data_in_frame[21] [0]), .O(n17));
    defparam i1_4_lut_adj_1025.LUT_INIT = 16'hdeed;
    SB_LUT4 i15_4_lut_adj_1026 (.I0(n17), .I1(n30_adj_4089), .I2(n26), 
            .I3(n18_adj_4084), .O(n31_adj_4090));
    defparam i15_4_lut_adj_1026.LUT_INIT = 16'hfffe;
    SB_LUT4 i13985_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35569), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n22388));
    defparam i13985_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n35118), .S(n35062));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n35158), .S(n35082));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n35156), .S(n35084));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n27009), .S(n27759));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n35154), .S(n35086));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n35200), .S(n34990));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n35186), .S(n35116));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n35152), .S(n35088));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n35150), .S(n35090));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n35148), .S(n35020));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n35146), .S(n35092));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n35144), .S(n35094));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n35142), .S(n35096));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n35140), .S(n35098));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n35138), .S(n35100));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n35136), .S(n35102));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n35134), .S(n35060));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n35132), .S(n35104));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n35130), .S(n35106));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n27007), .S(n27755));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n35128), .S(n35108));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n27005), .S(n27753));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n35126), .S(n35110));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n7_adj_4091), .S(n8_adj_4092));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n35124), .S(n35058));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n7_adj_4093), .S(n8_adj_4094));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n35122), .S(n35112));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n35120), .S(n35056));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(clk32MHz), 
            .D(n35048), .S(n35036));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1027 (.I0(n32949), .I1(n32920), .I2(GND_net), 
            .I3(GND_net), .O(n21278));
    defparam i1_2_lut_adj_1027.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1028 (.I0(\data_out_frame[18] [0]), .I1(n35881), 
            .I2(\data_out_frame[15] [5]), .I3(n21451), .O(n36151));
    defparam i3_4_lut_adj_1028.LUT_INIT = 16'h6996;
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(clk32MHz), 
            .E(n21961), .D(n35904));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_27 (.CI(n30703), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n30704));
    SB_LUT4 i1_2_lut_adj_1029 (.I0(\data_out_frame[24] [2]), .I1(\data_out_frame[24] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n35897));
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1030 (.I0(\data_out_frame[24] [5]), .I1(\data_out_frame[24] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n36087));
    defparam i1_2_lut_adj_1030.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1031 (.I0(n35840), .I1(n36151), .I2(GND_net), 
            .I3(GND_net), .O(n36272));
    defparam i1_2_lut_adj_1031.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1032 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[20] [0]), 
            .I2(\data_out_frame[17] [6]), .I3(n35878), .O(n33954));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1032.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1033 (.I0(n33954), .I1(\data_out_frame[20] [2]), 
            .I2(n35690), .I3(\data_out_frame[20] [1]), .O(n36317));
    defparam i3_4_lut_adj_1033.LUT_INIT = 16'h9669;
    SB_LUT4 i13986_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35569), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n22389));
    defparam i13986_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1034 (.I0(\data_out_frame[25] [7]), .I1(n36207), 
            .I2(n35912), .I3(n35904), .O(n21611));
    defparam i3_4_lut_adj_1034.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1035 (.I0(n35909), .I1(\data_out_frame[23] [1]), 
            .I2(n36247), .I3(n36317), .O(n32_adj_4095));
    defparam i12_4_lut_adj_1035.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1036 (.I0(n21586), .I1(n32_adj_4095), .I2(n22_adj_4096), 
            .I3(n35716), .O(n36_adj_4097));
    defparam i16_4_lut_adj_1036.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1037 (.I0(n36272), .I1(n35948), .I2(n36087), 
            .I3(n35897), .O(n34_adj_4098));
    defparam i14_4_lut_adj_1037.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1038 (.I0(\data_out_frame[23] [5]), .I1(n32964), 
            .I2(n32954), .I3(\data_out_frame[23] [7]), .O(n35_adj_4099));
    defparam i15_4_lut_adj_1038.LUT_INIT = 16'h6996;
    SB_LUT4 i13987_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35569), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n22390));
    defparam i13987_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13988_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35569), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n22391));
    defparam i13988_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_4_lut_adj_1039 (.I0(n35972), .I1(n32876), .I2(n35889), 
            .I3(\data_out_frame[24] [7]), .O(n33));
    defparam i13_4_lut_adj_1039.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut (.I0(n33), .I1(n35_adj_4099), .I2(n34_adj_4098), 
            .I3(n36_adj_4097), .O(n36090));
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13989_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35569), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n22392));
    defparam i13989_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1040 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[2] [3]), .I3(GND_net), .O(n21436));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1040.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1041 (.I0(\data_in_frame[4] [5]), .I1(n35702), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_943));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1041.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1042 (.I0(n20771), .I1(\FRAME_MATCHER.state_31__N_2565 [3]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(n17814), .O(n18082));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1042.LUT_INIT = 16'h4000;
    SB_LUT4 i18618_2_lut_3_lut (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [28]), 
            .I3(GND_net), .O(n27009));
    defparam i18618_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(clk32MHz), 
            .E(n21961), .D(n36210));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(clk32MHz), 
            .E(n21961), .D(n35912));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(clk32MHz), 
            .E(n21961), .D(n37142));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(clk32MHz), 
            .E(n21961), .D(n36207));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_4_lut_adj_1043 (.I0(\FRAME_MATCHER.state [0]), .I1(n18279), 
            .I2(n28068), .I3(n27756), .O(n13_adj_4100));
    defparam i5_4_lut_adj_1043.LUT_INIT = 16'hfffe;
    SB_LUT4 i30105_4_lut (.I0(n13_adj_4100), .I1(n11_adj_4101), .I2(n27954), 
            .I3(\FRAME_MATCHER.state [2]), .O(n21925));
    defparam i30105_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut_3_lut_adj_1044 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [29]), 
            .I3(GND_net), .O(n35156));
    defparam i1_2_lut_3_lut_adj_1044.LUT_INIT = 16'he0e0;
    SB_LUT4 mux_1315_i1_3_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n4915), .I3(GND_net), .O(n4916));
    defparam mux_1315_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(clk32MHz), 
            .E(n21961), .D(n35863));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(clk32MHz), 
            .E(n21961), .D(n32949));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(clk32MHz), 
            .E(n21961), .D(n21278));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(clk32MHz), 
            .E(n21961), .D(n37246));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(clk32MHz), 
            .E(n21961), .D(n37228));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(clk32MHz), 
            .E(n21961), .D(n36248));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(clk32MHz), 
            .E(n21961), .D(n36899));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(clk32MHz), 
            .E(n21961), .D(n38149));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(clk32MHz), 
            .E(n21961), .D(n36611));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(clk32MHz), 
            .E(n21961), .D(n37877));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(clk32MHz), 
            .E(n21961), .D(n36761));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_4058), .S(n3_adj_4078));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1045 (.I0(\data_out_frame[15] [4]), .I1(n36204), 
            .I2(n32865), .I3(GND_net), .O(n35878));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1045.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1046 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n21451));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1046.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1047 (.I0(n35871), .I1(n36148), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4102));
    defparam i1_2_lut_adj_1047.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1048 (.I0(n36801), .I1(n21451), .I2(n35878), 
            .I3(n6_adj_4102), .O(n37037));
    defparam i4_4_lut_adj_1048.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1049 (.I0(n35917), .I1(n36164), .I2(GND_net), 
            .I3(GND_net), .O(n32964));
    defparam i1_2_lut_adj_1049.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1050 (.I0(\data_out_frame[20] [2]), .I1(n37037), 
            .I2(GND_net), .I3(GND_net), .O(n35716));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1050.LUT_INIT = 16'h9999;
    SB_LUT4 i13990_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35569), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n22393));
    defparam i13990_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_26_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [24]), 
            .I2(GND_net), .I3(n30702), .O(n34660)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13991_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35569), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n22394));
    defparam i13991_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_127_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4087));   // verilog/coms.v(154[7:23])
    defparam equal_127_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 equal_118_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4103));   // verilog/coms.v(154[7:23])
    defparam equal_118_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_CARRY add_43_5 (.CI(n30681), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n30682));
    SB_LUT4 i4_4_lut_adj_1051 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[4] [3]), 
            .I2(n21436), .I3(n6_adj_4104), .O(Kp_23__N_940));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1051.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1052 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[3] [7]), 
            .I2(\data_in_frame[0] [0]), .I3(n35727), .O(n10_adj_4105));   // verilog/coms.v(70[16:69])
    defparam i4_4_lut_adj_1052.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(\data_in_frame[4] [2]), .I1(n10_adj_4105), .I2(\data_in_frame[4] [1]), 
            .I3(GND_net), .O(Kp_23__N_934));   // verilog/coms.v(70[16:69])
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1053 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n21048));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1053.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1054 (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[4] [3]), 
            .I2(\data_in_frame[2] [0]), .I3(GND_net), .O(n35684));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1054.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1055 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[2] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n35713));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1055.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1056 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35663));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1056.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1057 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[2] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n35802));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1057.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1058 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35768));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1058.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_1__7__I_0_2_lut (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_834));   // verilog/coms.v(78[16:27])
    defparam data_in_frame_1__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1059 (.I0(\data_in_frame[3] [3]), .I1(\data_in_frame[5] [4]), 
            .I2(\data_in_frame[3] [1]), .I3(n6_adj_4106), .O(n35624));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1059.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1060 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35738));
    defparam i1_2_lut_adj_1060.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1061 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[2] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35757));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1061.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1062 (.I0(n33327), .I1(n32945), .I2(\data_out_frame[25] [0]), 
            .I3(\data_out_frame[24] [6]), .O(n10_adj_4107));
    defparam i4_4_lut_adj_1062.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_4_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n30680), .O(n35244)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1063 (.I0(n32920), .I1(n35862), .I2(GND_net), 
            .I3(GND_net), .O(n35863));
    defparam i1_2_lut_adj_1063.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1064 (.I0(n35935), .I1(\data_out_frame[15] [5]), 
            .I2(\data_out_frame[17] [7]), .I3(n36115), .O(n10_adj_4108));
    defparam i4_4_lut_adj_1064.LUT_INIT = 16'h6996;
    SB_CARRY add_43_4 (.CI(n30680), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n30681));
    SB_LUT4 i5_3_lut_adj_1065 (.I0(n35871), .I1(n10_adj_4108), .I2(n36944), 
            .I3(GND_net), .O(n36801));
    defparam i5_3_lut_adj_1065.LUT_INIT = 16'h6969;
    SB_CARRY add_43_26 (.CI(n30702), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n30703));
    SB_LUT4 i3_4_lut_adj_1066 (.I0(\data_out_frame[18] [1]), .I1(n36801), 
            .I2(n36944), .I3(\data_out_frame[16] [1]), .O(n35917));
    defparam i3_4_lut_adj_1066.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_25_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [23]), 
            .I2(GND_net), .I3(n30701), .O(n34668)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_43_3_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n30679), .O(n35242)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_25 (.CI(n30701), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n30702));
    SB_LUT4 i2_3_lut_adj_1067 (.I0(n37644), .I1(n2208), .I2(\data_out_frame[23] [0]), 
            .I3(GND_net), .O(n35972));
    defparam i2_3_lut_adj_1067.LUT_INIT = 16'h6969;
    SB_CARRY add_43_3 (.CI(n30679), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n30680));
    SB_LUT4 i1_4_lut_adj_1068 (.I0(\data_out_frame[25] [1]), .I1(n32934), 
            .I2(n35972), .I3(n32942), .O(n35862));
    defparam i1_4_lut_adj_1068.LUT_INIT = 16'h9669;
    SB_LUT4 add_43_2_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n35240)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1069 (.I0(n35862), .I1(n35983), .I2(GND_net), 
            .I3(GND_net), .O(n36207));
    defparam i1_2_lut_adj_1069.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1070 (.I0(\data_out_frame[18] [3]), .I1(n35600), 
            .I2(GND_net), .I3(GND_net), .O(n36014));
    defparam i1_2_lut_adj_1070.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_24_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [22]), 
            .I2(GND_net), .I3(n30700), .O(n34672)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1071 (.I0(\data_out_frame[18] [2]), .I1(n32867), 
            .I2(n36259), .I3(n36115), .O(n36164));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_1071.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1072 (.I0(n19038), .I1(\data_out_frame[20] [4]), 
            .I2(n32876), .I3(GND_net), .O(n32945));
    defparam i2_3_lut_adj_1072.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1073 (.I0(\data_out_frame[25] [2]), .I1(n33064), 
            .I2(n32945), .I3(\data_out_frame[23] [1]), .O(n10_adj_4109));
    defparam i4_4_lut_adj_1073.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_4073), .S(n3_adj_4035));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_4075), .S(n3_adj_4033));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_4076), .S(n3_adj_4032));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n34638), .S(n3_adj_4031));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n34646), .S(n3_adj_4030));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n34650), .S(n3_adj_4029));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n34660), .S(n3_adj_4028));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n34668), .S(n3_adj_4027));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n34672), .S(n3_adj_4026));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n34684), .S(n3_adj_4025));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n34700), .S(n3_adj_4024));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1074 (.I0(\data_in_frame[5] [0]), .I1(\data_in_frame[2] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4110));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1074.LUT_INIT = 16'h6666;
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n34722), .S(n3_adj_4023));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n34746), .S(n3_adj_4022));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_24 (.CI(n30700), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n30701));
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n34766), .S(n3_adj_4021));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n34790), .S(n3_adj_4020));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n34816), .S(n3_adj_4019));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n34842), .S(n3_adj_4018));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n34866), .S(n3_adj_4017));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n34890), .S(n3_adj_4016));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n34920), .S(n3_adj_4015));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n34940), .S(n3_adj_4014));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n34962), .S(n3_adj_4013));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n34988), .S(n3_adj_4012));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n35022), .S(n3_adj_4011));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n35114), .S(n3_adj_4010));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n35184), .S(n3_adj_4009));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n35248), .S(n3_adj_4005));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n35246), .S(n3_adj_4004));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n35244), .S(n3_adj_4003));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n35242), .S(n3_adj_4002));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1075 (.I0(\data_out_frame[25] [3]), .I1(n35983), 
            .I2(n33979), .I3(GND_net), .O(n37142));
    defparam i2_3_lut_adj_1075.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1076 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(n33991), .I3(GND_net), .O(n36944));
    defparam i2_3_lut_adj_1076.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1077 (.I0(\data_out_frame[20] [5]), .I1(n36944), 
            .I2(n36008), .I3(n33961), .O(n35948));
    defparam i3_4_lut_adj_1077.LUT_INIT = 16'h9669;
    SB_LUT4 add_43_23_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [21]), 
            .I2(GND_net), .I3(n30699), .O(n34684)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n30679));
    SB_CARRY add_43_23 (.CI(n30699), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n30700));
    SB_LUT4 i2_3_lut_adj_1078 (.I0(\data_out_frame[23] [2]), .I1(n37273), 
            .I2(\data_out_frame[23] [1]), .I3(GND_net), .O(n33979));
    defparam i2_3_lut_adj_1078.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1079 (.I0(\data_out_frame[25] [3]), .I1(n35987), 
            .I2(n33979), .I3(GND_net), .O(n35912));
    defparam i2_3_lut_adj_1079.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1080 (.I0(\data_out_frame[23] [3]), .I1(\data_out_frame[23] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35909));
    defparam i1_2_lut_adj_1080.LUT_INIT = 16'h6666;
    SB_LUT4 add_43_22_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [20]), 
            .I2(GND_net), .I3(n30698), .O(n34700)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1081 (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[14] [1]), 
            .I2(n6_adj_4111), .I3(n35935), .O(n35600));
    defparam i1_4_lut_adj_1081.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1082 (.I0(\data_out_frame[18] [4]), .I1(n36011), 
            .I2(n35600), .I3(n32863), .O(n19038));
    defparam i3_4_lut_adj_1082.LUT_INIT = 16'h6996;
    SB_LUT4 i1418_2_lut (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n2206));   // verilog/coms.v(78[16:27])
    defparam i1418_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1083 (.I0(n2206), .I1(n19038), .I2(n33986), .I3(n6_adj_4112), 
            .O(n2208));
    defparam i4_4_lut_adj_1083.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1084 (.I0(n2208), .I1(n20475), .I2(GND_net), 
            .I3(GND_net), .O(n33015));
    defparam i1_2_lut_adj_1084.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n22407));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_4_lut_adj_1085 (.I0(\data_out_frame[25] [4]), .I1(n35909), 
            .I2(n6_adj_4113), .I3(n33939), .O(n35987));
    defparam i1_4_lut_adj_1085.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1086 (.I0(n35987), .I1(n36209), .I2(GND_net), 
            .I3(GND_net), .O(n36210));
    defparam i1_2_lut_adj_1086.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1087 (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[17] [2]), 
            .I2(n35932), .I3(n6_adj_4114), .O(n35618));   // verilog/coms.v(85[17:63])
    defparam i4_4_lut_adj_1087.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1088 (.I0(\data_out_frame[16] [7]), .I1(\data_out_frame[19] [3]), 
            .I2(n35777), .I3(n35618), .O(n10_adj_4115));
    defparam i4_4_lut_adj_1088.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1089 (.I0(\data_out_frame[15] [1]), .I1(n10_adj_4115), 
            .I2(\data_out_frame[15] [0]), .I3(GND_net), .O(n21586));
    defparam i5_3_lut_adj_1089.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1090 (.I0(\data_out_frame[8] [0]), .I1(n36051), 
            .I2(\data_out_frame[7] [6]), .I3(n20861), .O(n12_adj_4116));   // verilog/coms.v(85[17:70])
    defparam i5_4_lut_adj_1090.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1091 (.I0(\data_out_frame[5] [4]), .I1(n12_adj_4116), 
            .I2(\data_out_frame[14] [6]), .I3(n35656), .O(n35820));   // verilog/coms.v(85[17:70])
    defparam i6_4_lut_adj_1091.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1092 (.I0(n35820), .I1(n1519), .I2(\data_out_frame[12] [5]), 
            .I3(\data_out_frame[12] [4]), .O(n21789));   // verilog/coms.v(85[17:63])
    defparam i3_4_lut_adj_1092.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1093 (.I0(n35837), .I1(n21789), .I2(\data_out_frame[16] [7]), 
            .I3(n36133), .O(n10_adj_4117));
    defparam i4_4_lut_adj_1093.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1094 (.I0(\data_out_frame[18] [7]), .I1(n10_adj_4117), 
            .I2(n38156), .I3(GND_net), .O(n33986));
    defparam i5_3_lut_adj_1094.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1095 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n21015));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1095.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1096 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[15] [4]), .I3(GND_net), .O(n35881));
    defparam i2_3_lut_adj_1096.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n22406));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1097 (.I0(n36146), .I1(n35881), .I2(GND_net), 
            .I3(GND_net), .O(n32954));
    defparam i1_2_lut_adj_1097.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1098 (.I0(n32867), .I1(n35980), .I2(n33007), 
            .I3(GND_net), .O(n33991));
    defparam i2_3_lut_adj_1098.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1099 (.I0(\data_out_frame[7] [1]), .I1(n36222), 
            .I2(\data_out_frame[9] [4]), .I3(n21647), .O(n12_adj_4118));   // verilog/coms.v(71[16:62])
    defparam i5_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1100 (.I0(\data_out_frame[9] [3]), .I1(n12_adj_4118), 
            .I2(\data_out_frame[11] [5]), .I3(\data_out_frame[7] [3]), .O(n32867));   // verilog/coms.v(71[16:62])
    defparam i6_4_lut_adj_1100.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1101 (.I0(\data_out_frame[18] [0]), .I1(n33007), 
            .I2(\data_out_frame[18] [1]), .I3(\data_out_frame[17] [6]), 
            .O(n36148));
    defparam i3_4_lut_adj_1101.LUT_INIT = 16'h6996;
    SB_LUT4 i18738_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27129));
    defparam i18738_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12_4_lut_adj_1102 (.I0(\FRAME_MATCHER.state [19]), .I1(\FRAME_MATCHER.state [21]), 
            .I2(\FRAME_MATCHER.state [26]), .I3(\FRAME_MATCHER.state [28]), 
            .O(n28_adj_4119));
    defparam i12_4_lut_adj_1102.LUT_INIT = 16'hfffe;
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n22405));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n22404));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n22403));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n22402));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n22401));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n22400));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n22399));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n22398));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n22397));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n22396));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n22395));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n22394));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n22393));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n22392));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1103 (.I0(\data_out_frame[18] [5]), .I1(\data_out_frame[16] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n36011));
    defparam i1_2_lut_adj_1103.LUT_INIT = 16'h6666;
    SB_LUT4 i10_4_lut_adj_1104 (.I0(\FRAME_MATCHER.state [29]), .I1(\FRAME_MATCHER.state [31]), 
            .I2(\FRAME_MATCHER.state [16]), .I3(\FRAME_MATCHER.state [23]), 
            .O(n26_adj_4120));
    defparam i10_4_lut_adj_1104.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1105 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[15] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n36259));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1105.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_1106 (.I0(\FRAME_MATCHER.state [25]), .I1(\FRAME_MATCHER.state [30]), 
            .I2(\FRAME_MATCHER.state [17]), .I3(\FRAME_MATCHER.state [20]), 
            .O(n27_adj_4121));
    defparam i11_4_lut_adj_1106.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1107 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[16] [3]), 
            .I2(\data_out_frame[18] [4]), .I3(\data_out_frame[16] [1]), 
            .O(n36008));
    defparam i3_4_lut_adj_1107.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1108 (.I0(\data_out_frame[15] [1]), .I1(\data_out_frame[19] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n36167));
    defparam i1_2_lut_adj_1108.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut (.I0(\FRAME_MATCHER.state [27]), .I1(\FRAME_MATCHER.state [22]), 
            .I2(\FRAME_MATCHER.state [18]), .I3(\FRAME_MATCHER.state [24]), 
            .O(n25));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1109 (.I0(\data_out_frame[17] [0]), .I1(\data_out_frame[16] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n36133));
    defparam i1_2_lut_adj_1109.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1110 (.I0(\data_out_frame[15] [2]), .I1(\data_out_frame[17] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n36268));
    defparam i1_2_lut_adj_1110.LUT_INIT = 16'h6666;
    SB_LUT4 i15_4_lut_adj_1111 (.I0(n25), .I1(n27_adj_4121), .I2(n26_adj_4120), 
            .I3(n28_adj_4119), .O(n28068));
    defparam i15_4_lut_adj_1111.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1112 (.I0(\FRAME_MATCHER.state [4]), .I1(\FRAME_MATCHER.state [7]), 
            .I2(\FRAME_MATCHER.state [5]), .I3(\FRAME_MATCHER.state [6]), 
            .O(n27756));
    defparam i3_4_lut_adj_1112.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1113 (.I0(\FRAME_MATCHER.state [9]), .I1(\FRAME_MATCHER.state [15]), 
            .I2(\FRAME_MATCHER.state [11]), .I3(\FRAME_MATCHER.state [13]), 
            .O(n10_adj_4122));
    defparam i4_4_lut_adj_1113.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_2_lut (.I0(\FRAME_MATCHER.state [14]), .I1(\FRAME_MATCHER.state [8]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4123));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1114 (.I0(\FRAME_MATCHER.state [12]), .I1(n9_adj_4123), 
            .I2(\FRAME_MATCHER.state [10]), .I3(n10_adj_4122), .O(n27954));
    defparam i1_4_lut_adj_1114.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1115 (.I0(\data_out_frame[10] [7]), .I1(n36256), 
            .I2(n35615), .I3(n36034), .O(n12_adj_4124));
    defparam i5_4_lut_adj_1115.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1116 (.I0(\data_out_frame[4] [6]), .I1(n12_adj_4124), 
            .I2(\data_out_frame[13] [3]), .I3(n36109), .O(n35871));
    defparam i6_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1117 (.I0(n27954), .I1(n27756), .I2(n28068), 
            .I3(GND_net), .O(n20771));
    defparam i2_3_lut_adj_1117.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1118 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[4] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n35615));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1118.LUT_INIT = 16'h6666;
    SB_CARRY add_43_22 (.CI(n30698), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n30699));
    SB_LUT4 i1_2_lut_adj_1119 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4125));
    defparam i1_2_lut_adj_1119.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1120 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n20703));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_adj_1120.LUT_INIT = 16'hbbbb;
    SB_LUT4 i5_3_lut_adj_1121 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[13] [5]), 
            .I2(n35771), .I3(GND_net), .O(n14_adj_4126));   // verilog/coms.v(71[16:69])
    defparam i5_3_lut_adj_1121.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1122 (.I0(n21032), .I1(n1168), .I2(\data_out_frame[11] [3]), 
            .I3(n21647), .O(n15_adj_4127));   // verilog/coms.v(71[16:69])
    defparam i6_4_lut_adj_1122.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1123 (.I0(n15_adj_4127), .I1(n4_adj_4128), .I2(n14_adj_4126), 
            .I3(n4_adj_4125), .O(n33007));   // verilog/coms.v(71[16:69])
    defparam i8_4_lut_adj_1123.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1124 (.I0(n35745), .I1(\data_out_frame[12] [7]), 
            .I2(n35612), .I3(n36228), .O(n14_adj_4129));   // verilog/coms.v(73[16:42])
    defparam i6_4_lut_adj_1124.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1125 (.I0(n9_adj_4130), .I1(n14_adj_4129), .I2(\data_out_frame[8] [3]), 
            .I3(n21812), .O(n33493));   // verilog/coms.v(73[16:42])
    defparam i7_4_lut_adj_1125.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1126 (.I0(\data_out_frame[11] [2]), .I1(n21812), 
            .I2(\data_out_frame[7] [0]), .I3(GND_net), .O(n36109));
    defparam i2_3_lut_adj_1126.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1127 (.I0(n36212), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[4] [4]), .I3(\data_out_frame[5] [1]), .O(n14_adj_4131));   // verilog/coms.v(76[16:27])
    defparam i6_4_lut_adj_1127.LUT_INIT = 16'h6996;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(153[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i26392_2_lut (.I0(n20704), .I1(n20792), .I2(GND_net), .I3(GND_net), 
            .O(n36406));
    defparam i26392_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i7_4_lut_adj_1128 (.I0(\data_out_frame[11] [4]), .I1(n14_adj_4131), 
            .I2(n10_adj_4132), .I3(\data_out_frame[5] [0]), .O(n21032));   // verilog/coms.v(76[16:27])
    defparam i7_4_lut_adj_1128.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1129 (.I0(n35771), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[13] [4]), .I3(n36109), .O(n10_adj_4133));
    defparam i4_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1130 (.I0(n33493), .I1(\data_out_frame[13] [1]), 
            .I2(n33007), .I3(GND_net), .O(n35840));
    defparam i2_3_lut_adj_1130.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1131 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n36027));
    defparam i1_2_lut_adj_1131.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1132 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n36238));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1132.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1133 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n36034));
    defparam i1_2_lut_adj_1133.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1134 (.I0(\data_out_frame[8] [6]), .I1(n35638), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4134));   // verilog/coms.v(74[16:43])
    defparam i2_2_lut_adj_1134.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1135 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[9] [0]), 
            .I2(n36034), .I3(\data_out_frame[11] [0]), .O(n14_adj_4135));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1136 (.I0(\data_out_frame[13] [2]), .I1(n14_adj_4135), 
            .I2(n10_adj_4134), .I3(n36105), .O(n36204));   // verilog/coms.v(74[16:43])
    defparam i7_4_lut_adj_1136.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1137 (.I0(\data_out_frame[10] [3]), .I1(n36238), 
            .I2(n36044), .I3(n20824), .O(n20_adj_4136));   // verilog/coms.v(75[16:43])
    defparam i8_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1138 (.I0(\data_out_frame[13] [0]), .I1(n36302), 
            .I2(\data_out_frame[4] [1]), .I3(n32930), .O(n19_adj_4137));   // verilog/coms.v(75[16:43])
    defparam i7_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1139 (.I0(\data_out_frame[12] [6]), .I1(n20861), 
            .I2(n35650), .I3(n21026), .O(n21_adj_4138));   // verilog/coms.v(75[16:43])
    defparam i9_4_lut_adj_1139.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1140 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[4] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4139));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1140.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1141 (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[8] [5]), 
            .I2(\data_out_frame[8] [4]), .I3(n6_adj_4139), .O(n35638));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1141.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1142 (.I0(n21026), .I1(n21227), .I2(GND_net), 
            .I3(GND_net), .O(n36124));
    defparam i1_2_lut_adj_1142.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1143 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[11] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35629));
    defparam i1_2_lut_adj_1143.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1144 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n36096));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_1144.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1145 (.I0(n20804), .I1(n36030), .I2(GND_net), 
            .I3(GND_net), .O(n36228));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1145.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_1146 (.I0(n36096), .I1(\data_out_frame[10] [0]), 
            .I2(\data_out_frame[11] [2]), .I3(n33839), .O(n26_adj_4140));
    defparam i11_4_lut_adj_1146.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1147 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[11] [3]), 
            .I2(\data_out_frame[12] [2]), .I3(\data_out_frame[11] [5]), 
            .O(n24_adj_4141));
    defparam i9_4_lut_adj_1147.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1148 (.I0(n36174), .I1(\data_out_frame[11] [4]), 
            .I2(\data_out_frame[11] [1]), .I3(n36228), .O(n25_adj_4142));
    defparam i10_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_21_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [19]), 
            .I2(GND_net), .I3(n30697), .O(n34722)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i14_4_lut_adj_1149 (.I0(n23_adj_4143), .I1(n25_adj_4142), .I2(n24_adj_4141), 
            .I3(n26_adj_4140), .O(n37842));
    defparam i14_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1150 (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[14] [4]), 
            .I2(\data_out_frame[5] [5]), .I3(n35827), .O(n44));
    defparam i16_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1151 (.I0(n35681), .I1(\data_out_frame[14] [3]), 
            .I2(\data_out_frame[14] [7]), .I3(n36124), .O(n43));
    defparam i15_4_lut_adj_1151.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(n33815), .I1(\data_out_frame[10] [2]), .I2(n35612), 
            .I3(n35638), .O(n49));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(n36027), .I1(n36238), .I2(n35840), .I3(n35785), 
            .O(n48));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n22391));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i18_4_lut (.I0(\data_out_frame[12] [5]), .I1(n36296), .I2(n35871), 
            .I3(n35656), .O(n46));
    defparam i18_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n22390));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n22389));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n22388));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n22387));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n22386));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n22385));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i19_4_lut_adj_1152 (.I0(n37842), .I1(n35795), .I2(n36112), 
            .I3(\data_out_frame[8] [1]), .O(n47));
    defparam i19_4_lut_adj_1152.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1153 (.I0(n35629), .I1(\data_out_frame[14] [6]), 
            .I2(n32867), .I3(n33991), .O(n45));
    defparam i17_4_lut_adj_1153.LUT_INIT = 16'h9669;
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47), .I2(n46), .I3(n48), .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i25_3_lut (.I0(n49), .I1(n43), .I2(n44), .I3(GND_net), .O(n53));
    defparam i25_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i16_4_lut_adj_1154 (.I0(n36268), .I1(n36133), .I2(n36167), 
            .I3(n36008), .O(n40));
    defparam i16_4_lut_adj_1154.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1155 (.I0(\data_out_frame[16] [0]), .I1(n36259), 
            .I2(n36146), .I3(n36011), .O(n38));
    defparam i14_4_lut_adj_1155.LUT_INIT = 16'h9669;
    SB_LUT4 i15_4_lut_adj_1156 (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[19] [1]), 
            .I2(\data_out_frame[17] [7]), .I3(\data_out_frame[19] [4]), 
            .O(n39));
    defparam i15_4_lut_adj_1156.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n22384));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13_4_lut_adj_1157 (.I0(n35659), .I1(\data_out_frame[19] [2]), 
            .I2(\data_out_frame[19] [3]), .I3(n36148), .O(n37));
    defparam i13_4_lut_adj_1157.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1158 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[4] [6]), 
            .I2(\data_in_frame[5] [1]), .I3(n6_adj_4110), .O(n35699));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_1158.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1159 (.I0(\data_out_frame[15] [5]), .I1(\data_out_frame[18] [2]), 
            .I2(n53), .I3(n54), .O(n35_adj_4144));
    defparam i11_4_lut_adj_1159.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1160 (.I0(n36057), .I1(n36072), .I2(\data_in_frame[4] [7]), 
            .I3(\data_in_frame[0] [7]), .O(n10_adj_4145));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1160.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut (.I0(n37), .I1(n39), .I2(n38), .I3(n40), .O(n46_adj_4146));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1161 (.I0(\data_out_frame[17] [4]), .I1(\data_out_frame[17] [2]), 
            .I2(n21015), .I3(n33886), .O(n41));
    defparam i17_4_lut_adj_1161.LUT_INIT = 16'h9669;
    SB_LUT4 i23_4_lut (.I0(n41), .I1(n46_adj_4146), .I2(n35_adj_4144), 
            .I3(n36_adj_4147), .O(n21333));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1162 (.I0(n32867), .I1(n36197), .I2(n36027), 
            .I3(n6_adj_4148), .O(n33813));
    defparam i4_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1163 (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[14] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n35827));
    defparam i1_2_lut_adj_1163.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1164 (.I0(n34025), .I1(n35827), .I2(n33813), 
            .I3(GND_net), .O(n33961));
    defparam i2_3_lut_adj_1164.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1165 (.I0(\data_out_frame[17] [1]), .I1(\data_out_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4149));
    defparam i1_2_lut_adj_1165.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1166 (.I0(n4_adj_4149), .I1(n33961), .I2(\data_out_frame[16] [3]), 
            .I3(n35659), .O(n16_adj_4150));
    defparam i7_4_lut_adj_1166.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n22383));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n22382));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n22381));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i8_4_lut_adj_1167 (.I0(n36093), .I1(n16_adj_4150), .I2(n12_adj_4151), 
            .I3(\data_out_frame[16] [7]), .O(n32934));
    defparam i8_4_lut_adj_1167.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1168 (.I0(\data_out_frame[20] [7]), .I1(n33986), 
            .I2(n33963), .I3(n21333), .O(n20475));
    defparam i3_4_lut_adj_1168.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1169 (.I0(n20475), .I1(n32934), .I2(GND_net), 
            .I3(GND_net), .O(n33064));
    defparam i1_2_lut_adj_1169.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1170 (.I0(\data_out_frame[19] [1]), .I1(n33986), 
            .I2(GND_net), .I3(GND_net), .O(n21249));
    defparam i1_2_lut_adj_1170.LUT_INIT = 16'h9999;
    SB_LUT4 i9_4_lut_adj_1171 (.I0(n35699), .I1(n35757), .I2(n35738), 
            .I3(n35624), .O(n22_adj_4152));   // verilog/coms.v(78[16:27])
    defparam i9_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1172 (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n36296));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1172.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1173 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n36051));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1173.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1174 (.I0(n36194), .I1(n36051), .I2(\data_out_frame[14] [5]), 
            .I3(n36231), .O(n12_adj_4153));   // verilog/coms.v(74[16:27])
    defparam i5_4_lut_adj_1174.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1175 (.I0(n36017), .I1(n12_adj_4153), .I2(n36296), 
            .I3(n36024), .O(n21420));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1176 (.I0(\data_out_frame[9] [4]), .I1(n21216), 
            .I2(\data_out_frame[5] [1]), .I3(n6_adj_4154), .O(n21227));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_1176.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1177 (.I0(\FRAME_MATCHER.state [2]), .I1(n20789), 
            .I2(GND_net), .I3(GND_net), .O(n35539));
    defparam i1_2_lut_adj_1177.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_1178 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35533));
    defparam i1_2_lut_adj_1178.LUT_INIT = 16'h2222;
    SB_LUT4 i29474_3_lut (.I0(n35533), .I1(n35539), .I2(n20771), .I3(GND_net), 
            .O(n39281));
    defparam i29474_3_lut.LUT_INIT = 16'hcece;
    SB_LUT4 i2_4_lut_adj_1179 (.I0(n39281), .I1(n38292), .I2(n36420), 
            .I3(\FRAME_MATCHER.state [3]), .O(n36850));
    defparam i2_4_lut_adj_1179.LUT_INIT = 16'h3fbb;
    SB_LUT4 i2_2_lut_adj_1180 (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6));
    defparam i2_2_lut_adj_1180.LUT_INIT = 16'heeee;
    SB_LUT4 i18_4_lut_adj_1181 (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44_adj_4155));   // verilog/coms.v(154[7:23])
    defparam i18_4_lut_adj_1181.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1182 (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42_adj_4156));   // verilog/coms.v(154[7:23])
    defparam i16_4_lut_adj_1182.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1183 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43_adj_4157));   // verilog/coms.v(154[7:23])
    defparam i17_4_lut_adj_1183.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1184 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41_adj_4158));   // verilog/coms.v(154[7:23])
    defparam i15_4_lut_adj_1184.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1185 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40_adj_4159));   // verilog/coms.v(154[7:23])
    defparam i14_4_lut_adj_1185.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4160));   // verilog/coms.v(154[7:23])
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41_adj_4158), .I1(n43_adj_4157), .I2(n42_adj_4156), 
            .I3(n44_adj_4155), .O(n50));   // verilog/coms.v(154[7:23])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1186 (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45_adj_4161));   // verilog/coms.v(154[7:23])
    defparam i19_4_lut_adj_1186.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1187 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[11] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n36197));
    defparam i1_2_lut_adj_1187.LUT_INIT = 16'h6666;
    SB_CARRY add_43_21 (.CI(n30697), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n30698));
    SB_LUT4 add_43_20_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [18]), 
            .I2(GND_net), .I3(n30696), .O(n34746)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i25_4_lut (.I0(n45_adj_4161), .I1(n50), .I2(n39_adj_4160), 
            .I3(n40_adj_4159), .O(n20713));   // verilog/coms.v(154[7:23])
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1188 (.I0(n27129), .I1(n20713), .I2(\FRAME_MATCHER.i [4]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n20715));
    defparam i1_4_lut_adj_1188.LUT_INIT = 16'hfcec;
    SB_LUT4 i7_4_lut_adj_1189 (.I0(\data_in[2] [6]), .I1(\data_in[1] [2]), 
            .I2(n20768), .I3(\data_in[3] [2]), .O(n18_adj_4162));
    defparam i7_4_lut_adj_1189.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1190 (.I0(\data_in[1] [6]), .I1(n18_adj_4162), 
            .I2(\data_in[1] [3]), .I3(\data_in[2] [0]), .O(n20_adj_4163));
    defparam i9_4_lut_adj_1190.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut (.I0(\data_in[2] [5]), .I1(\data_in[0] [1]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4164));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1191 (.I0(n15_adj_4164), .I1(n20_adj_4163), .I2(\data_in[0] [5]), 
            .I3(\data_in[3] [7]), .O(n20620));
    defparam i10_4_lut_adj_1191.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_2_lut_adj_1192 (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4165));
    defparam i2_2_lut_adj_1192.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1193 (.I0(\data_in[0] [2]), .I1(\data_in[3] [5]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_4166));
    defparam i6_4_lut_adj_1193.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_1194 (.I0(\data_in[3] [6]), .I1(n14_adj_4166), 
            .I2(n10_adj_4165), .I3(\data_in[2] [1]), .O(n20762));
    defparam i7_4_lut_adj_1194.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_4_lut_adj_1195 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_4167));
    defparam i4_4_lut_adj_1195.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1196 (.I0(\data_in[3] [4]), .I1(n10_adj_4167), 
            .I2(\data_in[2] [7]), .I3(GND_net), .O(n20768));
    defparam i5_3_lut_adj_1196.LUT_INIT = 16'hdfdf;
    SB_LUT4 i28313_4_lut (.I0(\data_in[1] [5]), .I1(\data_in[1] [0]), .I2(\data_in[2] [2]), 
            .I3(\data_in[0] [3]), .O(n38341));
    defparam i28313_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_1197 (.I0(\data_in[2] [4]), .I1(\data_in[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4168));
    defparam i1_2_lut_adj_1197.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_1198 (.I0(n9_adj_4168), .I1(n38341), .I2(\data_in[3] [0]), 
            .I3(\data_in[0] [6]), .O(n20710));
    defparam i7_4_lut_adj_1198.LUT_INIT = 16'hffbf;
    SB_LUT4 i6_4_lut_adj_1199 (.I0(\data_in[0] [6]), .I1(\data_in[3] [0]), 
            .I2(\data_in[1] [4]), .I3(\data_in[1] [5]), .O(n16_adj_4169));
    defparam i6_4_lut_adj_1199.LUT_INIT = 16'hffdf;
    SB_LUT4 i7_4_lut_adj_1200 (.I0(\data_in[2] [2]), .I1(n20620), .I2(n20762), 
            .I3(\data_in[1] [0]), .O(n17_adj_4170));
    defparam i7_4_lut_adj_1200.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1201 (.I0(n17_adj_4170), .I1(\data_in[0] [3]), 
            .I2(n16_adj_4169), .I3(\data_in[2] [4]), .O(n63));
    defparam i9_4_lut_adj_1201.LUT_INIT = 16'hfeff;
    SB_LUT4 i3_4_lut_adj_1202 (.I0(\data_in[3] [3]), .I1(\data_in[2] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[3] [5]), .O(n37965));
    defparam i3_4_lut_adj_1202.LUT_INIT = 16'h8000;
    SB_LUT4 i5_4_lut_adj_1203 (.I0(\data_in[0] [7]), .I1(n20710), .I2(\data_in[3] [6]), 
            .I3(n37965), .O(n12_adj_4171));
    defparam i5_4_lut_adj_1203.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut_adj_1204 (.I0(\data_in[0] [2]), .I1(n12_adj_4171), 
            .I2(n20620), .I3(\data_in[2] [1]), .O(n63_adj_4045));
    defparam i6_4_lut_adj_1204.LUT_INIT = 16'hfdff;
    SB_LUT4 i3_4_lut_adj_1205 (.I0(\data_in[0] [5]), .I1(\data_in[1] [2]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [1]), .O(n37935));
    defparam i3_4_lut_adj_1205.LUT_INIT = 16'h8000;
    SB_LUT4 i6_4_lut_adj_1206 (.I0(\data_in[2] [5]), .I1(n20710), .I2(\data_in[1] [6]), 
            .I3(\data_in[3] [7]), .O(n16_adj_4172));
    defparam i6_4_lut_adj_1206.LUT_INIT = 16'hfffd;
    SB_LUT4 i7_4_lut_adj_1207 (.I0(n20768), .I1(n20762), .I2(\data_in[2] [6]), 
            .I3(n37935), .O(n17_adj_4173));
    defparam i7_4_lut_adj_1207.LUT_INIT = 16'hfeff;
    SB_LUT4 i9_4_lut_adj_1208 (.I0(n17_adj_4173), .I1(\data_in[2] [0]), 
            .I2(n16_adj_4172), .I3(\data_in[1] [3]), .O(n63_adj_4174));
    defparam i9_4_lut_adj_1208.LUT_INIT = 16'hfbff;
    SB_LUT4 i18852_2_lut (.I0(\FRAME_MATCHER.state [0]), .I1(n17985), .I2(GND_net), 
            .I3(GND_net), .O(\FRAME_MATCHER.state_31__N_2501 [0]));
    defparam i18852_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i3297_2_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(GND_net), .I3(GND_net), .O(n4_c));
    defparam i3297_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1209 (.I0(\FRAME_MATCHER.i [4]), .I1(n20713), .I2(GND_net), 
            .I3(GND_net), .O(n20617));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_adj_1209.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1210 (.I0(n20792), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.i [31]), .I3(n20619), .O(n26_adj_4175));
    defparam i1_4_lut_adj_1210.LUT_INIT = 16'h5054;
    SB_LUT4 i4_4_lut_adj_1211 (.I0(n20617), .I1(n4_c), .I2(n20792), .I3(\FRAME_MATCHER.state_31__N_2501 [0]), 
            .O(n10_adj_4176));
    defparam i4_4_lut_adj_1211.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1212 (.I0(n26_adj_4175), .I1(n20704), .I2(\FRAME_MATCHER.i [31]), 
            .I3(n20715), .O(n31_adj_4177));
    defparam i1_4_lut_adj_1212.LUT_INIT = 16'hbabb;
    SB_LUT4 i1_4_lut_adj_1213 (.I0(n20789), .I1(n6), .I2(\FRAME_MATCHER.state [3]), 
            .I3(n10_adj_4176), .O(n22_adj_4178));
    defparam i1_4_lut_adj_1213.LUT_INIT = 16'h7350;
    SB_LUT4 i1_2_lut_adj_1214 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35990));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1214.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1215 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state_31__N_2501 [0]), 
            .I2(n22_adj_4178), .I3(n31_adj_4177), .O(n35160));
    defparam i1_4_lut_adj_1215.LUT_INIT = 16'hdc50;
    SB_LUT4 i1_2_lut_adj_1216 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n36225));   // verilog/coms.v(71[16:62])
    defparam i1_2_lut_adj_1216.LUT_INIT = 16'h6666;
    SB_CARRY add_43_20 (.CI(n30696), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n30697));
    SB_LUT4 add_43_19_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [17]), 
            .I2(GND_net), .I3(n30695), .O(n34766)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1217 (.I0(byte_transmit_counter[6]), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4179));
    defparam i1_2_lut_adj_1217.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1218 (.I0(byte_transmit_counter[4]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[1]), 
            .O(n4_adj_4180));
    defparam i1_4_lut_adj_1218.LUT_INIT = 16'ha8a0;
    SB_LUT4 i30437_4_lut (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[7]), 
            .I2(n4_adj_4180), .I3(n4_adj_4179), .O(tx_transmit_N_3354));
    defparam i30437_4_lut.LUT_INIT = 16'h0013;
    SB_LUT4 i26467_3_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n20771), .I2(n36412), 
            .I3(GND_net), .O(n36486));
    defparam i26467_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mux_876_i1_4_lut (.I0(tx_transmit_N_3354), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n28158), .I3(n8_adj_4181), .O(n3412[0]));   // verilog/coms.v(145[4] 299[11])
    defparam mux_876_i1_4_lut.LUT_INIT = 16'h0cac;
    SB_LUT4 i2_4_lut_adj_1219 (.I0(\data_in_frame[5] [6]), .I1(n35844), 
            .I2(n10_adj_4145), .I3(\data_in_frame[5] [2]), .O(n15_adj_4182));   // verilog/coms.v(78[16:27])
    defparam i2_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 i13976_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35569), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n22379));
    defparam i13976_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_19 (.CI(n30695), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n30696));
    SB_LUT4 add_43_18_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [16]), 
            .I2(GND_net), .I3(n30694), .O(n34790)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1220 (.I0(\data_out_frame[9] [2]), .I1(\data_out_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n36212));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1220.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1221 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[8] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n35650));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1221.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1222 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35754));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1222.LUT_INIT = 16'h6666;
    SB_CARRY add_43_18 (.CI(n30694), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n30695));
    SB_LUT4 add_43_17_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [15]), 
            .I2(GND_net), .I3(n30693), .O(n34816)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_1223 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[4] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4128));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1223.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1224 (.I0(\data_out_frame[9] [4]), .I1(\data_out_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4183));   // verilog/coms.v(71[16:62])
    defparam i1_2_lut_adj_1224.LUT_INIT = 16'h6666;
    SB_LUT4 i18649_2_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n27040));
    defparam i18649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i26406_2_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n20789), .I2(GND_net), 
            .I3(GND_net), .O(n36420));
    defparam i26406_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_1225 (.I0(n36105), .I1(n35780), .I2(n20804), 
            .I3(\data_out_frame[4] [7]), .O(n18_adj_4184));
    defparam i7_4_lut_adj_1225.LUT_INIT = 16'h6996;
    SB_LUT4 i18612_2_lut (.I0(tx_active), .I1(r_SM_Main_2__N_3457[0]), .I2(GND_net), 
            .I3(GND_net), .O(n27000));
    defparam i18612_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_1226 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n20789), .I3(GND_net), .O(n35));
    defparam i2_3_lut_adj_1226.LUT_INIT = 16'hfbfb;
    SB_LUT4 i9_4_lut_adj_1227 (.I0(\data_out_frame[6] [5]), .I1(n18_adj_4184), 
            .I2(\data_out_frame[8] [5]), .I3(\data_out_frame[4] [6]), .O(n20_adj_4185));
    defparam i9_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1228 (.I0(n36241), .I1(n20_adj_4185), .I2(n16_adj_4186), 
            .I3(n36044), .O(n37915));
    defparam i10_4_lut_adj_1228.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1229 (.I0(n35754), .I1(\data_out_frame[8] [4]), 
            .I2(n35650), .I3(n18_adj_4183), .O(n30_adj_4187));   // verilog/coms.v(71[16:62])
    defparam i13_4_lut_adj_1229.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1230 (.I0(n35678), .I1(n36225), .I2(\data_out_frame[9] [5]), 
            .I3(\data_out_frame[7] [3]), .O(n28_adj_4188));   // verilog/coms.v(71[16:62])
    defparam i11_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1231 (.I0(n35990), .I1(n37915), .I2(\data_out_frame[8] [6]), 
            .I3(n36020), .O(n29_adj_4189));   // verilog/coms.v(71[16:62])
    defparam i12_4_lut_adj_1231.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1232 (.I0(n36212), .I1(n36256), .I2(\data_out_frame[9] [0]), 
            .I3(n36024), .O(n27_adj_4190));   // verilog/coms.v(71[16:62])
    defparam i10_4_lut_adj_1232.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1233 (.I0(n27_adj_4190), .I1(n29_adj_4189), .I2(n28_adj_4188), 
            .I3(n30_adj_4187), .O(n33839));   // verilog/coms.v(71[16:62])
    defparam i16_4_lut_adj_1233.LUT_INIT = 16'h6996;
    SB_LUT4 i13977_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35569), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n22380));
    defparam i13977_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1234 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[10] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n20824));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1234.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1235 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[12] [1]), .I3(GND_net), .O(n36191));
    defparam i2_3_lut_adj_1235.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1236 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35780));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1236.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1237 (.I0(n36112), .I1(\data_out_frame[8] [5]), 
            .I2(\data_out_frame[4] [1]), .I3(GND_net), .O(n21522));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1237.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1238 (.I0(\data_out_frame[10] [2]), .I1(n36305), 
            .I2(\data_out_frame[10] [1]), .I3(\data_out_frame[10] [6]), 
            .O(n35745));   // verilog/coms.v(85[17:63])
    defparam i3_4_lut_adj_1238.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1239 (.I0(n35745), .I1(n21522), .I2(\data_out_frame[10] [7]), 
            .I3(GND_net), .O(n36174));   // verilog/coms.v(85[17:63])
    defparam i2_3_lut_adj_1239.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1240 (.I0(\data_out_frame[5] [5]), .I1(n32930), 
            .I2(\data_out_frame[9] [7]), .I3(n6_adj_4191), .O(n35964));
    defparam i4_4_lut_adj_1240.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1241 (.I0(n36191), .I1(n20824), .I2(\data_out_frame[7] [5]), 
            .I3(\data_out_frame[14] [3]), .O(n16_adj_4192));
    defparam i6_4_lut_adj_1241.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1242 (.I0(n35961), .I1(n35754), .I2(\data_out_frame[8] [0]), 
            .I3(n36197), .O(n17_adj_4193));
    defparam i7_4_lut_adj_1242.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1243 (.I0(n17_adj_4193), .I1(\data_out_frame[5] [3]), 
            .I2(n16_adj_4192), .I3(n35964), .O(n38156));
    defparam i9_4_lut_adj_1243.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1244 (.I0(n36191), .I1(n36287), .I2(n21227), 
            .I3(\data_out_frame[11] [6]), .O(n10_adj_4194));
    defparam i4_4_lut_adj_1244.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1245 (.I0(n35964), .I1(n10_adj_4194), .I2(\data_out_frame[12] [0]), 
            .I3(GND_net), .O(n34025));
    defparam i5_3_lut_adj_1245.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1246 (.I0(n20912), .I1(n21420), .I2(GND_net), 
            .I3(GND_net), .O(n35837));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1246.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1247 (.I0(n34025), .I1(\data_out_frame[14] [2]), 
            .I2(n38156), .I3(GND_net), .O(n32863));
    defparam i2_3_lut_adj_1247.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n40897), .I2(n39278), .I3(byte_transmit_counter[4]), .O(n40924));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n40924_bdd_4_lut (.I0(n40924), .I1(n14_adj_4195), .I2(n7_adj_4196), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n40924_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n38348), .I2(n38349), .I3(byte_transmit_counter[2]), .O(n40918));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n40918_bdd_4_lut (.I0(n40918), .I1(n38358), .I2(n38357), .I3(byte_transmit_counter[2]), 
            .O(n14_adj_4197));
    defparam n40918_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n40912));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n40912_bdd_4_lut (.I0(n40912), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n40915));
    defparam n40912_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30837 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n40906));
    defparam byte_transmit_counter_0__bdd_4_lut_30837.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_adj_1248 (.I0(\data_out_frame[18] [7]), .I1(\data_out_frame[18] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(GND_net), .O(n35659));
    defparam i2_3_lut_adj_1248.LUT_INIT = 16'h9696;
    SB_LUT4 n40906_bdd_4_lut (.I0(n40906), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n40909));
    defparam n40906_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30832 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n40900));
    defparam byte_transmit_counter_0__bdd_4_lut_30832.LUT_INIT = 16'he4aa;
    SB_LUT4 n40900_bdd_4_lut (.I0(n40900), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n40903));
    defparam n40900_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30842 (.I0(byte_transmit_counter[1]), 
            .I1(n39279), .I2(n39280), .I3(byte_transmit_counter[2]), .O(n40894));
    defparam byte_transmit_counter_1__bdd_4_lut_30842.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1249 (.I0(\data_out_frame[19] [0]), .I1(n35659), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4198));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1249.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1250 (.I0(n32863), .I1(n35837), .I2(\data_out_frame[16] [4]), 
            .I3(n6_adj_4198), .O(n33939));   // verilog/coms.v(76[16:43])
    defparam i4_4_lut_adj_1250.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_in_frame[15] [7]), .I1(n21085), 
            .I2(\data_in_frame[9] [2]), .I3(n35764), .O(n36262));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1251 (.I0(Kp_23__N_829), .I1(\data_in_frame[3] [0]), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[1] [0]), .O(n21620));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1251.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1252 (.I0(\data_out_frame[10] [4]), .I1(n36302), 
            .I2(GND_net), .I3(GND_net), .O(n35795));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1252.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1253 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[8] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n36231));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1253.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1254 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n36305));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1254.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1255 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n36241));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1255.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1256 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[4] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n36044));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1256.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1257 (.I0(\data_out_frame[19] [6]), .I1(n36146), 
            .I2(n35881), .I3(n35975), .O(n6_adj_4081));
    defparam i1_2_lut_3_lut_4_lut_adj_1257.LUT_INIT = 16'h6996;
    SB_LUT4 n40894_bdd_4_lut (.I0(n40894), .I1(n17_adj_4199), .I2(n16_adj_4200), 
            .I3(byte_transmit_counter[2]), .O(n40897));
    defparam n40894_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30827 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n40888));
    defparam byte_transmit_counter_0__bdd_4_lut_30827.LUT_INIT = 16'he4aa;
    SB_LUT4 n40888_bdd_4_lut (.I0(n40888), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n40891));
    defparam n40888_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30817 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n40882));
    defparam byte_transmit_counter_0__bdd_4_lut_30817.LUT_INIT = 16'he4aa;
    SB_LUT4 n40882_bdd_4_lut (.I0(n40882), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n40885));
    defparam n40882_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30812 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n40876));
    defparam byte_transmit_counter_0__bdd_4_lut_30812.LUT_INIT = 16'he4aa;
    SB_LUT4 n40876_bdd_4_lut (.I0(n40876), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n40879));
    defparam n40876_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30807 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter[1]), .O(n40864));
    defparam byte_transmit_counter_0__bdd_4_lut_30807.LUT_INIT = 16'he4aa;
    SB_LUT4 n40864_bdd_4_lut (.I0(n40864), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter[1]), 
            .O(n40867));
    defparam n40864_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30797 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter[1]), .O(n40858));
    defparam byte_transmit_counter_0__bdd_4_lut_30797.LUT_INIT = 16'he4aa;
    SB_LUT4 n40858_bdd_4_lut (.I0(n40858), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter[1]), 
            .O(n40861));
    defparam n40858_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1258 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [4]), 
            .I2(\data_out_frame[20] [7]), .I3(\data_out_frame[20] [6]), 
            .O(n35690));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_3_lut_4_lut_adj_1258.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30792 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter[1]), .O(n40852));
    defparam byte_transmit_counter_0__bdd_4_lut_30792.LUT_INIT = 16'he4aa;
    SB_LUT4 n40852_bdd_4_lut (.I0(n40852), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter[1]), 
            .O(n40855));
    defparam n40852_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1259 (.I0(n2208), .I1(n20475), .I2(n37273), 
            .I3(\data_out_frame[24] [7]), .O(n32942));
    defparam i1_2_lut_3_lut_4_lut_adj_1259.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30787 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n40846));
    defparam byte_transmit_counter_0__bdd_4_lut_30787.LUT_INIT = 16'he4aa;
    SB_LUT4 n40846_bdd_4_lut (.I0(n40846), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n40849));
    defparam n40846_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1260 (.I0(n36241), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[8] [1]), .I3(n36305), .O(n10_adj_4201));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1260.LUT_INIT = 16'h6996;
    SB_LUT4 i13978_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35569), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n22381));
    defparam i13978_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1261 (.I0(\data_out_frame[13] [1]), .I1(n33493), 
            .I2(\data_out_frame[15] [2]), .I3(\data_out_frame[17] [3]), 
            .O(n35929));
    defparam i1_2_lut_3_lut_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30782 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n40828));
    defparam byte_transmit_counter_0__bdd_4_lut_30782.LUT_INIT = 16'he4aa;
    SB_LUT4 n40828_bdd_4_lut (.I0(n40828), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n40831));
    defparam n40828_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30767 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n40816));
    defparam byte_transmit_counter_0__bdd_4_lut_30767.LUT_INIT = 16'he4aa;
    SB_LUT4 n40816_bdd_4_lut (.I0(n40816), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n40819));
    defparam n40816_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30757 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter[1]), .O(n40810));
    defparam byte_transmit_counter_0__bdd_4_lut_30757.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1262 (.I0(\data_out_frame[8] [3]), .I1(n35681), 
            .I2(GND_net), .I3(GND_net), .O(n1519));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_1262.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1263 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[14] [7]), .I3(n36030), .O(n10_adj_4202));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_1263.LUT_INIT = 16'h6996;
    SB_LUT4 n40810_bdd_4_lut (.I0(n40810), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter[1]), 
            .O(n40813));
    defparam n40810_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30752 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter[1]), .O(n40804));
    defparam byte_transmit_counter_0__bdd_4_lut_30752.LUT_INIT = 16'he4aa;
    SB_LUT4 n40804_bdd_4_lut (.I0(n40804), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter[1]), 
            .O(n40807));
    defparam n40804_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30747 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter[1]), .O(n40798));
    defparam byte_transmit_counter_0__bdd_4_lut_30747.LUT_INIT = 16'he4aa;
    SB_LUT4 n40798_bdd_4_lut (.I0(n40798), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter[1]), 
            .O(n40801));
    defparam n40798_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30742 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter[1]), .O(n40792));
    defparam byte_transmit_counter_0__bdd_4_lut_30742.LUT_INIT = 16'he4aa;
    SB_LUT4 n40792_bdd_4_lut (.I0(n40792), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter[1]), 
            .O(n40795));
    defparam n40792_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30737 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter[1]), .O(n40786));
    defparam byte_transmit_counter_0__bdd_4_lut_30737.LUT_INIT = 16'he4aa;
    SB_LUT4 i11_4_lut_adj_1264 (.I0(n15_adj_4182), .I1(n22_adj_4152), .I2(n36054), 
            .I3(n35802), .O(n24_adj_4203));   // verilog/coms.v(78[16:27])
    defparam i11_4_lut_adj_1264.LUT_INIT = 16'h6996;
    SB_CARRY add_43_17 (.CI(n30693), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n30694));
    SB_LUT4 i12_4_lut_adj_1265 (.I0(n35713), .I1(n24_adj_4203), .I2(n20_adj_4204), 
            .I3(n35684), .O(n33636));   // verilog/coms.v(78[16:27])
    defparam i12_4_lut_adj_1265.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_16_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [14]), 
            .I2(GND_net), .I3(n30692), .O(n34842)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 n40786_bdd_4_lut (.I0(n40786), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter[1]), 
            .O(n40789));
    defparam n40786_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_30847 (.I0(byte_transmit_counter[3]), 
            .I1(n40663), .I2(n39274), .I3(byte_transmit_counter[4]), .O(n40780));
    defparam byte_transmit_counter_3__bdd_4_lut_30847.LUT_INIT = 16'he4aa;
    SB_LUT4 n40780_bdd_4_lut (.I0(n40780), .I1(n14_adj_4205), .I2(n7_adj_4206), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n40780_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_30727 (.I0(byte_transmit_counter[3]), 
            .I1(n40669), .I2(n39263), .I3(byte_transmit_counter[4]), .O(n40774));
    defparam byte_transmit_counter_3__bdd_4_lut_30727.LUT_INIT = 16'he4aa;
    SB_LUT4 n40774_bdd_4_lut (.I0(n40774), .I1(n14_adj_4197), .I2(n7_adj_4207), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n40774_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_30722 (.I0(byte_transmit_counter[3]), 
            .I1(n40675), .I2(n39260), .I3(byte_transmit_counter[4]), .O(n40768));
    defparam byte_transmit_counter_3__bdd_4_lut_30722.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1266 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[8] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n36017));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1266.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1267 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35792));
    defparam i1_2_lut_adj_1267.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1268 (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n36194));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1268.LUT_INIT = 16'h6666;
    SB_LUT4 n40768_bdd_4_lut (.I0(n40768), .I1(n14_adj_4208), .I2(n7_adj_4209), 
            .I3(byte_transmit_counter[4]), .O(tx_data[3]));
    defparam n40768_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_30717 (.I0(byte_transmit_counter[3]), 
            .I1(n40681), .I2(n39257), .I3(byte_transmit_counter[4]), .O(n40762));
    defparam byte_transmit_counter_3__bdd_4_lut_30717.LUT_INIT = 16'he4aa;
    SB_LUT4 n40762_bdd_4_lut (.I0(n40762), .I1(n14_adj_4210), .I2(n7_adj_4211), 
            .I3(byte_transmit_counter[4]), .O(tx_data[4]));
    defparam n40762_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_30712 (.I0(byte_transmit_counter[3]), 
            .I1(n40687), .I2(n39254), .I3(byte_transmit_counter[4]), .O(n40756));
    defparam byte_transmit_counter_3__bdd_4_lut_30712.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1269 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n20861));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1269.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1270 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[12] [2]), .I3(GND_net), .O(n35961));
    defparam i2_3_lut_adj_1270.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1271 (.I0(n36194), .I1(\data_out_frame[9] [7]), 
            .I2(n35792), .I3(\data_out_frame[10] [0]), .O(n14_adj_4212));   // verilog/coms.v(74[16:27])
    defparam i6_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1272 (.I0(\data_out_frame[14] [4]), .I1(n14_adj_4212), 
            .I2(n10_adj_4213), .I3(n35678), .O(n20912));   // verilog/coms.v(74[16:27])
    defparam i7_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 n40756_bdd_4_lut (.I0(n40756), .I1(n14_adj_4214), .I2(n7_adj_4215), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n40756_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_30707 (.I0(byte_transmit_counter[3]), 
            .I1(n40693), .I2(n39251), .I3(byte_transmit_counter[4]), .O(n40750));
    defparam byte_transmit_counter_3__bdd_4_lut_30707.LUT_INIT = 16'he4aa;
    SB_LUT4 n40750_bdd_4_lut (.I0(n40750), .I1(n14_adj_4216), .I2(n7_adj_4217), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n40750_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY add_43_16 (.CI(n30692), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n30693));
    SB_LUT4 i1_2_lut_adj_1273 (.I0(n33886), .I1(n20912), .I2(GND_net), 
            .I3(GND_net), .O(n36093));
    defparam i1_2_lut_adj_1273.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1274 (.I0(n21789), .I1(\data_out_frame[16] [6]), 
            .I2(n35777), .I3(n6_adj_4218), .O(n33963));
    defparam i4_4_lut_adj_1274.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1275 (.I0(\data_out_frame[19] [2]), .I1(n33963), 
            .I2(GND_net), .I3(GND_net), .O(n21240));
    defparam i1_2_lut_adj_1275.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1276 (.I0(n33939), .I1(\data_out_frame[23] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35889));
    defparam i1_2_lut_adj_1276.LUT_INIT = 16'h9999;
    SB_LUT4 i2_3_lut_adj_1277 (.I0(Kp_23__N_937), .I1(n21048), .I2(Kp_23__N_934), 
            .I3(GND_net), .O(n35751));
    defparam i2_3_lut_adj_1277.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1278 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n35578), .O(n35579));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1278.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_4_lut_adj_1279 (.I0(\data_out_frame[25] [5]), .I1(\data_out_frame[23] [4]), 
            .I2(n6_adj_4219), .I3(n21240), .O(n36209));
    defparam i1_4_lut_adj_1279.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1280 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n35560), .O(n35562));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1280.LUT_INIT = 16'hffbf;
    SB_LUT4 add_43_15_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [13]), 
            .I2(GND_net), .I3(n30691), .O(n34866)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i28302_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n15));
    defparam i28302_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n22380));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1281 (.I0(n36209), .I1(n35889), .I2(\data_out_frame[25] [6]), 
            .I3(n21240), .O(n10_adj_4221));
    defparam i4_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1282 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n35560), .O(n35561));
    defparam i1_2_lut_3_lut_4_lut_adj_1282.LUT_INIT = 16'hff7f;
    SB_LUT4 i14096_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35578), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n22499));
    defparam i14096_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14097_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35578), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n22500));
    defparam i14097_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1283 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n35578), .O(n35586));
    defparam i1_2_lut_3_lut_4_lut_adj_1283.LUT_INIT = 16'hff7f;
    SB_CARRY add_43_15 (.CI(n30691), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n30692));
    SB_LUT4 i14098_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35578), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n22501));
    defparam i14098_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14099_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35578), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n22502));
    defparam i14099_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14100_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35578), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n22503));
    defparam i14100_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14101_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35578), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n22504));
    defparam i14101_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1284 (.I0(\FRAME_MATCHER.state [2]), .I1(n20792), 
            .I2(GND_net), .I3(GND_net), .O(n20794));   // verilog/coms.v(222[5:21])
    defparam i1_2_lut_adj_1284.LUT_INIT = 16'hdddd;
    SB_LUT4 i14102_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35578), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n22505));
    defparam i14102_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14103_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35578), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n22506));
    defparam i14103_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n38425), .I3(n38423), .O(n7_adj_4223));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_adj_1285 (.I0(\FRAME_MATCHER.state [2]), .I1(n20792), 
            .I2(GND_net), .I3(GND_net), .O(n20793));   // verilog/coms.v(151[5:27])
    defparam i1_2_lut_adj_1285.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1286 (.I0(\data_out_frame[5] [0]), .I1(n1168), 
            .I2(\data_out_frame[6] [7]), .I3(\data_out_frame[4] [5]), .O(n21647));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_4_lut_adj_1286.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1287 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [7]), 
            .I2(n35647), .I3(n6_adj_4224), .O(Kp_23__N_810));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_1287.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1288 (.I0(\data_in_frame[0] [0]), .I1(Kp_23__N_810), 
            .I2(GND_net), .I3(GND_net), .O(n35811));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_adj_1288.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n38419), .I3(n38417), .O(n7_adj_4217));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i9_4_lut_adj_1289 (.I0(n20881), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[1] [2]), .I3(n35663), .O(n26_adj_4225));
    defparam i9_4_lut_adj_1289.LUT_INIT = 16'h1040;
    SB_LUT4 i13979_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35569), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n22382));
    defparam i13979_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i10_4_lut_adj_1290 (.I0(\data_in_frame[1] [5]), .I1(n18279), 
            .I2(\data_in_frame[1] [3]), .I3(\data_in_frame[1] [6]), .O(n27_adj_4226));
    defparam i10_4_lut_adj_1290.LUT_INIT = 16'h2000;
    SB_LUT4 i13_4_lut_adj_1291 (.I0(\data_in_frame[2] [0]), .I1(n26_adj_4225), 
            .I2(n5), .I3(n35811), .O(n30_adj_4227));
    defparam i13_4_lut_adj_1291.LUT_INIT = 16'h0804;
    SB_LUT4 i6_4_lut_adj_1292 (.I0(\data_in_frame[0] [7]), .I1(Kp_23__N_810), 
            .I2(\data_in_frame[1] [1]), .I3(\data_in_frame[2] [1]), .O(n23_adj_4228));
    defparam i6_4_lut_adj_1292.LUT_INIT = 16'h2184;
    SB_LUT4 i14_4_lut_adj_1293 (.I0(n27_adj_4226), .I1(\data_in_frame[1] [4]), 
            .I2(n22_adj_4229), .I3(n21436), .O(n31_adj_4230));
    defparam i14_4_lut_adj_1293.LUT_INIT = 16'h0080;
    SB_LUT4 i16_4_lut_adj_1294 (.I0(n31_adj_4230), .I1(n23_adj_4228), .I2(n30_adj_4227), 
            .I3(n38325), .O(\FRAME_MATCHER.state_31__N_2565 [3]));
    defparam i16_4_lut_adj_1294.LUT_INIT = 16'h0080;
    SB_LUT4 i2_3_lut_adj_1295 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n20771), .I3(GND_net), .O(n20795));   // verilog/coms.v(231[5:23])
    defparam i2_3_lut_adj_1295.LUT_INIT = 16'hfefe;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n38413), .I3(n38411), .O(n7_adj_4215));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 add_43_14_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [12]), 
            .I2(GND_net), .I3(n30690), .O(n34890)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n38407), .I3(n38405), .O(n7_adj_4211));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_CARRY add_43_14 (.CI(n30690), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n30691));
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n38401), .I3(n38399), .O(n7_adj_4209));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_4_lut_adj_1296 (.I0(\FRAME_MATCHER.state [3]), .I1(n20794), 
            .I2(n4_adj_4231), .I3(n18028), .O(n6_adj_4232));   // verilog/coms.v(115[11:12])
    defparam i1_4_lut_adj_1296.LUT_INIT = 16'ha2a0;
    SB_LUT4 i1_4_lut_adj_1297 (.I0(n20795), .I1(n6_adj_4232), .I2(\FRAME_MATCHER.state_31__N_2565 [3]), 
            .I3(n20703), .O(n35036));   // verilog/coms.v(115[11:12])
    defparam i1_4_lut_adj_1297.LUT_INIT = 16'hccdc;
    SB_LUT4 i13980_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35569), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n22383));
    defparam i13980_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n38386), .I3(n38384), .O(n7_adj_4196));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 add_43_13_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [11]), 
            .I2(GND_net), .I3(n30689), .O(n34920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n38389), .I3(n38387), .O(n7_adj_4206));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i13981_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35569), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n22384));
    defparam i13981_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i18653_2_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n10));
    defparam i18653_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1298 (.I0(\FRAME_MATCHER.state [4]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35056));
    defparam i1_2_lut_adj_1298.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1299 (.I0(\FRAME_MATCHER.state [5]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35112));
    defparam i1_2_lut_adj_1299.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(byte_transmit_counter[1]), .I2(n38395), .I3(n38393), .O(n7_adj_4207));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_CARRY add_43_11 (.CI(n30687), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n30688));
    SB_LUT4 i14064_3_lut_4_lut (.I0(n8), .I1(n35560), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n22467));
    defparam i14064_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14065_3_lut_4_lut (.I0(n8), .I1(n35560), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n22468));
    defparam i14065_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14066_3_lut_4_lut (.I0(n8), .I1(n35560), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n22469));
    defparam i14066_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1300 (.I0(n33950), .I1(n35914), .I2(n36188), 
            .I3(GND_net), .O(n36189));
    defparam i1_2_lut_3_lut_adj_1300.LUT_INIT = 16'h9696;
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk32MHz), 
            .E(n21904), .D(n8825[0]), .R(n22138));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1301 (.I0(\FRAME_MATCHER.state [6]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4094));
    defparam i1_2_lut_adj_1301.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_30702 (.I0(byte_transmit_counter[3]), 
            .I1(n40711), .I2(n39248), .I3(byte_transmit_counter[4]), .O(n40744));
    defparam byte_transmit_counter_3__bdd_4_lut_30702.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1302 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[3] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n36057));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1302.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1303 (.I0(\FRAME_MATCHER.state [7]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35058));
    defparam i1_2_lut_adj_1303.LUT_INIT = 16'h8888;
    SB_LUT4 i14067_3_lut_4_lut (.I0(n8), .I1(n35560), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n22470));
    defparam i14067_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n22379));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14068_3_lut_4_lut (.I0(n8), .I1(n35560), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n22471));
    defparam i14068_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_3_lut_4_lut (.I0(n7_adj_4234), .I1(n21797), .I2(n35849), 
            .I3(n4_adj_3992), .O(n23_adj_4235));
    defparam i7_3_lut_4_lut.LUT_INIT = 16'hbeeb;
    SB_LUT4 i14069_3_lut_4_lut (.I0(n8), .I1(n35560), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n22472));
    defparam i14069_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1304 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(n36072), .I3(\data_in_frame[4] [7]), .O(n18_adj_3994));
    defparam i1_2_lut_3_lut_4_lut_adj_1304.LUT_INIT = 16'h6996;
    SB_CARRY add_43_13 (.CI(n30689), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n30690));
    SB_LUT4 i5_4_lut_adj_1305 (.I0(\data_in_frame[4] [0]), .I1(n36057), 
            .I2(\data_in_frame[1] [6]), .I3(\data_in_frame[2] [0]), .O(n12_adj_4236));   // verilog/coms.v(78[16:27])
    defparam i5_4_lut_adj_1305.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1306 (.I0(n11), .I1(\FRAME_MATCHER.state [8]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4092));
    defparam i1_2_lut_adj_1306.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n22378));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n40744_bdd_4_lut (.I0(n40744), .I1(n14_adj_4237), .I2(n7_adj_4223), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n40744_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i30281_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n22128));
    defparam i30281_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i14070_3_lut_4_lut (.I0(n8), .I1(n35560), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n22473));
    defparam i14070_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n22377));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1307 (.I0(\FRAME_MATCHER.state [9]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35110));
    defparam i1_2_lut_adj_1307.LUT_INIT = 16'h8888;
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .E(n21925), .D(n4917));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1308 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [30]), 
            .I3(GND_net), .O(n35158));
    defparam i1_2_lut_3_lut_adj_1308.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_3_lut_4_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n36850), 
            .I2(n17985), .I3(n2), .O(n35048));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'haa20;
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n22376));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i19354_2_lut (.I0(\FRAME_MATCHER.state [10]), .I1(n11), .I2(GND_net), 
            .I3(GND_net), .O(n27753));
    defparam i19354_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_4_lut_adj_1309 (.I0(n3_adj_4000), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n20792), .I3(n17948), .O(n4_adj_4231));   // verilog/coms.v(115[11:12])
    defparam i1_3_lut_4_lut_adj_1309.LUT_INIT = 16'habaa;
    SB_LUT4 i1_2_lut_adj_1310 (.I0(\FRAME_MATCHER.state [11]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35108));
    defparam i1_2_lut_adj_1310.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1311 (.I0(\data_out_frame[17] [0]), .I1(n33886), 
            .I2(n20912), .I3(GND_net), .O(n6_adj_4218));
    defparam i1_2_lut_3_lut_adj_1311.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1312 (.I0(\data_out_frame[12] [5]), .I1(n35932), 
            .I2(\data_out_frame[8] [3]), .I3(n35681), .O(n33886));
    defparam i2_3_lut_4_lut_adj_1312.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1313 (.I0(n11), .I1(\FRAME_MATCHER.state [12]), 
            .I2(GND_net), .I3(GND_net), .O(n27755));
    defparam i1_2_lut_adj_1313.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_adj_1314 (.I0(n36486), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n28158), .I3(GND_net), .O(n20723));
    defparam i1_3_lut_adj_1314.LUT_INIT = 16'haeae;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[12] [2]), .I3(n20861), .O(n10_adj_4213));   // verilog/coms.v(74[16:27])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14071_3_lut_4_lut (.I0(n8), .I1(n35560), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n22474));
    defparam i14071_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i30113_3_lut (.I0(n36412), .I1(n20771), .I2(n20723), .I3(GND_net), 
            .O(n37904));
    defparam i30113_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i14056_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35560), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n22459));
    defparam i14056_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1315 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[8] [1]), 
            .I2(\data_out_frame[8] [0]), .I3(GND_net), .O(n35678));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1315.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[8] [2]), 
            .I2(n10_adj_4202), .I3(n35795), .O(n35932));   // verilog/coms.v(72[16:27])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut_4_lut_adj_1316 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[5] [7]), .O(n20_adj_4204));   // verilog/coms.v(78[16:27])
    defparam i7_3_lut_4_lut_adj_1316.LUT_INIT = 16'h6996;
    SB_LUT4 i14057_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35560), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n22460));
    defparam i14057_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i30278_4_lut (.I0(n20723), .I1(n28158), .I2(n5_adj_4238), 
            .I3(n6_adj_4239), .O(n35502));
    defparam i30278_4_lut.LUT_INIT = 16'h1115;
    SB_LUT4 i14058_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35560), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n22461));
    defparam i14058_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14059_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35560), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n22462));
    defparam i14059_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14060_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35560), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n22463));
    defparam i14060_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14061_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35560), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n22464));
    defparam i14061_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13982_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35569), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n22385));
    defparam i13982_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14062_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35560), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n22465));
    defparam i14062_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1317 (.I0(\data_in_frame[1] [7]), .I1(n12_adj_4236), 
            .I2(\data_in_frame[6] [2]), .I3(n35671), .O(n35798));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_1317.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1318 (.I0(n35798), .I1(\data_in_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4240));
    defparam i2_2_lut_adj_1318.LUT_INIT = 16'h6666;
    SB_LUT4 i14063_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35560), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n22466));
    defparam i14063_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14048_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35560), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n22451));
    defparam i14048_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13983_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35569), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n22386));
    defparam i13983_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14049_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35560), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n22452));
    defparam i14049_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14050_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35560), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n22453));
    defparam i14050_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14051_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35560), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n22454));
    defparam i14051_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1319 (.I0(n35663), .I1(n36072), .I2(\data_in_frame[5] [4]), 
            .I3(\data_in_frame[7] [6]), .O(n35814));
    defparam i2_3_lut_4_lut_adj_1319.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1320 (.I0(n35805), .I1(Kp_23__N_777), .I2(n35751), 
            .I3(n33636), .O(n14_adj_4241));
    defparam i6_4_lut_adj_1320.LUT_INIT = 16'h6996;
    SB_LUT4 i14052_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35560), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n22455));
    defparam i14052_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14053_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35560), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n22456));
    defparam i14053_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1321 (.I0(n20789), .I1(n36406), .I2(\FRAME_MATCHER.state [2]), 
            .I3(\FRAME_MATCHER.state [3]), .O(n2841));
    defparam i1_4_lut_adj_1321.LUT_INIT = 16'hccc8;
    SB_LUT4 select_400_Select_0_i3_2_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n2841), 
            .I2(GND_net), .I3(GND_net), .O(n3));
    defparam select_400_Select_0_i3_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14054_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35560), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n22457));
    defparam i14054_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n22375));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n22374));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n22373));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n22372));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n22371));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n22370));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n22369));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n22368));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n22367));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n22366));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n22365));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n22364));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n22363));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n22362));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n22361));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n22360));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n22359));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n22358));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n22357));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n22356));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n22355));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n22354));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n22353));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n22352));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n22351));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n22350));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n22349));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n22348));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n22347));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n22346));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30732 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter[1]), .O(n40738));
    defparam byte_transmit_counter_0__bdd_4_lut_30732.LUT_INIT = 16'he4aa;
    SB_LUT4 i30108_3_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n36486), .I2(n28158), 
            .I3(GND_net), .O(n37539));
    defparam i30108_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 add_43_12_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [10]), 
            .I2(GND_net), .I3(n30688), .O(n34940)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_12 (.CI(n30688), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n30689));
    SB_LUT4 i14055_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35560), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n22458));
    defparam i14055_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_11_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [9]), 
            .I2(GND_net), .I3(n30687), .O(n34962)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n22345));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i30586_4_lut (.I0(n36486), .I1(\FRAME_MATCHER.state [3]), .I2(n4902), 
            .I3(n28158), .O(n36508));
    defparam i30586_4_lut.LUT_INIT = 16'h5011;
    SB_LUT4 i14040_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35560), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n22443));
    defparam i14040_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1322 (.I0(Kp_23__N_940), .I1(n14_adj_4241), .I2(n10_adj_4240), 
            .I3(Kp_23__N_943), .O(n38079));
    defparam i7_4_lut_adj_1322.LUT_INIT = 16'h6996;
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .E(n21925), .D(n4918));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i30120_2_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n4902));   // verilog/coms.v(145[4] 299[11])
    defparam i30120_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 mux_1315_i24_3_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n4915), .I3(GND_net), .O(n4939));
    defparam mux_1315_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1315_i23_3_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n4915), .I3(GND_net), .O(n4938));
    defparam mux_1315_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .E(n21925), .D(n4919));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .E(n21925), .D(n4920));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .E(n21925), .D(n4921));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .E(n21925), .D(n4922));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .E(n21925), .D(n4923));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .E(n21925), .D(n4924));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .E(n21925), .D(n4925));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .E(n21925), 
            .D(n4926));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .E(n21925), 
            .D(n4927));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .E(n21925), 
            .D(n4928));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .E(n21925), 
            .D(n4929));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .E(n21925), 
            .D(n4930));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .E(n21925), 
            .D(n4931));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .E(n21925), 
            .D(n4932));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .E(n21925), 
            .D(n4933));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .E(n21925), 
            .D(n4934));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .E(n21925), 
            .D(n4935));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .E(n21925), 
            .D(n4936));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .E(n21925), 
            .D(n4937));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .E(n21925), 
            .D(n4938));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .E(n21925), 
            .D(n4939));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR driver_enable_3875 (.Q(DE_c), .C(clk32MHz), .E(n36508), 
            .D(n4902), .R(n37539));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1323 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [4]), .I3(GND_net), .O(n36112));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1323.LUT_INIT = 16'h9696;
    SB_LUT4 i10_4_lut_adj_1324 (.I0(n5_adj_4050), .I1(n11_adj_4061), .I2(n21100), 
            .I3(n20979), .O(n26_adj_4242));
    defparam i10_4_lut_adj_1324.LUT_INIT = 16'hfffe;
    SB_LUT4 i14041_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35560), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n22444));
    defparam i14041_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1315_i22_3_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n4915), .I3(GND_net), .O(n4937));
    defparam mux_1315_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30261_3_lut_4_lut (.I0(n20700), .I1(n35), .I2(tx_active), 
            .I3(r_SM_Main_2__N_3457[0]), .O(n21904));
    defparam i30261_3_lut_4_lut.LUT_INIT = 16'h3337;
    SB_LUT4 i11_4_lut_adj_1325 (.I0(n21085), .I1(n38079), .I2(n32987), 
            .I3(n8_adj_4056), .O(n27_adj_4243));
    defparam i11_4_lut_adj_1325.LUT_INIT = 16'hffef;
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n22344));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14042_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35560), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n22445));
    defparam i14042_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14043_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35560), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n22446));
    defparam i14043_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n22343));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n22342));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14044_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35560), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n22447));
    defparam i14044_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n22341));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n22340));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14045_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35560), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n22448));
    defparam i14045_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFFESR LED_3874 (.Q(LED_c), .C(clk32MHz), .E(n35502), .D(n22128), 
            .R(n37904));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14046_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35560), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n22449));
    defparam i14046_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14047_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35560), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n22450));
    defparam i14047_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13_4_lut_adj_1326 (.I0(n32855), .I1(n26_adj_4242), .I2(n18_adj_4244), 
            .I3(n20900), .O(n29_adj_4245));
    defparam i13_4_lut_adj_1326.LUT_INIT = 16'hfffe;
    SB_LUT4 i14032_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35560), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n22435));
    defparam i14032_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14033_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35560), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n22436));
    defparam i14033_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14034_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35560), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n22437));
    defparam i14034_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14035_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35560), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n22438));
    defparam i14035_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15_4_lut_adj_1327 (.I0(n29_adj_4245), .I1(n27_adj_4243), .I2(n23_adj_4235), 
            .I3(n38300), .O(n31));
    defparam i15_4_lut_adj_1327.LUT_INIT = 16'hfeff;
    SB_LUT4 i14036_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35560), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n22439));
    defparam i14036_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1315_i21_3_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n4915), .I3(GND_net), .O(n4936));
    defparam mux_1315_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1315_i20_3_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n4915), .I3(GND_net), .O(n4935));
    defparam mux_1315_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1315_i19_3_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n4915), .I3(GND_net), .O(n4934));
    defparam mux_1315_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_9 (.CI(n30685), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n30686));
    SB_LUT4 i14037_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35560), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n22440));
    defparam i14037_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14038_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35560), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n22441));
    defparam i14038_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_adj_1328 (.I0(n20961), .I1(n33841), .I2(n35993), 
            .I3(GND_net), .O(n8_adj_4067));
    defparam i3_3_lut_adj_1328.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1315_i18_3_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n4915), .I3(GND_net), .O(n4933));
    defparam mux_1315_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_4_lut_adj_1329 (.I0(n21223), .I1(\data_in_frame[19] [4]), 
            .I2(\data_in_frame[21] [6]), .I3(\data_in_frame[19] [5]), .O(n38098));   // verilog/coms.v(268[9:85])
    defparam i2_4_lut_adj_1329.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1315_i17_3_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n4915), .I3(GND_net), .O(n4932));
    defparam mux_1315_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1315_i16_3_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n4915), .I3(GND_net), .O(n4931));
    defparam mux_1315_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1315_i15_3_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n4915), .I3(GND_net), .O(n4930));
    defparam mux_1315_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1315_i14_3_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n4915), .I3(GND_net), .O(n4929));
    defparam mux_1315_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14039_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35560), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n22442));
    defparam i14039_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1315_i13_3_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n4915), .I3(GND_net), .O(n4928));
    defparam mux_1315_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1315_i12_3_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n4915), .I3(GND_net), .O(n4927));
    defparam mux_1315_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n40738_bdd_4_lut (.I0(n40738), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter[1]), 
            .O(n40741));
    defparam n40738_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1315_i11_3_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n4915), .I3(GND_net), .O(n4926));
    defparam mux_1315_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1315_i10_3_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n4915), .I3(GND_net), .O(n4925));
    defparam mux_1315_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13968_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35569), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n22371));
    defparam i13968_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1315_i9_3_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n4915), .I3(GND_net), .O(n4924));
    defparam mux_1315_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1315_i8_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n4915), .I3(GND_net), .O(n4923));
    defparam mux_1315_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1315_i7_3_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n4915), .I3(GND_net), .O(n4922));
    defparam mux_1315_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1315_i6_3_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n4915), .I3(GND_net), .O(n4921));
    defparam mux_1315_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13969_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35569), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n22372));
    defparam i13969_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1315_i5_3_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n4915), .I3(GND_net), .O(n4920));
    defparam mux_1315_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1315_i4_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n4915), .I3(GND_net), .O(n4919));
    defparam mux_1315_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30693 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter[1]), .O(n40732));
    defparam byte_transmit_counter_0__bdd_4_lut_30693.LUT_INIT = 16'he4aa;
    SB_LUT4 i13970_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35569), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n22373));
    defparam i13970_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13971_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35569), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n22374));
    defparam i13971_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n40732_bdd_4_lut (.I0(n40732), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter[1]), 
            .O(n40735));
    defparam n40732_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13972_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35569), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n22375));
    defparam i13972_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13973_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35569), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n22376));
    defparam i13973_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13974_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35569), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n22377));
    defparam i13974_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13975_3_lut_4_lut (.I0(n8_adj_4222), .I1(n35569), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n22378));
    defparam i13975_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1330 (.I0(\data_in_frame[20] [3]), .I1(n36155), 
            .I2(n35886), .I3(n33841), .O(n37091));
    defparam i3_4_lut_adj_1330.LUT_INIT = 16'h9669;
    SB_LUT4 equal_125_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4222));   // verilog/coms.v(154[7:23])
    defparam equal_125_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1331 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n35569), .I3(\FRAME_MATCHER.i [0]), .O(n35575));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1331.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_3_lut_4_lut_adj_1332 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n20789), .I3(n20700), .O(n22179));   // verilog/coms.v(127[12] 300[6])
    defparam i2_3_lut_4_lut_adj_1332.LUT_INIT = 16'h0200;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1333 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n35578), .I3(\FRAME_MATCHER.i [0]), .O(n35585));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1333.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1334 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n35560), .I3(\FRAME_MATCHER.i [0]), .O(n35568));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1334.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_2_lut_3_lut_adj_1335 (.I0(n20629), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n20700));   // verilog/coms.v(212[5:16])
    defparam i1_2_lut_3_lut_adj_1335.LUT_INIT = 16'hbfbf;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[6] [6]), 
            .I2(\data_out_frame[4] [5]), .I3(GND_net), .O(n36105));   // verilog/coms.v(76[16:27])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_4_lut (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(n1_adj_4246), .I3(\FRAME_MATCHER.state [2]), .O(n5_adj_4238));   // verilog/coms.v(145[4] 299[11])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h50bb;
    SB_LUT4 i2_4_lut_4_lut (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state_31__N_2565 [3]), .I3(\FRAME_MATCHER.state [2]), 
            .O(n6_adj_4239));   // verilog/coms.v(145[4] 299[11])
    defparam i2_4_lut_4_lut.LUT_INIT = 16'haa04;
    SB_LUT4 equal_1505_i8_3_lut_4_lut (.I0(\data_in_frame[6] [5]), .I1(Kp_23__N_940), 
            .I2(\data_in_frame[8] [7]), .I3(n35696), .O(n8_adj_4056));   // verilog/coms.v(76[16:43])
    defparam equal_1505_i8_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1336 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [31]), 
            .I3(GND_net), .O(n35118));
    defparam i1_2_lut_3_lut_adj_1336.LUT_INIT = 16'he0e0;
    SB_LUT4 i4_4_lut_adj_1337 (.I0(\data_in_frame[18] [3]), .I1(n36155), 
            .I2(\data_in_frame[20] [4]), .I3(\data_in_frame[18] [2]), .O(n10_adj_4083));
    defparam i4_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1338 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n6_adj_4224));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1338.LUT_INIT = 16'h9696;
    SB_LUT4 i28298_3_lut_4_lut (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[2] [7]), .I3(n21440), .O(n38325));   // verilog/coms.v(77[16:27])
    defparam i28298_3_lut_4_lut.LUT_INIT = 16'hff96;
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n22840));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n22839));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n22838));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n22837));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n22836));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n22835));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n22834));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n22833));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n22832));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n22831));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n22830));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n22829));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n22828));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n22827));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n22826));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n22825));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n22824));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n22823));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n22822));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n22821));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n22820));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n22819));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n22818));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 mux_1315_i3_3_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n4915), .I3(GND_net), .O(n4918));
    defparam mux_1315_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_1505_i7_3_lut_4_lut (.I0(\data_in_frame[6] [5]), .I1(Kp_23__N_940), 
            .I2(n36069), .I3(\data_in_frame[8] [6]), .O(n7_adj_4234));   // verilog/coms.v(76[16:43])
    defparam equal_1505_i7_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n22783));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n22782));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_4_lut_4_lut_adj_1339 (.I0(\FRAME_MATCHER.state [3]), .I1(n36412), 
            .I2(n35533), .I3(\FRAME_MATCHER.state [2]), .O(n17814));
    defparam i1_4_lut_4_lut_adj_1339.LUT_INIT = 16'h2272;
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n22781));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n22780));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n22779));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n22778));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n22777));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n22776));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n22775));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n22774));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n22773));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n22772));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n22771));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14120_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35578), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n22523));
    defparam i14120_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n22770));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n22769));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n22768));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n22767));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n22766));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n22765));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n22764));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1340 (.I0(\FRAME_MATCHER.state [3]), .I1(n36412), 
            .I2(n20771), .I3(\FRAME_MATCHER.state [1]), .O(n21961));
    defparam i2_3_lut_4_lut_adj_1340.LUT_INIT = 16'h0002;
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n22763));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n22762));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n22761));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n22760));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_10_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [8]), 
            .I2(GND_net), .I3(n30686), .O(n34988)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n22759));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n22758));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n22757));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n22756));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n22755));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n22754));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n22753));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n22752));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n22751));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n22750));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n22749));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n22748));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n22747));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n22746));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(clk32MHz), .D(n22745));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(clk32MHz), .D(n22744));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(clk32MHz), .D(n22743));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(clk32MHz), .D(n22742));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(clk32MHz), .D(n22741));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(clk32MHz), .D(n22740));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(clk32MHz), .D(n22739));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(clk32MHz), .D(n22738));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n22737));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n22736));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n22735));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n22734));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n22733));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n22732));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n22731));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(clk32MHz), .D(n22730));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(clk32MHz), .D(n22729));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(clk32MHz), .D(n22728));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(clk32MHz), .D(n22727));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(clk32MHz), .D(n22726));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(clk32MHz), .D(n22725));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(clk32MHz), .D(n22724));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(clk32MHz), .D(n22721));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(clk32MHz), 
           .D(n22720));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk32MHz), 
           .D(n22719));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_10 (.CI(n30686), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n30687));
    SB_DFF data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(clk32MHz), 
           .D(n22718));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(clk32MHz), 
           .D(n22717));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(clk32MHz), 
           .D(n22716));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(clk32MHz), 
           .D(n22715));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(clk32MHz), 
           .D(n22714));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(clk32MHz), 
           .D(n22713));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n22712));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n22711));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk32MHz), 
           .D(n22710));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n22709));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n22708));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n22707));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n22706));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n22705));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n22704));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n22703));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n22702));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n22701));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n22700));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n22699));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n22698));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n22697));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n22696));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1341 (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[6] [2]), 
            .I2(\data_out_frame[4] [1]), .I3(\data_out_frame[6] [1]), .O(n20804));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1341.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n22695));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n22694));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n22693));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n22692));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n22691));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1342 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(n36020), .I3(GND_net), .O(n36222));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1342.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n22690));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n22689));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n22688));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n22687));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n22686));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n22685));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n22684));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n22683));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n22682));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n22681));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n22680));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n22679));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n22678));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n22677));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n22676));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n22675));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n22674));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n22673));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n22672));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n22671));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n22670));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n22669));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n22668));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n22667));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1343 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[8] [4]), .I3(\data_out_frame[10] [5]), .O(n36302));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1343.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n22666));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_3971_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n30716), .O(n8825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_9_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n22665));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n22664));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n22663));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n22662));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n22661));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_4_lut_adj_1344 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[7] [7]), .I3(n10_adj_4201), .O(n35681));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_4_lut_adj_1344.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut (.I0(n36112), .I1(\data_out_frame[8] [5]), .I2(\data_out_frame[4] [1]), 
            .I3(\data_out_frame[9] [1]), .O(n36256));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n22660));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n22659));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n22658));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_3971_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n30715), .O(n8825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_8_lut.LUT_INIT = 16'hC33C;
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n22657));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_3_lut_4_lut (.I0(\data_out_frame[10] [5]), .I1(n36174), 
            .I2(\data_out_frame[10] [0]), .I3(n21026), .O(n32930));
    defparam i1_3_lut_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n22656));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1345 (.I0(\data_out_frame[10] [5]), .I1(n36174), 
            .I2(\data_out_frame[7] [6]), .I3(GND_net), .O(n6_adj_4191));
    defparam i1_2_lut_3_lut_adj_1345.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1346 (.I0(\FRAME_MATCHER.state [3]), .I1(n35539), 
            .I2(n18279), .I3(n31_adj_4090), .O(n21865));
    defparam i3_4_lut_adj_1346.LUT_INIT = 16'h0004;
    SB_LUT4 i3_3_lut_4_lut (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(n27000), .O(n8_adj_4181));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1347 (.I0(n21026), .I1(\data_out_frame[10] [0]), 
            .I2(n32930), .I3(GND_net), .O(n35612));
    defparam i1_2_lut_3_lut_adj_1347.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1348 (.I0(\FRAME_MATCHER.state [0]), .I1(n17985), 
            .I2(n35589), .I3(GND_net), .O(n35046));
    defparam i1_2_lut_3_lut_adj_1348.LUT_INIT = 16'hb0b0;
    SB_LUT4 i1_3_lut_4_lut_adj_1349 (.I0(n8), .I1(\FRAME_MATCHER.i [4]), 
            .I2(n20713), .I3(\FRAME_MATCHER.i [3]), .O(n20619));
    defparam i1_3_lut_4_lut_adj_1349.LUT_INIT = 16'hfefc;
    SB_CARRY add_3971_8 (.CI(n30715), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n30716));
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n22339));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i28265_2_lut_4_lut (.I0(n20704), .I1(n20792), .I2(n20629), 
            .I3(n27040), .O(n38292));
    defparam i28265_2_lut_4_lut.LUT_INIT = 16'h8088;
    SB_LUT4 i5_2_lut_3_lut (.I0(\data_out_frame[5] [0]), .I1(n1168), .I2(\data_out_frame[6] [7]), 
            .I3(GND_net), .O(n16_adj_4186));   // verilog/coms.v(85[17:70])
    defparam i5_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i14121_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35578), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n22524));
    defparam i14121_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_3971_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n30714), .O(n8825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_7 (.CI(n30714), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n30715));
    SB_LUT4 i2_3_lut_4_lut_adj_1350 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[7] [3]), .I3(\data_out_frame[4] [7]), .O(n21216));   // verilog/coms.v(73[16:34])
    defparam i2_3_lut_4_lut_adj_1350.LUT_INIT = 16'h6996;
    SB_LUT4 add_43_9_lut (.I0(n6_adj_4059), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n30685), .O(n35022)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n22338));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n22337));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n22336));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n22335));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n22334));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n22333));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk32MHz), 
           .D(n41163));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk32MHz), 
           .D(n41164));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n22315));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n22314));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n22313));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(clk32MHz), .D(n22312));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n22311));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n22310));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n22309));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n22655));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n22654));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n22653));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n22652));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n22651));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n22650));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n22649));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n22648));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n22647));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n22646));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n22645));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n22644));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n22643));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n22642));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n22641));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n22640));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n22639));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n22638));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n22637));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n22636));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n22635));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n22634));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n22633));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n22632));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n22631));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n22630));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n22629));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n22628));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n22627));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n22626));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n22625));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1351 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(n36222), .I3(GND_net), .O(n1168));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_3_lut_adj_1351.LUT_INIT = 16'h9696;
    SB_LUT4 i14122_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35578), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n22525));
    defparam i14122_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14123_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35578), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n22526));
    defparam i14123_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1352 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[5] [5]), .I3(GND_net), .O(n36020));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1352.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1353 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[9] [7]), .I3(\data_out_frame[7] [5]), .O(n36024));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut_adj_1353.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1354 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[9] [6]), .I3(GND_net), .O(n36287));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1354.LUT_INIT = 16'h9696;
    SB_LUT4 i26398_2_lut_3_lut (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n36412));
    defparam i26398_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_1355 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n20771), .I3(\FRAME_MATCHER.state [2]), .O(n28158));
    defparam i2_3_lut_4_lut_adj_1355.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1356 (.I0(\data_out_frame[9] [5]), .I1(n21216), 
            .I2(\data_out_frame[7] [4]), .I3(n35792), .O(n21026));
    defparam i2_3_lut_4_lut_adj_1356.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1357 (.I0(\data_out_frame[9] [5]), .I1(n21216), 
            .I2(n36287), .I3(GND_net), .O(n6_adj_4148));
    defparam i1_2_lut_3_lut_adj_1357.LUT_INIT = 16'h9696;
    SB_LUT4 i18595_2_lut_3_lut (.I0(n63_adj_4045), .I1(n63), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n92[1]));   // verilog/coms.v(139[4] 141[7])
    defparam i18595_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 add_3971_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n30713), .O(n8825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut_3_lut_adj_1358 (.I0(n63_adj_4045), .I1(n63), .I2(n63_adj_4174), 
            .I3(GND_net), .O(n17985));   // verilog/coms.v(139[4] 141[7])
    defparam i2_2_lut_3_lut_adj_1358.LUT_INIT = 16'h8080;
    SB_LUT4 i12_2_lut_3_lut (.I0(n36146), .I1(n35881), .I2(n21420), .I3(GND_net), 
            .O(n36_adj_4147));
    defparam i12_2_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 equal_112_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4034));
    defparam equal_112_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 mux_1315_i2_3_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n4915), .I3(GND_net), .O(n4917));
    defparam mux_1315_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 equal_113_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [2]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));
    defparam equal_113_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n22624));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n22623));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n22622));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n22621));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n22620));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n22619));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n22618));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n22617));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n22616));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n22615));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n22614));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n22613));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n22612));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n22611));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n22610));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n22609));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n22608));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n22607));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n22606));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n22605));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n22604));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n22603));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n22602));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n22601));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n22600));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n22599));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n22598));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n22597));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n22596));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n22595));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n22594));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n22593));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n22592));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n22591));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n22590));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n22589));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n22588));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n22587));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1359 (.I0(tx_transmit_N_3354), .I1(n27000), 
            .I2(n20700), .I3(n36850), .O(n35589));   // verilog/coms.v(214[11:56])
    defparam i1_3_lut_4_lut_adj_1359.LUT_INIT = 16'h0eff;
    SB_LUT4 i14124_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35578), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n22527));
    defparam i14124_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n22586));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n22585));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(clk32MHz), 
           .D(n22584));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(clk32MHz), 
           .D(n22583));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(clk32MHz), 
           .D(n22582));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(clk32MHz), 
           .D(n22581));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(clk32MHz), 
           .D(n22580));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(clk32MHz), 
           .D(n22579));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1360 (.I0(tx_transmit_N_3354), .I1(n27000), 
            .I2(n17985), .I3(n20700), .O(n3_adj_4000));   // verilog/coms.v(214[11:56])
    defparam i1_3_lut_4_lut_adj_1360.LUT_INIT = 16'h00e0;
    SB_LUT4 i5_3_lut_4_lut_adj_1361 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[11] [3]), .I3(n10_adj_4133), .O(n32865));   // verilog/coms.v(85[17:28])
    defparam i5_3_lut_4_lut_adj_1361.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(clk32MHz), 
           .D(n22578));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(clk32MHz), 
           .D(n22577));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(clk32MHz), 
           .D(n22576));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(clk32MHz), 
           .D(n22575));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(clk32MHz), 
           .D(n22574));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(clk32MHz), 
           .D(n22573));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(clk32MHz), 
           .D(n22572));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(clk32MHz), 
           .D(n22571));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(clk32MHz), 
           .D(n22570));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(clk32MHz), 
           .D(n22569));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(clk32MHz), 
           .D(n22568));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(clk32MHz), 
           .D(n22567));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(clk32MHz), 
           .D(n22566));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(clk32MHz), 
           .D(n22565));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(clk32MHz), 
           .D(n22564));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(clk32MHz), 
           .D(n22563));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n22292));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(clk32MHz), 
           .D(n22562));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14125_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35578), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n22528));
    defparam i14125_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1362 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[7] [2]), .I3(GND_net), .O(n6_adj_4154));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1362.LUT_INIT = 16'h9696;
    SB_CARRY add_3971_6 (.CI(n30713), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n30714));
    SB_LUT4 i28397_4_lut (.I0(\data_out_frame[6] [7]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [7]), 
            .O(n38425));
    defparam i28397_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 add_3971_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n30712), .O(n8825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14126_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35578), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n22529));
    defparam i14126_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i28395_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n38423));
    defparam i28395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1363 (.I0(\FRAME_MATCHER.state [14]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35104));
    defparam i1_2_lut_adj_1363.LUT_INIT = 16'h8888;
    SB_LUT4 i2_2_lut_3_lut_adj_1364 (.I0(n21249), .I1(n33064), .I2(n33015), 
            .I3(GND_net), .O(n6_adj_4113));
    defparam i2_2_lut_3_lut_adj_1364.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i16_3_lut (.I0(\data_out_frame[16] [1]), 
            .I1(\data_out_frame[17] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4247));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i8_3_lut_4_lut (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[8] [3]), 
            .I2(\data_out_frame[11] [6]), .I3(\data_out_frame[12] [3]), 
            .O(n23_adj_4143));
    defparam i8_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1980746_i1_3_lut (.I0(n40813), .I1(n40807), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4237));
    defparam i1980746_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_3_lut_adj_1365 (.I0(n21249), .I1(n33064), .I2(\data_out_frame[23] [3]), 
            .I3(GND_net), .O(n6_adj_4219));
    defparam i2_2_lut_3_lut_adj_1365.LUT_INIT = 16'h9696;
    SB_LUT4 i18633_2_lut_4_lut (.I0(n20704), .I1(n20792), .I2(rx_data_ready), 
            .I3(\FRAME_MATCHER.rx_data_ready_prev ), .O(n27024));
    defparam i18633_2_lut_4_lut.LUT_INIT = 16'h0070;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i17_3_lut (.I0(\data_out_frame[18] [1]), 
            .I1(\data_out_frame[19] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4248));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_2_lut_3_lut_adj_1366 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[6] [6]), .I3(GND_net), .O(n10_adj_4132));   // verilog/coms.v(76[16:27])
    defparam i2_2_lut_3_lut_adj_1366.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1367 (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[8] [7]), 
            .I2(\data_out_frame[7] [1]), .I3(\data_out_frame[9] [2]), .O(n35771));   // verilog/coms.v(71[16:69])
    defparam i2_3_lut_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_LUT4 i29503_2_lut (.I0(\data_out_frame[23] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39277));
    defparam i29503_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1368 (.I0(n20629), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n20704));   // verilog/coms.v(254[5:25])
    defparam i1_2_lut_3_lut_adj_1368.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_adj_1369 (.I0(\FRAME_MATCHER.state [13]), .I1(n11), 
            .I2(GND_net), .I3(GND_net), .O(n35106));
    defparam i1_2_lut_adj_1369.LUT_INIT = 16'h8888;
    SB_LUT4 i14127_3_lut_4_lut (.I0(n8_adj_4034), .I1(n35578), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n22530));
    defparam i14127_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i29502_2_lut (.I0(\data_out_frame[20] [1]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39276));
    defparam i29502_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1370 (.I0(n33939), .I1(n21333), .I2(n33963), 
            .I3(GND_net), .O(n6_adj_4112));
    defparam i1_2_lut_3_lut_adj_1370.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1371 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[4] [3]), 
            .I2(\data_out_frame[6] [4]), .I3(\data_out_frame[8] [6]), .O(n21812));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1371.LUT_INIT = 16'h6996;
    SB_CARRY add_3971_5 (.CI(n30712), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n30713));
    SB_LUT4 i3_2_lut_3_lut (.I0(n33939), .I1(n21333), .I2(\data_out_frame[18] [5]), 
            .I3(GND_net), .O(n12_adj_4151));
    defparam i3_2_lut_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[3] ), 
            .I3(\state[2] ), .O(n3957));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h001a;
    SB_LUT4 i19545_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(n15_adj_3), .O(scl_enable_N_3958));
    defparam i19545_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i14112_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35578), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n22515));
    defparam i14112_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1372 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[11] [0]), 
            .I2(\data_out_frame[4] [4]), .I3(n4_adj_4125), .O(n9_adj_4130));   // verilog/coms.v(73[16:42])
    defparam i1_3_lut_4_lut_adj_1372.LUT_INIT = 16'h6996;
    SB_LUT4 i14113_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35578), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n22516));
    defparam i14113_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i16_3_lut (.I0(\data_out_frame[16] [2]), 
            .I1(\data_out_frame[17] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4250));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1373 (.I0(n1), .I1(n20792), .I2(n11_adj_3975), 
            .I3(\FRAME_MATCHER.state [17]), .O(n35100));
    defparam i1_2_lut_4_lut_adj_1373.LUT_INIT = 16'hba00;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i17_3_lut (.I0(\data_out_frame[18] [2]), 
            .I1(\data_out_frame[19] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4251));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3971_4_lut (.I0(GND_net), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(n30711), .O(n8825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29507_2_lut (.I0(\data_out_frame[23] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39265));
    defparam i29507_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29509_2_lut (.I0(\data_out_frame[20] [2]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39264));
    defparam i29509_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14114_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35578), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n22517));
    defparam i14114_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i16_3_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\data_out_frame[17] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4252));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1374 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n27024), .O(n35578));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1374.LUT_INIT = 16'hfeff;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i17_3_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\data_out_frame[19] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4253));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29511_2_lut (.I0(\data_out_frame[23] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39262));
    defparam i29511_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29513_2_lut (.I0(\data_out_frame[20] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39261));
    defparam i29513_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_3971_4 (.CI(n30711), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n30712));
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(clk32MHz), 
           .D(n22561));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1375 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n27024), .O(n35560));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1375.LUT_INIT = 16'hefff;
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(clk32MHz), .D(n22560));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1376 (.I0(n21_adj_4138), .I1(n19_adj_4137), 
            .I2(n20_adj_4136), .I3(n35820), .O(n6_adj_4114));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i16_3_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\data_out_frame[17] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4254));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i17_3_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\data_out_frame[19] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4255));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29514_2_lut (.I0(\data_out_frame[23] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39259));
    defparam i29514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29516_2_lut (.I0(\data_out_frame[20] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39258));
    defparam i29516_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i16_3_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\data_out_frame[17] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4256));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i17_3_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\data_out_frame[19] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4257));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29517_2_lut (.I0(\data_out_frame[23] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39256));
    defparam i29517_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29519_2_lut (.I0(\data_out_frame[20] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39255));
    defparam i29519_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_adj_1377 (.I0(n21_adj_4138), .I1(n19_adj_4137), 
            .I2(n20_adj_4136), .I3(n36204), .O(n33815));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i16_3_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\data_out_frame[17] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4258));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i17_3_lut (.I0(\data_out_frame[18] [6]), 
            .I1(\data_out_frame[19] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4259));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29520_2_lut (.I0(\data_out_frame[23] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39253));
    defparam i29520_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29522_2_lut (.I0(\data_out_frame[20] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39252));
    defparam i29522_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_2_lut_3_lut_adj_1378 (.I0(\data_out_frame[13] [6]), .I1(n21032), 
            .I2(n33813), .I3(GND_net), .O(n6_adj_4111));
    defparam i2_2_lut_3_lut_adj_1378.LUT_INIT = 16'h9696;
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(clk32MHz), .D(n22559));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(clk32MHz), .D(n22558));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1379 (.I0(\data_out_frame[13] [6]), .I1(n21032), 
            .I2(n32865), .I3(GND_net), .O(n35785));
    defparam i1_2_lut_3_lut_adj_1379.LUT_INIT = 16'h9696;
    SB_LUT4 add_3971_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n30710), .O(n8825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(clk32MHz), .D(n22557));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(clk32MHz), .D(n22556));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(clk32MHz), .D(n22555));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(clk32MHz), .D(n22554));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(clk32MHz), .D(n22553));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(clk32MHz), .D(n22552));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i16_3_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\data_out_frame[17] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4260));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(clk32MHz), .D(n22551));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(clk32MHz), .D(n22550));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(clk32MHz), .D(n22549));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(clk32MHz), .D(n22548));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(clk32MHz), .D(n22547));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(clk32MHz), .D(n22546));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(clk32MHz), .D(n22545));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i17_3_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\data_out_frame[19] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4261));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(clk32MHz), .D(n22544));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(clk32MHz), .D(n22543));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(clk32MHz), .D(n22542));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(clk32MHz), .D(n22541));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(clk32MHz), .D(n22540));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(clk32MHz), .D(n22539));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(clk32MHz), .D(n22538));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n22537));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n22536));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n22535));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n22534));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n22533));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14115_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35578), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n22518));
    defparam i14115_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n22532));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14116_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35578), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n22519));
    defparam i14116_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n22531));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n22530));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n22529));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n22528));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n22527));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n22526));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n22525));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n22524));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n22523));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n22522));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n22521));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n22520));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n22519));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n22518));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n22517));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n22516));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n22515));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n22514));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n22513));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n22512));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i29523_2_lut (.I0(\data_out_frame[23] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39250));
    defparam i29523_2_lut.LUT_INIT = 16'h8888;
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n22511));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n22510));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n22509));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i29527_2_lut (.I0(\data_out_frame[20] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39249));
    defparam i29527_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n22508));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n22507));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n22506));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n22505));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n22504));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n22503));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n22502));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n22501));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n22500));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n22499));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n22498));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n22497));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n22496));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n22495));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n22494));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n22493));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n22492));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n22491));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n22490));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n22489));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n22488));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n22487));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n22486));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n22485));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n22484));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n22483));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n22482));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n22481));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n22480));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n22479));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n22478));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n22477));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n22476));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n22475));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n22474));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n22473));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n22472));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n22471));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14117_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35578), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n22520));
    defparam i14117_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n22470));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1380 (.I0(\FRAME_MATCHER.state [1]), 
            .I1(n20771), .I2(\FRAME_MATCHER.state [0]), .I3(\FRAME_MATCHER.state [3]), 
            .O(n20792));   // verilog/coms.v(151[5:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1380.LUT_INIT = 16'hffef;
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n22469));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n22468));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i29499_2_lut (.I0(n40879), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n39248));
    defparam i29499_2_lut.LUT_INIT = 16'h2222;
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n22467));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n22466));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1381 (.I0(\FRAME_MATCHER.state [1]), .I1(n20771), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n20789));   // verilog/coms.v(151[5:27])
    defparam i1_2_lut_3_lut_adj_1381.LUT_INIT = 16'hfefe;
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n22465));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1382 (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n5180));
    defparam i1_2_lut_3_lut_adj_1382.LUT_INIT = 16'h0202;
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n22464));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n22463));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n22462));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n22461));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n22460));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n22459));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n22458));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n22457));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n22456));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n22455));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n22454));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n22453));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n22452));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n22451));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n22450));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n22449));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n22448));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n22447));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n22446));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n22445));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1383 (.I0(\FRAME_MATCHER.state [3]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n20771), .I3(GND_net), .O(n20629));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1383.LUT_INIT = 16'hfbfb;
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n22444));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i13735_2_lut (.I0(n35), .I1(n20700), .I2(GND_net), .I3(GND_net), 
            .O(n22138));   // verilog/coms.v(127[12] 300[6])
    defparam i13735_2_lut.LUT_INIT = 16'h4444;
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n22443));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n22442));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n22441));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n22440));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n22439));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n22438));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n22437));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n22436));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n22435));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n22434));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n22433));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n22432));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14118_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35578), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n22521));
    defparam i14118_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_3971_3 (.CI(n30710), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n30711));
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n22431));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n22430));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n22429));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i14119_3_lut_4_lut (.I0(n8_adj_4087), .I1(n35578), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n22522));
    defparam i14119_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n22428));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n22427));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n22426));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1384 (.I0(\data_out_frame[13] [1]), .I1(n33493), 
            .I2(n35871), .I3(GND_net), .O(n36146));
    defparam i1_2_lut_3_lut_adj_1384.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1385 (.I0(\data_out_frame[23] [5]), .I1(n21249), 
            .I2(n35945), .I3(\data_out_frame[24] [0]), .O(n6_adj_4080));
    defparam i1_2_lut_3_lut_4_lut_adj_1385.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n22425));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n22424));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_4_lut_adj_1386 (.I0(\data_out_frame[23] [5]), .I1(n21249), 
            .I2(n21586), .I3(n10_adj_4221), .O(n35904));
    defparam i5_3_lut_4_lut_adj_1386.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30822 (.I0(byte_transmit_counter[1]), 
            .I1(n39249), .I2(n39250), .I3(byte_transmit_counter[2]), .O(n40708));
    defparam byte_transmit_counter_1__bdd_4_lut_30822.LUT_INIT = 16'he4aa;
    SB_LUT4 n40708_bdd_4_lut (.I0(n40708), .I1(n17_adj_4261), .I2(n16_adj_4260), 
            .I3(byte_transmit_counter[2]), .O(n40711));
    defparam n40708_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_out_frame[23] [5]), .I1(n21249), 
            .I2(\data_out_frame[23] [6]), .I3(\data_out_frame[24] [0]), 
            .O(n22_adj_4096));
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1387 (.I0(n33064), .I1(\data_out_frame[20] [6]), 
            .I2(n36014), .I3(n36164), .O(n32876));
    defparam i2_3_lut_4_lut_adj_1387.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1388 (.I0(n33064), .I1(\data_out_frame[20] [6]), 
            .I2(n19038), .I3(n35948), .O(n37273));
    defparam i2_3_lut_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1389 (.I0(n33015), .I1(n37273), .I2(n10_adj_4109), 
            .I3(\data_out_frame[23] [0]), .O(n35983));
    defparam i5_3_lut_4_lut_adj_1389.LUT_INIT = 16'h9669;
    SB_LUT4 i14104_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35578), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n22507));
    defparam i14104_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14105_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35578), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n22508));
    defparam i14105_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14106_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35578), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n22509));
    defparam i14106_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1390 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [4]), 
            .I2(n36014), .I3(n35917), .O(n37644));   // verilog/coms.v(85[17:63])
    defparam i2_3_lut_4_lut_adj_1390.LUT_INIT = 16'h6996;
    SB_LUT4 i14107_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35578), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n22510));
    defparam i14107_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1391 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[3] [7]), .I3(\data_in_frame[4] [0]), .O(n35844));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1392 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(n36136), .I3(n36200), .O(n33831));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_4_lut_adj_1392.LUT_INIT = 16'h9669;
    SB_LUT4 i14108_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35578), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n22511));
    defparam i14108_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14109_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35578), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n22512));
    defparam i14109_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1393 (.I0(\data_in_frame[1] [5]), .I1(n35768), 
            .I2(n35844), .I3(\data_in_frame[1] [6]), .O(Kp_23__N_777));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_4_lut_adj_1393.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1394 (.I0(n1), .I1(n20792), .I2(n11_adj_3975), 
            .I3(\FRAME_MATCHER.state [26]), .O(n34990));
    defparam i1_2_lut_4_lut_adj_1394.LUT_INIT = 16'hba00;
    SB_LUT4 i5644_2_lut_3_lut (.I0(n32519), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n63_adj_4174), .I3(GND_net), .O(n13961));   // verilog/coms.v(157[9:60])
    defparam i5644_2_lut_3_lut.LUT_INIT = 16'hd0d0;
    SB_LUT4 i14110_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35578), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n22513));
    defparam i14110_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1395 (.I0(\data_in_frame[1] [5]), .I1(n35768), 
            .I2(\data_in_frame[6] [0]), .I3(\data_in_frame[3] [6]), .O(n36102));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1395.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1396 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[6] [6]), 
            .I2(\data_in_frame[6] [1]), .I3(\data_in_frame[6] [5]), .O(n35805));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1396.LUT_INIT = 16'h6996;
    SB_LUT4 i14111_3_lut_4_lut (.I0(n8_adj_4103), .I1(n35578), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n22514));
    defparam i14111_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1397 (.I0(\data_in_frame[6] [7]), .I1(\data_in_frame[6] [6]), 
            .I2(n10_adj_4072), .I3(\data_in_frame[4] [6]), .O(n21085));   // verilog/coms.v(85[17:28])
    defparam i5_3_lut_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1398 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [4]), 
            .I3(GND_net), .O(n35120));
    defparam i1_2_lut_3_lut_adj_1398.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30688 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n40696));
    defparam byte_transmit_counter_0__bdd_4_lut_30688.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1399 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[3] [2]), 
            .I2(n36081), .I3(GND_net), .O(n6_adj_4057));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1399.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1400 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[3] [2]), 
            .I2(\data_in_frame[5] [5]), .I3(GND_net), .O(n36072));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1400.LUT_INIT = 16'h9696;
    SB_LUT4 i19064_2_lut_4_lut (.I0(n31_adj_4090), .I1(n31), .I2(\FRAME_MATCHER.state [1]), 
            .I3(n18279), .O(n1_adj_4246));
    defparam i19064_2_lut_4_lut.LUT_INIT = 16'hffca;
    SB_LUT4 i3_2_lut_4_lut (.I0(n31_adj_4090), .I1(n31), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state [3]), .O(n11_adj_4101));
    defparam i3_2_lut_4_lut.LUT_INIT = 16'hffca;
    SB_LUT4 i1_2_lut_3_lut_adj_1401 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [5]), 
            .I3(GND_net), .O(n35122));
    defparam i1_2_lut_3_lut_adj_1401.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1402 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [6]), 
            .I3(GND_net), .O(n7_adj_4093));
    defparam i1_2_lut_3_lut_adj_1402.LUT_INIT = 16'he0e0;
    SB_LUT4 n40696_bdd_4_lut (.I0(n40696), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n40699));
    defparam n40696_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1403 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[8] [2]), .I3(GND_net), .O(n35656));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1403.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1404 (.I0(\data_out_frame[11] [6]), .I1(n21026), 
            .I2(n21227), .I3(\data_out_frame[14] [0]), .O(n35980));
    defparam i2_3_lut_4_lut_adj_1404.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1405 (.I0(n37037), .I1(\data_out_frame[24] [4]), 
            .I2(\data_out_frame[24] [3]), .I3(GND_net), .O(n36247));
    defparam i1_2_lut_3_lut_adj_1405.LUT_INIT = 16'h6969;
    SB_LUT4 i2_2_lut_3_lut_adj_1406 (.I0(n37037), .I1(\data_out_frame[24] [4]), 
            .I2(\data_out_frame[24] [5]), .I3(GND_net), .O(n7_adj_4086));
    defparam i2_2_lut_3_lut_adj_1406.LUT_INIT = 16'h6969;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30669 (.I0(byte_transmit_counter[1]), 
            .I1(n39252), .I2(n39253), .I3(byte_transmit_counter[2]), .O(n40690));
    defparam byte_transmit_counter_1__bdd_4_lut_30669.LUT_INIT = 16'he4aa;
    SB_LUT4 i5_3_lut_4_lut_adj_1407 (.I0(\data_in_frame[2] [4]), .I1(n35647), 
            .I2(n35811), .I3(\data_in_frame[1] [7]), .O(n22_adj_4229));   // verilog/coms.v(166[9:87])
    defparam i5_3_lut_4_lut_adj_1407.LUT_INIT = 16'h0990;
    SB_LUT4 i2_3_lut_4_lut_adj_1408 (.I0(\data_in_frame[2] [4]), .I1(n35647), 
            .I2(\data_in_frame[4] [4]), .I3(n21440), .O(n35702));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1409 (.I0(\data_in_frame[2] [4]), .I1(n35647), 
            .I2(\data_in_frame[7] [2]), .I3(n10_adj_4070), .O(n11_adj_4061));   // verilog/coms.v(166[9:87])
    defparam i5_3_lut_4_lut_adj_1409.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1410 (.I0(\data_in_frame[2] [4]), .I1(n35647), 
            .I2(n21436), .I3(\data_in_frame[4] [5]), .O(n21797));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_4_lut_adj_1410.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1411 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [7]), 
            .I3(GND_net), .O(n35124));
    defparam i1_2_lut_3_lut_adj_1411.LUT_INIT = 16'he0e0;
    SB_LUT4 n40690_bdd_4_lut (.I0(n40690), .I1(n17_adj_4259), .I2(n16_adj_4258), 
            .I3(byte_transmit_counter[2]), .O(n40693));
    defparam n40690_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1412 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [8]), 
            .I3(GND_net), .O(n7_adj_4091));
    defparam i1_2_lut_3_lut_adj_1412.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1413 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [9]), 
            .I3(GND_net), .O(n35126));
    defparam i1_2_lut_3_lut_adj_1413.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_2_lut_3_lut_adj_1414 (.I0(n21420), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[15] [0]), .I3(GND_net), .O(n35777));
    defparam i2_2_lut_3_lut_adj_1414.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1415 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[11] [6]), 
            .I2(n36124), .I3(\data_out_frame[14] [0]), .O(n35935));
    defparam i1_2_lut_4_lut_adj_1415.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1416 (.I0(\data_out_frame[16] [0]), .I1(\data_out_frame[13] [6]), 
            .I2(n21032), .I3(n32865), .O(n36115));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_4_lut_adj_1416.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1417 (.I0(n37273), .I1(\data_out_frame[24] [7]), 
            .I2(n10_adj_4107), .I3(GND_net), .O(n32920));
    defparam i5_3_lut_4_lut_adj_1417.LUT_INIT = 16'h6969;
    SB_LUT4 i18616_2_lut_3_lut (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [10]), 
            .I3(GND_net), .O(n27005));
    defparam i18616_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut_adj_1418 (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[1] [5]), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[1] [6]), .O(n6_adj_4106));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_4_lut_adj_1418.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1419 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [6]), .I3(GND_net), .O(n35727));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_3_lut_adj_1419.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1420 (.I0(n32519), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n17985), .I3(GND_net), .O(n17948));   // verilog/coms.v(157[9:60])
    defparam i1_2_lut_3_lut_adj_1420.LUT_INIT = 16'hd0d0;
    SB_LUT4 i1_2_lut_3_lut_adj_1421 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [11]), 
            .I3(GND_net), .O(n35128));
    defparam i1_2_lut_3_lut_adj_1421.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1422 (.I0(\data_in_frame[3] [0]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(GND_net), .O(n36054));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1422.LUT_INIT = 16'h9696;
    SB_LUT4 i18617_2_lut_3_lut (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [12]), 
            .I3(GND_net), .O(n27007));
    defparam i18617_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_4_lut_adj_1423 (.I0(n21440), .I1(n35684), .I2(\data_in_frame[1] [7]), 
            .I3(\data_in_frame[1] [6]), .O(Kp_23__N_937));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_4_lut_adj_1423.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1424 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n21440));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1424.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1425 (.I0(n33928), .I1(\data_out_frame[20] [2]), 
            .I2(n37037), .I3(GND_net), .O(n33327));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1425.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1426 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [13]), 
            .I3(GND_net), .O(n35130));
    defparam i1_2_lut_3_lut_adj_1426.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30655 (.I0(byte_transmit_counter[1]), 
            .I1(n39255), .I2(n39256), .I3(byte_transmit_counter[2]), .O(n40684));
    defparam byte_transmit_counter_1__bdd_4_lut_30655.LUT_INIT = 16'he4aa;
    SB_LUT4 n40684_bdd_4_lut (.I0(n40684), .I1(n17_adj_4257), .I2(n16_adj_4256), 
            .I3(byte_transmit_counter[2]), .O(n40687));
    defparam n40684_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1427 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [14]), 
            .I3(GND_net), .O(n35132));
    defparam i1_2_lut_3_lut_adj_1427.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30650 (.I0(byte_transmit_counter[1]), 
            .I1(n39258), .I2(n39259), .I3(byte_transmit_counter[2]), .O(n40678));
    defparam byte_transmit_counter_1__bdd_4_lut_30650.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1428 (.I0(\data_out_frame[20] [3]), .I1(n35917), 
            .I2(n36164), .I3(GND_net), .O(n33928));
    defparam i1_2_lut_3_lut_adj_1428.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_3_lut_4_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[4] [2]), .I3(\data_out_frame[5] [7]), .O(n36030));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1429 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[4] [4]), 
            .I2(\data_in_frame[2] [1]), .I3(GND_net), .O(n6_adj_4104));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1429.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1430 (.I0(\data_out_frame[24] [5]), .I1(\data_out_frame[24] [6]), 
            .I2(n36178), .I3(GND_net), .O(n6_adj_4088));
    defparam i1_2_lut_3_lut_adj_1430.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1431 (.I0(n35840), .I1(n36151), .I2(\data_out_frame[20] [1]), 
            .I3(\data_out_frame[19] [7]), .O(n36178));
    defparam i2_3_lut_4_lut_adj_1431.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1432 (.I0(n33954), .I1(n35975), .I2(\data_out_frame[19] [7]), 
            .I3(\data_out_frame[19] [6]), .O(n32951));
    defparam i2_3_lut_4_lut_adj_1432.LUT_INIT = 16'h6996;
    SB_LUT4 n40678_bdd_4_lut (.I0(n40678), .I1(n17_adj_4255), .I2(n16_adj_4254), 
            .I3(byte_transmit_counter[2]), .O(n40681));
    defparam n40678_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1433 (.I0(n36146), .I1(n35881), .I2(n35975), 
            .I3(GND_net), .O(n35926));
    defparam i1_2_lut_3_lut_adj_1433.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30645 (.I0(byte_transmit_counter[1]), 
            .I1(n39261), .I2(n39262), .I3(byte_transmit_counter[2]), .O(n40672));
    defparam byte_transmit_counter_1__bdd_4_lut_30645.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1434 (.I0(n33886), .I1(\data_out_frame[15] [1]), 
            .I2(\data_out_frame[19] [5]), .I3(GND_net), .O(n36278));
    defparam i1_2_lut_3_lut_adj_1434.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1435 (.I0(\data_in_frame[8] [5]), .I1(n35751), 
            .I2(n7_adj_4234), .I3(GND_net), .O(n35644));
    defparam i1_2_lut_3_lut_adj_1435.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1436 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [15]), 
            .I3(GND_net), .O(n35134));
    defparam i1_2_lut_3_lut_adj_1436.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_4_lut_adj_1437 (.I0(\data_in_frame[8] [5]), .I1(n35751), 
            .I2(n32855), .I3(\data_in_frame[9] [0]), .O(n36078));
    defparam i2_3_lut_4_lut_adj_1437.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1438 (.I0(\data_in_frame[8] [5]), .I1(n35751), 
            .I2(\data_in_frame[12] [7]), .I3(GND_net), .O(n35789));
    defparam i1_2_lut_3_lut_adj_1438.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1439 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [16]), 
            .I3(GND_net), .O(n35136));
    defparam i1_2_lut_3_lut_adj_1439.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_4_lut_adj_1440 (.I0(\data_in_frame[8] [5]), .I1(n35751), 
            .I2(\data_in_frame[8] [0]), .I3(n33831), .O(n18_adj_4244));
    defparam i2_3_lut_4_lut_adj_1440.LUT_INIT = 16'hf66f;
    SB_LUT4 i1_2_lut_3_lut_adj_1441 (.I0(\data_out_frame[24] [2]), .I1(\data_out_frame[24] [1]), 
            .I2(n33872), .I3(GND_net), .O(n6_adj_4082));
    defparam i1_2_lut_3_lut_adj_1441.LUT_INIT = 16'h9696;
    SB_LUT4 n40672_bdd_4_lut (.I0(n40672), .I1(n17_adj_4253), .I2(n16_adj_4252), 
            .I3(byte_transmit_counter[2]), .O(n40675));
    defparam n40672_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30640 (.I0(byte_transmit_counter[1]), 
            .I1(n39264), .I2(n39265), .I3(byte_transmit_counter[2]), .O(n40666));
    defparam byte_transmit_counter_1__bdd_4_lut_30640.LUT_INIT = 16'he4aa;
    SB_LUT4 i5_3_lut_4_lut_adj_1442 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(n10_adj_4066), .I3(n35671), .O(n20900));   // verilog/coms.v(76[16:43])
    defparam i5_3_lut_4_lut_adj_1442.LUT_INIT = 16'h6996;
    SB_LUT4 i28273_2_lut_3_lut (.I0(n21181), .I1(n35814), .I2(n21127), 
            .I3(GND_net), .O(n38300));
    defparam i28273_2_lut_3_lut.LUT_INIT = 16'h6060;
    SB_LUT4 n40666_bdd_4_lut (.I0(n40666), .I1(n17_adj_4251), .I2(n16_adj_4250), 
            .I3(byte_transmit_counter[2]), .O(n40669));
    defparam n40666_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_30635 (.I0(byte_transmit_counter[1]), 
            .I1(n39276), .I2(n39277), .I3(byte_transmit_counter[2]), .O(n40660));
    defparam byte_transmit_counter_1__bdd_4_lut_30635.LUT_INIT = 16'he4aa;
    SB_LUT4 n40660_bdd_4_lut (.I0(n40660), .I1(n17_adj_4248), .I2(n16_adj_4247), 
            .I3(byte_transmit_counter[2]), .O(n40663));
    defparam n40660_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30660 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n40648));
    defparam byte_transmit_counter_0__bdd_4_lut_30660.LUT_INIT = 16'he4aa;
    SB_LUT4 n40648_bdd_4_lut (.I0(n40648), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n40651));
    defparam n40648_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_4_lut_adj_1443 (.I0(n21181), .I1(n35814), .I2(n21127), 
            .I3(Kp_23__N_1147), .O(n32664));
    defparam i2_3_lut_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1444 (.I0(n21181), .I1(n35814), .I2(n36099), 
            .I3(n4_adj_4069), .O(n36308));
    defparam i1_2_lut_3_lut_4_lut_adj_1444.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1445 (.I0(\data_out_frame[19] [2]), .I1(n33963), 
            .I2(n10_adj_4079), .I3(\data_out_frame[25] [6]), .O(n36761));
    defparam i5_3_lut_4_lut_adj_1445.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1446 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[4] [5]), 
            .I2(n35702), .I3(GND_net), .O(n35696));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1446.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1447 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[2] [5]), .I3(GND_net), .O(n20881));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1447.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1448 (.I0(n32987), .I1(n11_adj_4061), .I2(\data_in_frame[11] [5]), 
            .I3(GND_net), .O(n35858));
    defparam i1_2_lut_3_lut_adj_1448.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut_adj_1449 (.I0(n32987), .I1(n11_adj_4061), .I2(n36130), 
            .I3(n33933), .O(n8_adj_4054));
    defparam i3_3_lut_4_lut_adj_1449.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1450 (.I0(\data_in_frame[6] [1]), .I1(Kp_23__N_777), 
            .I2(\data_in_frame[8] [3]), .I3(GND_net), .O(n4_adj_4069));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1450.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1451 (.I0(n32987), .I1(n11_adj_4061), .I2(\data_in_frame[9] [4]), 
            .I3(GND_net), .O(n33890));
    defparam i1_2_lut_3_lut_adj_1451.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1452 (.I0(\data_in_frame[3] [5]), .I1(\data_in_frame[5] [6]), 
            .I2(n21181), .I3(GND_net), .O(n36200));
    defparam i1_2_lut_3_lut_adj_1452.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1453 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(GND_net), .O(n21181));
    defparam i1_2_lut_3_lut_adj_1453.LUT_INIT = 16'h9696;
    SB_LUT4 i3_2_lut_4_lut_adj_1454 (.I0(Kp_23__N_1162), .I1(\data_in_frame[9] [1]), 
            .I2(\data_in_frame[11] [3]), .I3(\data_in_frame[15] [5]), .O(n12_adj_4065));   // verilog/coms.v(75[16:43])
    defparam i3_2_lut_4_lut_adj_1454.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1455 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [17]), 
            .I3(GND_net), .O(n35138));
    defparam i1_2_lut_3_lut_adj_1455.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut_adj_1456 (.I0(Kp_23__N_1162), .I1(\data_in_frame[9] [1]), 
            .I2(\data_in_frame[11] [3]), .I3(\data_in_frame[13] [5]), .O(n36127));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1457 (.I0(n21100), .I1(n11_adj_4061), .I2(\data_in_frame[9] [3]), 
            .I3(GND_net), .O(n20847));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1457.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1458 (.I0(n32987), .I1(n21127), .I2(n11_adj_4061), 
            .I3(n8_adj_4056), .O(n36130));
    defparam i2_3_lut_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1459 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(\data_in_frame[11] [1]), .I3(n33933), .O(n36250));
    defparam i2_3_lut_4_lut_adj_1459.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1460 (.I0(n32987), .I1(n21127), .I2(n33890), 
            .I3(\data_in_frame[9] [5]), .O(n33849));
    defparam i2_3_lut_4_lut_adj_1460.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1461 (.I0(n21085), .I1(n21100), .I2(n36142), 
            .I3(\data_in_frame[11] [4]), .O(n33843));
    defparam i2_3_lut_4_lut_adj_1461.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1462 (.I0(\data_in_frame[11] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(\data_in_frame[9] [2]), .I3(GND_net), .O(n6_adj_4060));   // verilog/coms.v(72[16:41])
    defparam i2_2_lut_3_lut_adj_1462.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1463 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [4]), 
            .I2(n35858), .I3(\data_in_frame[13] [6]), .O(n36142));
    defparam i2_3_lut_4_lut_adj_1463.LUT_INIT = 16'h6996;
    SB_LUT4 i28391_4_lut (.I0(\data_out_frame[6] [6]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [6]), 
            .O(n38419));
    defparam i28391_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i5_3_lut_4_lut_adj_1464 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[10] [7]), 
            .I2(n10_adj_3979), .I3(\data_in_frame[14] [7]), .O(n21568));   // verilog/coms.v(71[16:27])
    defparam i5_3_lut_4_lut_adj_1464.LUT_INIT = 16'h6996;
    SB_LUT4 i28389_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n38417));
    defparam i28389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1465 (.I0(\data_in_frame[11] [2]), .I1(\data_in_frame[9] [0]), 
            .I2(Kp_23__N_1151), .I3(GND_net), .O(n21479));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1465.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1466 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n36078), .I3(GND_net), .O(n6_adj_4055));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_3_lut_adj_1466.LUT_INIT = 16'h9696;
    SB_LUT4 i1981349_i1_3_lut (.I0(n40741), .I1(n40867), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4216));
    defparam i1981349_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29526_2_lut (.I0(n40885), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n39251));
    defparam i29526_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_4_lut_adj_1467 (.I0(\data_in_frame[11] [0]), .I1(\data_in_frame[10] [7]), 
            .I2(\data_in_frame[13] [2]), .I3(n7_adj_4234), .O(n35635));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1467.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1468 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[8] [0]), 
            .I2(n33831), .I3(GND_net), .O(n36265));
    defparam i1_2_lut_3_lut_adj_1468.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1469 (.I0(\data_in_frame[8] [1]), .I1(\data_in_frame[8] [0]), 
            .I2(\data_in_frame[12] [0]), .I3(n32664), .O(n14_adj_4039));
    defparam i5_3_lut_4_lut_adj_1469.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1470 (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[15] [4]), 
            .I2(n33683), .I3(\data_in_frame[13] [2]), .O(n36219));
    defparam i2_3_lut_4_lut_adj_1470.LUT_INIT = 16'h9669;
    SB_LUT4 i28384_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n38412));
    defparam i28384_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1471 (.I0(n63_adj_4045), .I1(n63), .I2(\FRAME_MATCHER.state [1]), 
            .I3(n63_adj_4174), .O(n35587));
    defparam i1_2_lut_4_lut_adj_1471.LUT_INIT = 16'h80ff;
    SB_LUT4 i28385_4_lut (.I0(n38412), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n38413));
    defparam i28385_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i28383_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n38411));
    defparam i28383_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 select_428_Select_2_i7_3_lut_4_lut (.I0(\FRAME_MATCHER.state_31__N_2501 [2]), 
            .I1(n20629), .I2(n20703), .I3(n4452), .O(n7_adj_4047));
    defparam select_428_Select_2_i7_3_lut_4_lut.LUT_INIT = 16'h0302;
    SB_LUT4 i1_2_lut_4_lut_adj_1472 (.I0(\FRAME_MATCHER.state [2]), .I1(n63), 
            .I2(n63_adj_4045), .I3(n63_adj_4174), .O(\FRAME_MATCHER.state_31__N_2501 [2]));   // verilog/coms.v(142[7:84])
    defparam i1_2_lut_4_lut_adj_1472.LUT_INIT = 16'hb300;
    SB_LUT4 i1981952_i1_3_lut (.I0(n40735), .I1(n40789), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4214));
    defparam i1981952_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1473 (.I0(n21085), .I1(\data_in_frame[9] [2]), 
            .I2(n11_adj_4061), .I3(\data_in_frame[9] [3]), .O(n20844));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_4_lut_adj_1473.LUT_INIT = 16'h6996;
    SB_LUT4 i29521_2_lut (.I0(n40891), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n39254));
    defparam i29521_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i28378_3_lut (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[7] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n38406));
    defparam i28378_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28379_4_lut (.I0(n38406), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n38407));
    defparam i28379_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 i28377_3_lut (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[5] [4]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n38405));
    defparam i28377_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1474 (.I0(\data_in_frame[9] [1]), .I1(n32987), 
            .I2(n11_adj_4061), .I3(\data_in_frame[11] [5]), .O(n33950));
    defparam i1_2_lut_4_lut_adj_1474.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_4_lut_adj_1475 (.I0(n35866), .I1(\data_in_frame[8] [5]), 
            .I2(n35751), .I3(n7_adj_4234), .O(n10_adj_4037));
    defparam i2_2_lut_4_lut_adj_1475.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1476 (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_829), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[2] [7]), .O(n21296));
    defparam i1_2_lut_4_lut_adj_1476.LUT_INIT = 16'h6996;
    SB_LUT4 i14128_3_lut_4_lut (.I0(n8), .I1(n35578), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n22531));
    defparam i14128_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1477 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [18]), 
            .I3(GND_net), .O(n35140));
    defparam i1_2_lut_3_lut_adj_1477.LUT_INIT = 16'he0e0;
    SB_LUT4 i14129_3_lut_4_lut (.I0(n8), .I1(n35578), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n22532));
    defparam i14129_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1982555_i1_3_lut (.I0(n40849), .I1(n40831), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4210));
    defparam i1982555_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29518_2_lut (.I0(n40645), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n39257));
    defparam i29518_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i14130_3_lut_4_lut (.I0(n8), .I1(n35578), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n22533));
    defparam i14130_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14131_3_lut_4_lut (.I0(n8), .I1(n35578), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n22534));
    defparam i14131_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14132_3_lut_4_lut (.I0(n8), .I1(n35578), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n22535));
    defparam i14132_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14133_3_lut_4_lut (.I0(n8), .I1(n35578), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n22536));
    defparam i14133_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_4_lut_adj_1478 (.I0(\data_in_frame[8] [5]), .I1(n35751), 
            .I2(\data_in_frame[12] [7]), .I3(\data_in_frame[13] [0]), .O(n10_adj_4007));
    defparam i2_2_lut_4_lut_adj_1478.LUT_INIT = 16'h6996;
    SB_LUT4 i28372_3_lut (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[7] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n38400));
    defparam i28372_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1479 (.I0(n20900), .I1(\data_in_frame[10] [4]), 
            .I2(n35798), .I3(n4_adj_4069), .O(n21171));
    defparam i2_3_lut_4_lut_adj_1479.LUT_INIT = 16'h6996;
    SB_LUT4 i28373_4_lut (.I0(n38400), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n38401));
    defparam i28373_4_lut.LUT_INIT = 16'hafa3;
    SB_LUT4 i28371_3_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[5] [3]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n38399));
    defparam i28371_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_4_lut_adj_1480 (.I0(n21797), .I1(n35849), .I2(n10_c), 
            .I3(n35814), .O(n33952));
    defparam i5_3_lut_4_lut_adj_1480.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_30622 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n40642));
    defparam byte_transmit_counter_0__bdd_4_lut_30622.LUT_INIT = 16'he4aa;
    SB_LUT4 i5_3_lut_4_lut_adj_1481 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[16] [0]), 
            .I2(n10_adj_3999), .I3(n35957), .O(n36155));
    defparam i5_3_lut_4_lut_adj_1481.LUT_INIT = 16'h6996;
    SB_LUT4 i14134_3_lut_4_lut (.I0(n8), .I1(n35578), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n22537));
    defparam i14134_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1984163_i1_3_lut (.I0(n40819), .I1(n40915), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4208));
    defparam i1984163_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29515_2_lut (.I0(n40651), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n39260));
    defparam i29515_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i28366_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n38394));
    defparam i28366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28367_4_lut (.I0(n38394), .I1(byte_transmit_counter[0]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n38395));
    defparam i28367_4_lut.LUT_INIT = 16'ha0a3;
    SB_LUT4 i28365_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n38393));
    defparam i28365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29512_2_lut (.I0(n40699), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n39263));
    defparam i29512_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i28361_4_lut (.I0(\data_out_frame[6] [1]), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[2]), .I3(\data_out_frame[7] [1]), 
            .O(n38389));
    defparam i28361_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i28359_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n38387));
    defparam i28359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1482 (.I0(\data_in_frame[12] [3]), .I1(n36290), 
            .I2(\data_in_frame[10] [1]), .I3(\data_in_frame[9] [7]), .O(n36158));
    defparam i1_2_lut_4_lut_adj_1482.LUT_INIT = 16'h6996;
    SB_LUT4 i1985369_i1_3_lut (.I0(n40801), .I1(n40795), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4205));
    defparam i1985369_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29530_2_lut (.I0(n40903), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n39274));
    defparam i29530_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i13910_3_lut_4_lut (.I0(n8), .I1(n35578), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n22313));
    defparam i13910_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1483 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [19]), 
            .I3(GND_net), .O(n35142));
    defparam i1_2_lut_3_lut_adj_1483.LUT_INIT = 16'he0e0;
    SB_LUT4 i5_3_lut_4_lut_adj_1484 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n10_adj_3982), .I3(\data_in_frame[12] [2]), .O(n37804));
    defparam i5_3_lut_4_lut_adj_1484.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1485 (.I0(n4_adj_4069), .I1(n36099), .I2(\data_in_frame[10] [5]), 
            .I3(\data_in_frame[15] [0]), .O(n36275));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1485.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1486 (.I0(n20900), .I1(\data_in_frame[10] [4]), 
            .I2(n20979), .I3(n36060), .O(n6_adj_3981));
    defparam i1_2_lut_4_lut_adj_1486.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1487 (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[14] [4]), 
            .I2(n10_adj_3980), .I3(n32886), .O(n36060));
    defparam i5_3_lut_4_lut_adj_1487.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1488 (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[16] [7]), 
            .I2(n10_adj_3978), .I3(n33879), .O(n35687));
    defparam i5_3_lut_4_lut_adj_1488.LUT_INIT = 16'h6996;
    SB_LUT4 n40642_bdd_4_lut (.I0(n40642), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n40645));
    defparam n40642_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1489 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [20]), 
            .I3(GND_net), .O(n35144));
    defparam i1_2_lut_3_lut_adj_1489.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1490 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [21]), 
            .I3(GND_net), .O(n35146));
    defparam i1_2_lut_3_lut_adj_1490.LUT_INIT = 16'he0e0;
    SB_LUT4 i19376_1_lut_2_lut (.I0(n20704), .I1(n20792), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4059));
    defparam i19376_1_lut_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i16_3_lut (.I0(\data_out_frame[16] [0]), 
            .I1(\data_out_frame[17] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4200));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i17_3_lut (.I0(\data_out_frame[18] [0]), 
            .I1(\data_out_frame[19] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4199));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_3_lut_4_lut_adj_1491 (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[17] [6]), 
            .I2(n36244), .I3(n33683), .O(n20));   // verilog/coms.v(70[16:27])
    defparam i7_3_lut_4_lut_adj_1491.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1492 (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[17] [6]), 
            .I2(n20847), .I3(GND_net), .O(n7));   // verilog/coms.v(70[16:27])
    defparam i2_2_lut_3_lut_adj_1492.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1493 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [22]), 
            .I3(GND_net), .O(n35148));
    defparam i1_2_lut_3_lut_adj_1493.LUT_INIT = 16'he0e0;
    SB_LUT4 i29475_2_lut (.I0(\data_out_frame[23] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39280));
    defparam i29475_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i29473_2_lut (.I0(\data_out_frame[20] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39279));
    defparam i29473_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i28329_3_lut (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[9] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n38357));
    defparam i28329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28330_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n38358));
    defparam i28330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28321_3_lut (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n38349));
    defparam i28321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28320_3_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n38348));
    defparam i28320_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1494 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [23]), 
            .I3(GND_net), .O(n35150));
    defparam i1_2_lut_3_lut_adj_1494.LUT_INIT = 16'he0e0;
    SB_LUT4 i28357_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n38385));
    defparam i28357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i28358_4_lut (.I0(n38385), .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n38386));
    defparam i28358_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i1_2_lut_3_lut_adj_1495 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [24]), 
            .I3(GND_net), .O(n35152));
    defparam i1_2_lut_3_lut_adj_1495.LUT_INIT = 16'he0e0;
    SB_LUT4 i28356_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n38384));
    defparam i28356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_4_lut_4_lut (.I0(n36090), .I1(n21611), .I2(n37644), 
            .I3(n35716), .O(n32949));
    defparam i4_4_lut_4_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1496 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [25]), 
            .I3(GND_net), .O(n35186));
    defparam i1_2_lut_3_lut_adj_1496.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1497 (.I0(n3_adj_4000), .I1(n2), .I2(\FRAME_MATCHER.state [26]), 
            .I3(GND_net), .O(n35200));
    defparam i1_2_lut_3_lut_adj_1497.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1498 (.I0(n19152), .I1(\data_in_frame[5] [5]), 
            .I2(\data_in_frame[7] [7]), .I3(GND_net), .O(n4_adj_3992));
    defparam i1_2_lut_3_lut_adj_1498.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_4_lut_adj_1499 (.I0(n36850), .I1(n17985), .I2(n36527), 
            .I3(n20792), .O(n11));
    defparam i1_4_lut_4_lut_adj_1499.LUT_INIT = 16'h444c;
    SB_LUT4 i1_3_lut_4_lut_adj_1500 (.I0(n20629), .I1(n20703), .I2(n17985), 
            .I3(n4452), .O(n2));
    defparam i1_3_lut_4_lut_adj_1500.LUT_INIT = 16'h0010;
    SB_LUT4 i1_2_lut_3_lut_adj_1501 (.I0(n20619), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n17985), .I3(GND_net), .O(n18028));   // verilog/coms.v(227[6] 229[9])
    defparam i1_2_lut_3_lut_adj_1501.LUT_INIT = 16'hd0d0;
    SB_LUT4 i1987178_i1_3_lut (.I0(n40861), .I1(n40855), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n14_adj_4195));
    defparam i1987178_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29505_2_lut (.I0(n40909), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n39278));
    defparam i29505_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_4_lut_adj_1502 (.I0(\data_in_frame[6] [4]), .I1(n21440), 
            .I2(n35684), .I3(Kp_23__N_834), .O(n36069));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_4_lut_adj_1502.LUT_INIT = 16'h6996;
    uart_tx tx (.n21920(n21920), .clk32MHz(clk32MHz), .n22195(n22195), 
            .r_SM_Main({r_SM_Main}), .\r_SM_Main_2__N_3454[1] (\r_SM_Main_2__N_3454[1] ), 
            .tx_o(tx_o), .tx_data({tx_data}), .\r_SM_Main_2__N_3457[0] (r_SM_Main_2__N_3457[0]), 
            .n13920(n13920), .GND_net(GND_net), .VCC_net(VCC_net), .\r_Bit_Index[0] (\r_Bit_Index[0] ), 
            .n4(n4), .n22817(n22817), .n22319(n22319), .tx_active(tx_active), 
            .n41168(n41168), .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(107[10:70])
    uart_rx rx (.clk32MHz(clk32MHz), .n22012(n22012), .n22193(n22193), 
            .n26980(n26980), .GND_net(GND_net), .n4(n4_adj_4), .n4_adj_1(n4_adj_5), 
            .\r_Bit_Index[0] (\r_Bit_Index[0]_adj_6 ), .n20781(n20781), 
            .r_Rx_Data(r_Rx_Data), .RX_N_10(RX_N_10), .VCC_net(VCC_net), 
            .n20776(n20776), .n4_adj_2(n4_adj_7), .n22843(n22843), .rx_data_ready(rx_data_ready), 
            .n22847(n22847), .rx_data({rx_data}), .n22308(n22308), .n22307(n22307), 
            .n22306(n22306), .n22305(n22305), .n22304(n22304), .n22303(n22303), 
            .n22302(n22302)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(93[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (n21920, clk32MHz, n22195, r_SM_Main, \r_SM_Main_2__N_3454[1] , 
            tx_o, tx_data, \r_SM_Main_2__N_3457[0] , n13920, GND_net, 
            VCC_net, \r_Bit_Index[0] , n4, n22817, n22319, tx_active, 
            n41168, tx_enable) /* synthesis syn_module_defined=1 */ ;
    output n21920;
    input clk32MHz;
    output n22195;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3454[1] ;
    output tx_o;
    input [7:0]tx_data;
    input \r_SM_Main_2__N_3457[0] ;
    output n13920;
    input GND_net;
    input VCC_net;
    output \r_Bit_Index[0] ;
    output n4;
    input n22817;
    input n22319;
    output tx_active;
    input n41168;
    output tx_enable;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [2:0]n307;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    
    wire n22161, n3, n1, n18035;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n15784;
    wire [8:0]n41;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n31682, n31681, n31680, n31679, n31678, n31677, n31676, 
        n31675, n27562, n15783, n40873, n40717, o_Tx_Serial_N_3485, 
        n10, n37667, n40870, n3_adj_3974, n40714;
    
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .E(n21920), 
            .D(n307[2]), .R(n22195));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .E(n21920), 
            .D(n307[1]), .R(n22195));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i30123_4_lut (.I0(r_SM_Main[2]), .I1(\r_SM_Main_2__N_3454[1] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n22161));
    defparam i30123_4_lut.LUT_INIT = 16'h4445;
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .E(n1), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n18035), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n15784), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i5605_2_lut (.I0(\r_SM_Main_2__N_3457[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n13920));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5605_2_lut.LUT_INIT = 16'h2222;
    SB_DFFESR r_Clock_Count_1513__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), 
            .E(n1), .D(n41[0]), .R(n22161));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1513__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), 
            .E(n1), .D(n41[1]), .R(n22161));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 r_Clock_Count_1513_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n31682), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1513_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1513_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n31681), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1513_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1513_add_4_9 (.CI(n31681), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n31682));
    SB_LUT4 r_Clock_Count_1513_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n31680), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1513_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1513_add_4_8 (.CI(n31680), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n31681));
    SB_LUT4 r_Clock_Count_1513_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n31679), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1513_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1513_add_4_7 (.CI(n31679), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n31680));
    SB_LUT4 r_Clock_Count_1513_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n31678), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1513_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1513_add_4_6 (.CI(n31678), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n31679));
    SB_LUT4 r_Clock_Count_1513_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n31677), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1513_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1513_add_4_5 (.CI(n31677), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n31678));
    SB_LUT4 r_Clock_Count_1513_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n31676), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1513_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1513_add_4_4 (.CI(n31676), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n31677));
    SB_LUT4 r_Clock_Count_1513_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n31675), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1513_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1513_add_4_3 (.CI(n31675), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n31676));
    SB_LUT4 r_Clock_Count_1513_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1513_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1513_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n31675));
    SB_LUT4 i7459_4_lut (.I0(\r_SM_Main_2__N_3457[0] ), .I1(n27562), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3454[1] ), .O(n15783));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7459_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i7460_3_lut (.I0(n15783), .I1(\r_SM_Main_2__N_3454[1] ), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n15784));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i7460_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFESR r_Clock_Count_1513__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), 
            .E(n1), .D(n41[8]), .R(n22161));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1985972_i1_3_lut (.I0(n40873), .I1(n40717), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_3485));
    defparam i1985972_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3485), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_DFFESR r_Clock_Count_1513__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), 
            .E(n1), .D(n41[7]), .R(n22161));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1513__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), 
            .E(n1), .D(n41[6]), .R(n22161));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1513__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), 
            .E(n1), .D(n41[5]), .R(n22161));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1513__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), 
            .E(n1), .D(n41[4]), .R(n22161));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i1611_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n307[1]));   // verilog/uart_tx.v(98[36:51])
    defparam i1611_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n27562));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[0]), 
            .I3(r_Clock_Count[5]), .O(n10));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[3]), .I1(n10), .I2(r_Clock_Count[4]), 
            .I3(GND_net), .O(n37667));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i3_4_lut (.I0(n37667), .I1(r_Clock_Count[8]), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[7]), .O(\r_SM_Main_2__N_3454[1] ));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13792_3_lut (.I0(n21920), .I1(n27562), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n22195));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13792_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1618_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n307[2]));   // verilog/uart_tx.v(98[36:51])
    defparam i1618_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n40870));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n40870_bdd_4_lut (.I0(n40870), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n40873));
    defparam n40870_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFFESR r_Clock_Count_1513__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), 
            .E(n1), .D(n41[3]), .R(n22161));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1513__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), 
            .E(n1), .D(n41[2]), .R(n22161));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(\r_SM_Main_2__N_3454[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n18035), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n18035), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n18035), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n18035), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n18035), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n18035), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n18035), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n3_adj_3974), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i9463_2_lut_3_lut (.I0(\r_SM_Main_2__N_3454[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_3974));
    defparam i9463_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk32MHz), .D(n22817));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3457[0] ), 
            .I3(r_SM_Main[1]), .O(n18035));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_30802 (.I0(\r_Bit_Index[0] ), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n40714));
    defparam r_Bit_Index_0__bdd_4_lut_30802.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3454[1] ), .O(n21920));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n22319));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(n41168));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 n40714_bdd_4_lut (.I0(n40714), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n40717));
    defparam n40714_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (clk32MHz, n22012, n22193, n26980, GND_net, n4, n4_adj_1, 
            \r_Bit_Index[0] , n20781, r_Rx_Data, RX_N_10, VCC_net, 
            n20776, n4_adj_2, n22843, rx_data_ready, n22847, rx_data, 
            n22308, n22307, n22306, n22305, n22304, n22303, n22302) /* synthesis syn_module_defined=1 */ ;
    input clk32MHz;
    output n22012;
    output n22193;
    output n26980;
    input GND_net;
    output n4;
    output n4_adj_1;
    output \r_Bit_Index[0] ;
    output n20781;
    output r_Rx_Data;
    input RX_N_10;
    input VCC_net;
    output n20776;
    output n4_adj_2;
    input n22843;
    output rx_data_ready;
    input n22847;
    output [7:0]rx_data;
    input n22308;
    input n22307;
    input n22306;
    input n22305;
    input n22304;
    input n22303;
    input n22302;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [7:0]n37;
    
    wire n21972;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n22159;
    wire [2:0]n326;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main_2__N_3383;
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n35545, n20583, n14, r_Rx_Data_R, n31674, n31673, n31672, 
        n31671, n31670, n31669, n31668, n27558, n27846, n13, n36, 
        n5, n25159, n25166, n8, n27922, n35192, n21911, n39267;
    
    SB_DFFESR r_Clock_Count_1511__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), 
            .E(n21972), .D(n37[7]), .R(n22159));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1511__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), 
            .E(n21972), .D(n37[6]), .R(n22159));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1511__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), 
            .E(n21972), .D(n37[5]), .R(n22159));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1511__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), 
            .E(n21972), .D(n37[4]), .R(n22159));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1511__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), 
            .E(n21972), .D(n37[3]), .R(n22159));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1511__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), 
            .E(n21972), .D(n37[2]), .R(n22159));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1511__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), 
            .E(n21972), .D(n37[1]), .R(n22159));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .E(n22012), 
            .D(n326[2]), .R(n22193));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .E(n22012), 
            .D(n326[1]), .R(n22193));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(r_SM_Main_2__N_3383[2]), 
            .R(n35545));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i18592_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n26980));
    defparam i18592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_141_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_141_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_142_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_142_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut (.I0(n20583), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n20781));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n14), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(RX_N_10));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFFESR r_Clock_Count_1511__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), 
            .E(n21972), .D(n37[0]), .R(n22159));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 r_Clock_Count_1511_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n31674), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1511_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1511_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n31673), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1511_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1511_add_4_8 (.CI(n31673), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n31674));
    SB_LUT4 r_Clock_Count_1511_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n31672), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1511_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1511_add_4_7 (.CI(n31672), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n31673));
    SB_LUT4 r_Clock_Count_1511_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n31671), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1511_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1511_add_4_6 (.CI(n31671), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n31672));
    SB_LUT4 r_Clock_Count_1511_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n31670), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1511_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1511_add_4_5 (.CI(n31670), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n31671));
    SB_LUT4 r_Clock_Count_1511_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n31669), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1511_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1511_add_4_4 (.CI(n31669), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n31670));
    SB_LUT4 r_Clock_Count_1511_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n31668), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1511_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1511_add_4_3 (.CI(n31668), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n31669));
    SB_LUT4 r_Clock_Count_1511_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1511_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1511_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n31668));
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(n27558), .I1(r_SM_Main_2__N_3383[2]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n27846));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc7c7;
    SB_LUT4 i18_3_lut (.I0(n13), .I1(n27846), .I2(r_SM_Main[1]), .I3(GND_net), 
            .O(n14));   // verilog/uart_rx.v(30[17:26])
    defparam i18_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1589_2_lut (.I0(r_Bit_Index[1]), .I1(\r_Bit_Index[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i1589_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n27558));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i13790_3_lut (.I0(n22012), .I1(n27558), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n22193));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13790_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main_2__N_3383[2]), .I2(r_SM_Main[0]), 
            .I3(r_SM_Main[1]), .O(n22012));
    defparam i2_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i1596_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(\r_Bit_Index[0] ), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i1596_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i2_4_lut_adj_838 (.I0(r_SM_Main[2]), .I1(r_SM_Main_2__N_3383[2]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n20583));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i2_4_lut_adj_838.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_2_lut_adj_839 (.I0(\r_Bit_Index[0] ), .I1(n20583), .I2(GND_net), 
            .I3(GND_net), .O(n20776));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_839.LUT_INIT = 16'heeee;
    SB_LUT4 equal_144_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_144_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[5]), .I2(n36), 
            .I3(n5), .O(n25159));
    defparam i3_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_adj_840 (.I0(n25159), .I1(r_SM_Main[0]), .I2(GND_net), 
            .I3(GND_net), .O(n25166));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_adj_840.LUT_INIT = 16'hbbbb;
    SB_LUT4 i3_4_lut_adj_841 (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[4]), 
            .I2(r_Clock_Count[3]), .I3(r_Clock_Count[0]), .O(n5));
    defparam i3_4_lut_adj_841.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_842 (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[6]), 
            .I2(GND_net), .I3(GND_net), .O(n36));   // verilog/uart_rx.v(120[34:51])
    defparam i1_2_lut_adj_842.LUT_INIT = 16'heeee;
    SB_LUT4 i19164_4_lut (.I0(r_Clock_Count[2]), .I1(n36), .I2(r_Clock_Count[5]), 
            .I3(n5), .O(r_SM_Main_2__N_3383[2]));
    defparam i19164_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i13756_3_lut (.I0(n21972), .I1(r_SM_Main[2]), .I2(n8), .I3(GND_net), 
            .O(n22159));   // verilog/uart_rx.v(120[34:51])
    defparam i13756_3_lut.LUT_INIT = 16'h8a8a;
    SB_LUT4 i1_4_lut (.I0(r_Rx_Data), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(n25166), .O(n21972));   // verilog/uart_rx.v(30[17:26])
    defparam i1_4_lut.LUT_INIT = 16'h3331;
    SB_LUT4 i17_3_lut_4_lut_3_lut (.I0(r_SM_Main[0]), .I1(n25159), .I2(r_Rx_Data), 
            .I3(GND_net), .O(n13));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i17_3_lut_4_lut_3_lut.LUT_INIT = 16'h8d8d;
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n27922), 
            .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(\r_Bit_Index[0] ), .C(clk32MHz), .D(n22843));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .D(n35192));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n22847));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i19_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(n25159), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_3383[2]), .O(n8));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i19_3_lut_4_lut.LUT_INIT = 16'h08f8;
    SB_LUT4 i21_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_3383[2]), 
            .I3(r_SM_Main[0]), .O(n21911));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i21_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n21911), 
            .I3(rx_data_ready), .O(n35192));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 i30275_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n35545));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i30275_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n22308));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n22307));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n22306));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n22305));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n22304));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n22303));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n22302));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i29370_2_lut (.I0(r_SM_Main_2__N_3383[2]), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n39267));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i29370_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(n25166), .I1(n39267), 
            .I2(r_SM_Main[1]), .I3(r_Rx_Data), .O(n27922));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'h3035;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (encoder1_position, GND_net, clk32MHz, 
            data_o, n37217, reg_B, VCC_net, ENCODER1_A_c_1, ENCODER1_B_c_0, 
            n22849, n22320) /* synthesis syn_module_defined=1 */ ;
    output [23:0]encoder1_position;
    input GND_net;
    input clk32MHz;
    output [1:0]data_o;
    output n37217;
    output [1:0]reg_B;
    input VCC_net;
    input ENCODER1_A_c_1;
    input ENCODER1_B_c_0;
    input n22849;
    input n22320;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n2992;
    
    wire n2969, n30969, n30968, n30967, n30966, count_enable, B_delayed, 
        A_delayed, n30965, n30964, n30963, n30962, n30961, n30960, 
        n30959, n30958, n30957, n30956, n30955, n30954, n30953, 
        n30952, n30951, n30950, n30949, n30948, n30947, count_direction, 
        n30946;
    
    SB_LUT4 add_687_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2969), 
            .I3(n30969), .O(n2992[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_687_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2969), 
            .I3(n30968), .O(n2992[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_24 (.CI(n30968), .I0(encoder1_position[22]), .I1(n2969), 
            .CO(n30969));
    SB_LUT4 add_687_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2969), 
            .I3(n30967), .O(n2992[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_23 (.CI(n30967), .I0(encoder1_position[21]), .I1(n2969), 
            .CO(n30968));
    SB_LUT4 add_687_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2969), 
            .I3(n30966), .O(n2992[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_22_lut.LUT_INIT = 16'hC33C;
    SB_DFFE count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[0]));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_CARRY add_687_22 (.CI(n30966), .I0(encoder1_position[20]), .I1(n2969), 
            .CO(n30967));
    SB_LUT4 add_687_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2969), 
            .I3(n30965), .O(n2992[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_21 (.CI(n30965), .I0(encoder1_position[19]), .I1(n2969), 
            .CO(n30966));
    SB_LUT4 add_687_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2969), 
            .I3(n30964), .O(n2992[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_20 (.CI(n30964), .I0(encoder1_position[18]), .I1(n2969), 
            .CO(n30965));
    SB_LUT4 add_687_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2969), 
            .I3(n30963), .O(n2992[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_19 (.CI(n30963), .I0(encoder1_position[17]), .I1(n2969), 
            .CO(n30964));
    SB_LUT4 add_687_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2969), 
            .I3(n30962), .O(n2992[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_18_lut.LUT_INIT = 16'hC33C;
    SB_DFFE count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[23]));   // quad.v(35[10] 41[6])
    SB_CARRY add_687_18 (.CI(n30962), .I0(encoder1_position[16]), .I1(n2969), 
            .CO(n30963));
    SB_LUT4 add_687_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2969), 
            .I3(n30961), .O(n2992[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_17 (.CI(n30961), .I0(encoder1_position[15]), .I1(n2969), 
            .CO(n30962));
    SB_LUT4 add_687_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2969), 
            .I3(n30960), .O(n2992[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_16_lut.LUT_INIT = 16'hC33C;
    SB_DFFE count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[22]));   // quad.v(35[10] 41[6])
    SB_CARRY add_687_16 (.CI(n30960), .I0(encoder1_position[14]), .I1(n2969), 
            .CO(n30961));
    SB_LUT4 add_687_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2969), 
            .I3(n30959), .O(n2992[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_15 (.CI(n30959), .I0(encoder1_position[13]), .I1(n2969), 
            .CO(n30960));
    SB_LUT4 add_687_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2969), 
            .I3(n30958), .O(n2992[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_14 (.CI(n30958), .I0(encoder1_position[12]), .I1(n2969), 
            .CO(n30959));
    SB_LUT4 add_687_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2969), 
            .I3(n30957), .O(n2992[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_13 (.CI(n30957), .I0(encoder1_position[11]), .I1(n2969), 
            .CO(n30958));
    SB_LUT4 add_687_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2969), 
            .I3(n30956), .O(n2992[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_12 (.CI(n30956), .I0(encoder1_position[10]), .I1(n2969), 
            .CO(n30957));
    SB_DFFE count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[21]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[20]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[19]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[18]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[17]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[16]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[15]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[14]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[13]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[12]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[11]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[10]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[9]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[8]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[7]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[6]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[5]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[4]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[3]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[2]));   // quad.v(35[10] 41[6])
    SB_DFFE count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .E(count_enable), 
            .D(n2992[1]));   // quad.v(35[10] 41[6])
    SB_LUT4 add_687_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2969), 
            .I3(n30955), .O(n2992[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_11 (.CI(n30955), .I0(encoder1_position[9]), .I1(n2969), 
            .CO(n30956));
    SB_LUT4 add_687_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2969), 
            .I3(n30954), .O(n2992[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_10 (.CI(n30954), .I0(encoder1_position[8]), .I1(n2969), 
            .CO(n30955));
    SB_LUT4 add_687_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2969), 
            .I3(n30953), .O(n2992[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_9 (.CI(n30953), .I0(encoder1_position[7]), .I1(n2969), 
            .CO(n30954));
    SB_LUT4 add_687_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2969), 
            .I3(n30952), .O(n2992[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_8 (.CI(n30952), .I0(encoder1_position[6]), .I1(n2969), 
            .CO(n30953));
    SB_LUT4 add_687_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2969), 
            .I3(n30951), .O(n2992[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_7 (.CI(n30951), .I0(encoder1_position[5]), .I1(n2969), 
            .CO(n30952));
    SB_LUT4 add_687_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2969), 
            .I3(n30950), .O(n2992[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_6 (.CI(n30950), .I0(encoder1_position[4]), .I1(n2969), 
            .CO(n30951));
    SB_LUT4 add_687_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2969), 
            .I3(n30949), .O(n2992[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_5 (.CI(n30949), .I0(encoder1_position[3]), .I1(n2969), 
            .CO(n30950));
    SB_LUT4 add_687_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2969), 
            .I3(n30948), .O(n2992[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_4 (.CI(n30948), .I0(encoder1_position[2]), .I1(n2969), 
            .CO(n30949));
    SB_LUT4 add_687_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2969), 
            .I3(n30947), .O(n2992[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_3 (.CI(n30947), .I0(encoder1_position[1]), .I1(n2969), 
            .CO(n30948));
    SB_LUT4 add_687_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n30946), .O(n2992[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_687_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_687_2 (.CI(n30946), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n30947));
    SB_CARRY add_687_1 (.CI(GND_net), .I0(n2969), .I1(n2969), .CO(n30946));
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1142_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2969));   // quad.v(37[5] 40[8])
    defparam i1142_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,100)  debounce (.GND_net(GND_net), .n37217(n37217), 
            .reg_B({reg_B}), .VCC_net(VCC_net), .ENCODER1_A_c_1(ENCODER1_A_c_1), 
            .clk32MHz(clk32MHz), .ENCODER1_B_c_0(ENCODER1_B_c_0), .n22849(n22849), 
            .data_o({data_o}), .n22320(n22320));   // quad.v(15[37] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,100) 
//

module \grp_debouncer(2,100)  (GND_net, n37217, reg_B, VCC_net, ENCODER1_A_c_1, 
            clk32MHz, ENCODER1_B_c_0, n22849, data_o, n22320);
    input GND_net;
    output n37217;
    output [1:0]reg_B;
    input VCC_net;
    input ENCODER1_A_c_1;
    input clk32MHz;
    input ENCODER1_B_c_0;
    input n22849;
    output [1:0]data_o;
    input n22320;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire n31692;
    wire [6:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire n31693;
    wire [6:0]n33;
    
    wire n31691, n12;
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_6__N_3697, n31690, n31689, n31694;
    
    SB_CARRY cnt_reg_1515_add_4_6 (.CI(n31692), .I0(GND_net), .I1(cnt_reg[4]), 
            .CO(n31693));
    SB_LUT4 cnt_reg_1515_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[3]), 
            .I3(n31691), .O(n33[3])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1515_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1515_add_4_5 (.CI(n31691), .I0(GND_net), .I1(cnt_reg[3]), 
            .CO(n31692));
    SB_LUT4 i5_4_lut (.I0(cnt_reg[5]), .I1(cnt_reg[3]), .I2(cnt_reg[6]), 
            .I3(cnt_reg[4]), .O(n12));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(170[42:59])
    defparam i5_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i6_4_lut (.I0(cnt_reg[1]), .I1(n12), .I2(cnt_reg[2]), .I3(cnt_reg[0]), 
            .O(n37217));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(170[42:59])
    defparam i6_4_lut.LUT_INIT = 16'hffef;
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n37217), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_6__N_3697));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 cnt_reg_1515_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[2]), 
            .I3(n31690), .O(n33[2])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1515_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1515_add_4_4 (.CI(n31690), .I0(GND_net), .I1(cnt_reg[2]), 
            .CO(n31691));
    SB_LUT4 cnt_reg_1515_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[1]), 
            .I3(n31689), .O(n33[1])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1515_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1515_add_4_3 (.CI(n31689), .I0(GND_net), .I1(cnt_reg[1]), 
            .CO(n31690));
    SB_LUT4 cnt_reg_1515_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[0]), 
            .I3(VCC_net), .O(n33[0])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1515_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1515_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(cnt_reg[0]), 
            .CO(n31689));
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(ENCODER1_A_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1515__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n33[0]), 
            .R(cnt_next_6__N_3697));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(ENCODER1_B_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n22849));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n22320));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1515__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n33[1]), 
            .R(cnt_next_6__N_3697));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1515__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n33[2]), 
            .R(cnt_next_6__N_3697));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1515__i3 (.Q(cnt_reg[3]), .C(clk32MHz), .D(n33[3]), 
            .R(cnt_next_6__N_3697));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1515__i4 (.Q(cnt_reg[4]), .C(clk32MHz), .D(n33[4]), 
            .R(cnt_next_6__N_3697));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1515__i5 (.Q(cnt_reg[5]), .C(clk32MHz), .D(n33[5]), 
            .R(cnt_next_6__N_3697));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1515__i6 (.Q(cnt_reg[6]), .C(clk32MHz), .D(n33[6]), 
            .R(cnt_next_6__N_3697));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 cnt_reg_1515_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[6]), 
            .I3(n31694), .O(n33[6])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1515_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 cnt_reg_1515_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[5]), 
            .I3(n31693), .O(n33[5])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1515_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY cnt_reg_1515_add_4_7 (.CI(n31693), .I0(GND_net), .I1(cnt_reg[5]), 
            .CO(n31694));
    SB_LUT4 cnt_reg_1515_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(cnt_reg[4]), 
            .I3(n31692), .O(n33[4])) /* synthesis syn_instantiated=1 */ ;
    defparam cnt_reg_1515_add_4_6_lut.LUT_INIT = 16'hC33C;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (n39932, VCC_net, INHA_c, clk32MHz, n20604, GND_net, 
            n20602, \pwm_counter[6] , \pwm_counter[8] , \pwm_counter[7] , 
            \pwm_counter[13] , \pwm_counter[10] , \pwm_counter[9] , \pwm_counter[17] , 
            \pwm_counter[22] , \pwm_counter[14] , \pwm_counter[18] , \pwm_counter[21] , 
            \pwm_counter[16] , \pwm_counter[12] , \pwm_counter[15] , \pwm_counter[19] , 
            \pwm_counter[11] , \pwm_counter[20] , \pwm_counter[31] , \pwm_counter[0] , 
            \pwm_counter[5] , \pwm_counter[4] , \pwm_counter[3] , \pwm_counter[2] , 
            \pwm_counter[1] ) /* synthesis syn_module_defined=1 */ ;
    input n39932;
    input VCC_net;
    output INHA_c;
    input clk32MHz;
    input n20604;
    input GND_net;
    output n20602;
    output \pwm_counter[6] ;
    output \pwm_counter[8] ;
    output \pwm_counter[7] ;
    output \pwm_counter[13] ;
    output \pwm_counter[10] ;
    output \pwm_counter[9] ;
    output \pwm_counter[17] ;
    output \pwm_counter[22] ;
    output \pwm_counter[14] ;
    output \pwm_counter[18] ;
    output \pwm_counter[21] ;
    output \pwm_counter[16] ;
    output \pwm_counter[12] ;
    output \pwm_counter[15] ;
    output \pwm_counter[19] ;
    output \pwm_counter[11] ;
    output \pwm_counter[20] ;
    output \pwm_counter[31] ;
    output \pwm_counter[0] ;
    output \pwm_counter[5] ;
    output \pwm_counter[4] ;
    output \pwm_counter[3] ;
    output \pwm_counter[2] ;
    output \pwm_counter[1] ;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [31:0]pwm_counter;   // verilog/pwm.v(11[9:20])
    
    wire n10, n14, n37494, n18, n24, n22, n26, n21, pwm_counter_31__N_652;
    wire [31:0]n133;
    
    wire n31667, n31666, n31665, n31664, n31663, n31662, n31661, 
        n31660, n31659, n31658, n31657, n31656, n31655, n31654, 
        n31653, n31652, n31651, n31650, n31649, n31648, n31647, 
        n31646, n31645, n31644, n31643, n31642, n31641, n31640, 
        n31639, n31638, n31637;
    
    SB_DFFESR pwm_out_12 (.Q(INHA_c), .C(clk32MHz), .E(VCC_net), .D(n39932), 
            .R(n20604));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 i2_2_lut (.I0(pwm_counter[27]), .I1(pwm_counter[28]), .I2(GND_net), 
            .I3(GND_net), .O(n10));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut (.I0(pwm_counter[23]), .I1(pwm_counter[29]), .I2(pwm_counter[25]), 
            .I3(pwm_counter[26]), .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(pwm_counter[30]), .I1(n14), .I2(n10), .I3(pwm_counter[24]), 
            .O(n20602));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(\pwm_counter[6] ), .I1(\pwm_counter[8] ), .I2(\pwm_counter[7] ), 
            .I3(GND_net), .O(n37494));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(n37494), .I1(\pwm_counter[13] ), .I2(\pwm_counter[10] ), 
            .I3(\pwm_counter[9] ), .O(n18));
    defparam i4_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i10_4_lut (.I0(\pwm_counter[17] ), .I1(\pwm_counter[22] ), .I2(\pwm_counter[14] ), 
            .I3(\pwm_counter[18] ), .O(n24));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(\pwm_counter[21] ), .I1(n20602), .I2(\pwm_counter[16] ), 
            .I3(\pwm_counter[12] ), .O(n22));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(\pwm_counter[15] ), .I1(n24), .I2(n18), .I3(\pwm_counter[19] ), 
            .O(n26));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_2_lut (.I0(\pwm_counter[11] ), .I1(\pwm_counter[20] ), .I2(GND_net), 
            .I3(GND_net), .O(n21));
    defparam i7_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i18764_4_lut (.I0(n21), .I1(\pwm_counter[31] ), .I2(n26), 
            .I3(n22), .O(pwm_counter_31__N_652));   // verilog/pwm.v(18[8:40])
    defparam i18764_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 pwm_counter_1509_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[31] ), 
            .I3(n31667), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_counter_1509_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[30]), 
            .I3(n31666), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_32 (.CI(n31666), .I0(GND_net), .I1(pwm_counter[30]), 
            .CO(n31667));
    SB_LUT4 pwm_counter_1509_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[29]), 
            .I3(n31665), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_31 (.CI(n31665), .I0(GND_net), .I1(pwm_counter[29]), 
            .CO(n31666));
    SB_LUT4 pwm_counter_1509_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[28]), 
            .I3(n31664), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_30 (.CI(n31664), .I0(GND_net), .I1(pwm_counter[28]), 
            .CO(n31665));
    SB_LUT4 pwm_counter_1509_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[27]), 
            .I3(n31663), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_29 (.CI(n31663), .I0(GND_net), .I1(pwm_counter[27]), 
            .CO(n31664));
    SB_LUT4 pwm_counter_1509_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[26]), 
            .I3(n31662), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_28 (.CI(n31662), .I0(GND_net), .I1(pwm_counter[26]), 
            .CO(n31663));
    SB_LUT4 pwm_counter_1509_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[25]), 
            .I3(n31661), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_27 (.CI(n31661), .I0(GND_net), .I1(pwm_counter[25]), 
            .CO(n31662));
    SB_LUT4 pwm_counter_1509_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[24]), 
            .I3(n31660), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_26 (.CI(n31660), .I0(GND_net), .I1(pwm_counter[24]), 
            .CO(n31661));
    SB_LUT4 pwm_counter_1509_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n31659), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_25 (.CI(n31659), .I0(GND_net), .I1(pwm_counter[23]), 
            .CO(n31660));
    SB_LUT4 pwm_counter_1509_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[22] ), 
            .I3(n31658), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_24 (.CI(n31658), .I0(GND_net), .I1(\pwm_counter[22] ), 
            .CO(n31659));
    SB_LUT4 pwm_counter_1509_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[21] ), 
            .I3(n31657), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_23 (.CI(n31657), .I0(GND_net), .I1(\pwm_counter[21] ), 
            .CO(n31658));
    SB_LUT4 pwm_counter_1509_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[20] ), 
            .I3(n31656), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_22 (.CI(n31656), .I0(GND_net), .I1(\pwm_counter[20] ), 
            .CO(n31657));
    SB_LUT4 pwm_counter_1509_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[19] ), 
            .I3(n31655), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_21 (.CI(n31655), .I0(GND_net), .I1(\pwm_counter[19] ), 
            .CO(n31656));
    SB_LUT4 pwm_counter_1509_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[18] ), 
            .I3(n31654), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_20 (.CI(n31654), .I0(GND_net), .I1(\pwm_counter[18] ), 
            .CO(n31655));
    SB_LUT4 pwm_counter_1509_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[17] ), 
            .I3(n31653), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_19 (.CI(n31653), .I0(GND_net), .I1(\pwm_counter[17] ), 
            .CO(n31654));
    SB_LUT4 pwm_counter_1509_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[16] ), 
            .I3(n31652), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_18 (.CI(n31652), .I0(GND_net), .I1(\pwm_counter[16] ), 
            .CO(n31653));
    SB_LUT4 pwm_counter_1509_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[15] ), 
            .I3(n31651), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_17 (.CI(n31651), .I0(GND_net), .I1(\pwm_counter[15] ), 
            .CO(n31652));
    SB_LUT4 pwm_counter_1509_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[14] ), 
            .I3(n31650), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_16 (.CI(n31650), .I0(GND_net), .I1(\pwm_counter[14] ), 
            .CO(n31651));
    SB_LUT4 pwm_counter_1509_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[13] ), 
            .I3(n31649), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_15 (.CI(n31649), .I0(GND_net), .I1(\pwm_counter[13] ), 
            .CO(n31650));
    SB_LUT4 pwm_counter_1509_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[12] ), 
            .I3(n31648), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_14 (.CI(n31648), .I0(GND_net), .I1(\pwm_counter[12] ), 
            .CO(n31649));
    SB_LUT4 pwm_counter_1509_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[11] ), 
            .I3(n31647), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_13 (.CI(n31647), .I0(GND_net), .I1(\pwm_counter[11] ), 
            .CO(n31648));
    SB_LUT4 pwm_counter_1509_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[10] ), 
            .I3(n31646), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_12 (.CI(n31646), .I0(GND_net), .I1(\pwm_counter[10] ), 
            .CO(n31647));
    SB_LUT4 pwm_counter_1509_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[9] ), 
            .I3(n31645), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_11 (.CI(n31645), .I0(GND_net), .I1(\pwm_counter[9] ), 
            .CO(n31646));
    SB_LUT4 pwm_counter_1509_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[8] ), 
            .I3(n31644), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_10 (.CI(n31644), .I0(GND_net), .I1(\pwm_counter[8] ), 
            .CO(n31645));
    SB_DFFSR pwm_counter_1509__i0 (.Q(\pwm_counter[0] ), .C(clk32MHz), .D(n133[0]), 
            .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_LUT4 pwm_counter_1509_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[7] ), 
            .I3(n31643), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_9 (.CI(n31643), .I0(GND_net), .I1(\pwm_counter[7] ), 
            .CO(n31644));
    SB_LUT4 pwm_counter_1509_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[6] ), 
            .I3(n31642), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_8 (.CI(n31642), .I0(GND_net), .I1(\pwm_counter[6] ), 
            .CO(n31643));
    SB_LUT4 pwm_counter_1509_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[5] ), 
            .I3(n31641), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_7 (.CI(n31641), .I0(GND_net), .I1(\pwm_counter[5] ), 
            .CO(n31642));
    SB_LUT4 pwm_counter_1509_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[4] ), 
            .I3(n31640), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_6 (.CI(n31640), .I0(GND_net), .I1(\pwm_counter[4] ), 
            .CO(n31641));
    SB_LUT4 pwm_counter_1509_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[3] ), 
            .I3(n31639), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_5 (.CI(n31639), .I0(GND_net), .I1(\pwm_counter[3] ), 
            .CO(n31640));
    SB_LUT4 pwm_counter_1509_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[2] ), 
            .I3(n31638), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_4 (.CI(n31638), .I0(GND_net), .I1(\pwm_counter[2] ), 
            .CO(n31639));
    SB_LUT4 pwm_counter_1509_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[1] ), 
            .I3(n31637), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_3 (.CI(n31637), .I0(GND_net), .I1(\pwm_counter[1] ), 
            .CO(n31638));
    SB_LUT4 pwm_counter_1509_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\pwm_counter[0] ), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1509_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1509_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\pwm_counter[0] ), 
            .CO(n31637));
    SB_DFFSR pwm_counter_1509__i1 (.Q(\pwm_counter[1] ), .C(clk32MHz), .D(n133[1]), 
            .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i2 (.Q(\pwm_counter[2] ), .C(clk32MHz), .D(n133[2]), 
            .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i3 (.Q(\pwm_counter[3] ), .C(clk32MHz), .D(n133[3]), 
            .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i4 (.Q(\pwm_counter[4] ), .C(clk32MHz), .D(n133[4]), 
            .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i5 (.Q(\pwm_counter[5] ), .C(clk32MHz), .D(n133[5]), 
            .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i6 (.Q(\pwm_counter[6] ), .C(clk32MHz), .D(n133[6]), 
            .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i7 (.Q(\pwm_counter[7] ), .C(clk32MHz), .D(n133[7]), 
            .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i8 (.Q(\pwm_counter[8] ), .C(clk32MHz), .D(n133[8]), 
            .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i9 (.Q(\pwm_counter[9] ), .C(clk32MHz), .D(n133[9]), 
            .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i10 (.Q(\pwm_counter[10] ), .C(clk32MHz), 
            .D(n133[10]), .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i11 (.Q(\pwm_counter[11] ), .C(clk32MHz), 
            .D(n133[11]), .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i12 (.Q(\pwm_counter[12] ), .C(clk32MHz), 
            .D(n133[12]), .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i13 (.Q(\pwm_counter[13] ), .C(clk32MHz), 
            .D(n133[13]), .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i14 (.Q(\pwm_counter[14] ), .C(clk32MHz), 
            .D(n133[14]), .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i15 (.Q(\pwm_counter[15] ), .C(clk32MHz), 
            .D(n133[15]), .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i16 (.Q(\pwm_counter[16] ), .C(clk32MHz), 
            .D(n133[16]), .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i17 (.Q(\pwm_counter[17] ), .C(clk32MHz), 
            .D(n133[17]), .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i18 (.Q(\pwm_counter[18] ), .C(clk32MHz), 
            .D(n133[18]), .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i19 (.Q(\pwm_counter[19] ), .C(clk32MHz), 
            .D(n133[19]), .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i20 (.Q(\pwm_counter[20] ), .C(clk32MHz), 
            .D(n133[20]), .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i21 (.Q(\pwm_counter[21] ), .C(clk32MHz), 
            .D(n133[21]), .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i22 (.Q(\pwm_counter[22] ), .C(clk32MHz), 
            .D(n133[22]), .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n133[23]), 
            .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i24 (.Q(pwm_counter[24]), .C(clk32MHz), .D(n133[24]), 
            .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i25 (.Q(pwm_counter[25]), .C(clk32MHz), .D(n133[25]), 
            .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i26 (.Q(pwm_counter[26]), .C(clk32MHz), .D(n133[26]), 
            .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i27 (.Q(pwm_counter[27]), .C(clk32MHz), .D(n133[27]), 
            .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i28 (.Q(pwm_counter[28]), .C(clk32MHz), .D(n133[28]), 
            .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i29 (.Q(pwm_counter[29]), .C(clk32MHz), .D(n133[29]), 
            .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i30 (.Q(pwm_counter[30]), .C(clk32MHz), .D(n133[30]), 
            .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1509__i31 (.Q(\pwm_counter[31] ), .C(clk32MHz), 
            .D(n133[31]), .R(pwm_counter_31__N_652));   // verilog/pwm.v(17[20:33])
    
endmodule
