// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Sun Oct 27 08:59:01 2019
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, PIN_1, PIN_2, PIN_3, PIN_4, 
            PIN_5, PIN_6, PIN_7, PIN_8, PIN_9, PIN_10, PIN_11, 
            PIN_12, PIN_13, PIN_14, PIN_15, PIN_16, PIN_17, PIN_18, 
            PIN_19, PIN_20, PIN_21, PIN_22, PIN_23, PIN_24) /* synthesis syn_preserve=0, syn_noprune=0, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input PIN_1 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(6[9:14])
    input PIN_2 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(7[9:14])
    inout PIN_3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(8[9:14])
    inout PIN_4 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(9[9:14])
    inout PIN_5 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input PIN_6 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input PIN_7 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    output PIN_8 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(13[9:14])
    inout PIN_9 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(14[9:14])
    inout PIN_10 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(15[9:15])
    inout PIN_11 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[9:15])
    inout PIN_12 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(17[9:15])
    input PIN_13 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(18[9:15])
    input PIN_14 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(19[9:15])
    input PIN_15 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(20[9:15])
    input PIN_16 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(21[9:15])
    input PIN_17 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:15])
    input PIN_18 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(23[9:15])
    output PIN_19 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(24[9:15])
    output PIN_20 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(25[9:15])
    output PIN_21 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(26[9:15])
    output PIN_22 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(27[9:15])
    output PIN_23 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(28[9:15])
    output PIN_24 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(29[9:15])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire LED_c /* synthesis SET_AS_NETWORK=LED_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(4[10:13])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire GND_net, VCC_net, PIN_1_c_1, PIN_2_c_0, PIN_6_c_0, PIN_7_c_1, 
        PIN_8_c, PIN_13_c, PIN_19_c_0, PIN_20_c, PIN_21_c, PIN_22_c, 
        PIN_23_c;
    wire [31:0]communication_counter;   // verilog/TinyFPGA_B.v(42[9:30])
    
    wire n1253;
    wire [23:0]color;   // verilog/TinyFPGA_B.v(43[12:17])
    
    wire blink, hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(117[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(118[21:25])
    
    wire tx_o, tx_enable, ID0, ID1, ID2, n4;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(182[22:39])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(183[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(184[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(185[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(186[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(187[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(189[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(190[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(191[22:35])
    wire [23:0]gearBoxRatio;   // verilog/TinyFPGA_B.v(193[22:34])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(218[22:33])
    
    wire n30786;
    wire [7:0]color_23__N_164;
    
    wire n30944, n30943, n18602, n30619, n1155, n1154, n7, n38245, 
        n1153, n1152, n1151, blink_N_255;
    wire [22:0]pwm_setpoint_22__N_57;
    
    wire PIN_13_N_105;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    
    wire n1222;
    wire [31:0]motor_state_23__N_106;
    wire [24:0]displacement_23__N_229;
    wire [23:0]displacement_23__N_80;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire start, \neo_pixel_transmitter.done ;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n30618, n30942, n30617, n30785, n30784;
    wire [3:0]state_3__N_362;
    
    wire n30941, n19265, n30616, n19266, n19267, n30940, n19268, 
        n19269, n19272;
    wire [31:0]one_wire_N_513;
    
    wire n18, n16, n44557, n13, n30939, n30938, n30615, n30937, 
        n30783, n30614, n30782, n30936, n30781, n30780, n30935, 
        n30779, n12501, n45113, n14, n1257, n30934, n30778, n30777, 
        n43084, n10, n2889, n2888, n30933, n30932, n17272, n30931, 
        n45109, n45108, n2816, n22, n23, n34, n33, n1258, n30930, 
        n2887, n2886, n2817, n32, n2885, n2884, n2883, n2882, 
        n2881, n24, n17268, n21, n2819, n2818, n2880, n2879, 
        n2878, n2877, n43631, n2876, n2875, n2874, n2873, n2872, 
        n2871, n2870, n31, n2869, n2868, n2867, n2866, n2839, 
        n2838, n2837, n2836, n2835, n2834, n2833, n30, n30776, 
        n30775, n2832, n2831, n2830, n30774, n30929, n30928, n30927, 
        n30926, n30925, n30924, n17264, n17293, n30923, n1125, 
        n1124, n1123, n1122, n1121, n1120, n45095, n43625, n35929, 
        n2829, n2828, n2;
    wire [9:0]half_duty_new;   // vhdl/pwm.vhd(53[12:25])
    
    wire n30773, n3;
    wire [9:0]\half_duty[0] ;   // vhdl/pwm.vhd(55[11:20])
    
    wire n45089, n45110, n2827, n2826, n30772, n45085, n4_adj_4326, 
        n19201, n30922, n30921, n3_adj_4327, n4_adj_4328, n5, n6, 
        n7_adj_4329, n8, n9, n10_adj_4330, n11, n12, n13_adj_4331, 
        n14_adj_4332, n15, n16_adj_4333, n17, n18_adj_4334, n19, 
        n20, n21_adj_4335, n22_adj_4336, n23_adj_4337, n24_adj_4338, 
        n25, n17299, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(89[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(93[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(93[12:19])
    
    wire n30771, n30920;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(94[12:25])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(95[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(95[12:26])
    
    wire n43622;
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(95[12:26])
    
    wire tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(110[11:16])
    
    wire n43616, n393, n392, n391, n390, n389, n388, n387, n386, 
        n385, n384, n383, n382, n381, n380, n379, n378, n30770, 
        n30919, n4_adj_4339, n30918, n30917, n30916, n30769, n30915, 
        n30768, n30914, n30767, n30766, n30913, n30912, n13_adj_4340, 
        n17250, n30765, n30911, n30764, n45112, n43613, n30763, 
        n30762, n30761, n11_adj_4341, n45094, n44580, n2825, n44321, 
        n20_adj_4342, n19_adj_4343, n18_adj_4344, n45054, n45052, 
        n43601, n40, n45051, n45048, n39, n45046, n38, n30760, 
        n38270, n30910, n45045, n30909, n37, n30908, n740, n30759, 
        n30907, n6_adj_4345, n35, n30758, n30906, n30905, n30904, 
        n30757, n30903, n8_adj_4346, n34_adj_4347, n30756, n30755, 
        n30902, n30901, n30754, n30753, n30900, n30899, n45030, 
        n44997, n44325, n17244, n30898, n30897, n30752, n44981, 
        n44979, n30751, n30750, n27, n30749, n30748, n30896, n44975, 
        n17241, n30747, n30746, n30745, n38308, n30895, n30744, 
        n30743, n30742, n30894, n38279, n44971, n44965, n30741, 
        n17236, n30740, n17231, n30739, n30738, n43587, n30737, 
        n30736, n30735, n30734, n44955, n30893, n43583, n30892, 
        n43579, n30733, n30732, n30891, n30731, n30890, n30889, 
        n30730, n6_adj_4348, n30729, n30888, n30887, n30728, n4_adj_4349, 
        n17200, n30886, n30727, n30885, n30884, n17195, n43577, 
        n30726, n44934, n30883, n30725, n30882, n30881, n30724, 
        n17269, n30723, n10_adj_4350, n17202, n20874, n20896, n42, 
        n38295, n95, n2824, n2823, n1220, n41, n40_adj_4351, n2822, 
        n39_adj_4352, n2821, n30880, n30879, n37_adj_4353, n30722, 
        n36, n30721, n44912, n30570, n2857, n44909, n44908, n30569, 
        n30720, n30568, n30567, n38249, n17225, n30719, n29, n44901, 
        n44900, n30566, n30718, n30878, n26349, n1219, n30717, 
        n30565, n30454, n3761, n30716, n30715, n43564, n20639, 
        n43562, n24_adj_4354, n45043, n44883, n22_adj_4355, n30714, 
        n30877, n20_adj_4356, n30713, n30876, n16_adj_4357, n43552, 
        n30453, n44879, n43539, n43537, n44956, n44569, n44866, 
        n44857, n44855, n44853, n44851, n30712, n44849, n44847, 
        n44843, n44841, n44840, n30875, n1225, n30711, n1224, 
        n30710, n2820, n30452, n5_adj_4358, n15_adj_4359, n1223, 
        n30874, n30564, n19145, n19144, n19143, n19142, n43515, 
        n19141, n19140, n19139, n19138, n19137, n19136, n19135, 
        n19134, n19133, n19132, n19131, n19130, n19129, n19128, 
        n19127, n19126, n19125, n19124, n19123, n19122, n19121, 
        n19120, n19119, n19118, n19117, n19116, n19115, n19114, 
        n19113, n19112, n19111, n19110, n19109, n19108, n19107, 
        n19106, n19105, n19104, n19103, n19102, n19101, n19100, 
        n19099, n19098, n19097, n19096, n19095, n19094, n19093, 
        n19092, n19091, n19090, n19089, n19088, n19087, n19086, 
        n19085, n19084, n19083, n19082, n19081, n19080, n19079, 
        n19078, n19077, n19076, n19075, n19074, n19073, n19072, 
        n19071, n19070, n19069, n19068, n19067, n19066, n19065, 
        n19064, n19063, n19062, n19061, n19060, n19059, n19058, 
        n19057, n19056, n19055, n19054, n19053, n19052, n19051, 
        n19050, n19049, n19048, n19047, n19046, n19045, n19044, 
        n19043, n19042, n19041, n19040, n19039, n19038, n19037, 
        n19036, n19035, n19034, n19033, n19032, n19031, n19030, 
        n19029, n19028, n19027, n19026, n19025, n19024, n19023, 
        n19022, n19021, n19020, n19019, n19018, n19017, n19014, 
        n19013, n19012, n19011, n19010, n19009, n19008, n19007, 
        n19006, n19005, n19004, n19003, n19002, n19001, n19000, 
        n18999, n18998, n18997, n18996, n18995, n18994, n18993, 
        n18992, n18991, n18990, n18989, n18988, n18987, n18986, 
        n18985, n18984, n18983, n18982, n18981, n18943, n18940, 
        n18939, n18938, n377, n376, n375, n374, n373, n372, 
        n371, n370, n369, n1085, n30563, n37368, n17311, n249, 
        n248, n224, n44825, n1058, n1057, n1056, n1055, n1054, 
        n1053, n1052, n44823, n44575, n44819, n44967, n1025, n1024, 
        n1023, n1022, n1021, n30562, n2664, n30709, n1111, n99, 
        n98, n97, n96, n95_adj_4360, n94, n93, n92, n91, n90, 
        n89, n88, n87, n86, n85, n84, n83, n82, n81, n80, 
        n43509, n17305, n30873, n30872, n44738, n43507, n43505, 
        n18584, n30708, n30451, n44347, n30871, n4682, n4681, 
        n4680, n4679, n4678, n4677, n4676, n4675, n4674, n4673, 
        n4672, n4671, n4670, n4669, n4668, n4667, n4666, n4665, 
        n4664, n4663, n4662, n4661, n4660, n4659, n30450, n30707, 
        n4926, n4754, n1254, n15_adj_4361, n19271, n30706, n23_adj_4362, 
        n15_adj_4363, n25_adj_4364, n4_adj_4365, n12_adj_4366, n15_adj_4367, 
        n30705, n30561, n15_adj_4368, n8_adj_4369, n9_adj_4370, n19270, 
        n6899, quadA_debounced, quadB_debounced, count_enable, n6898, 
        n1252, n79, n78, n77, n75, n74, n73, n72, n71, n70, 
        n69, n68, n67, n66, n65, n64, n63, n62, n61, n60, 
        n59, n58, n57, n56, n55, n3_adj_4371, n1221, n1105, 
        quadA_debounced_adj_4372, quadB_debounced_adj_4373, count_enable_adj_4374, 
        n6897, n13_adj_4375, n54, n53, n17199, n30870, n44704, 
        n44810, n33_adj_4376, n32_adj_4377, n31_adj_4378, n30_adj_4379, 
        n29_adj_4380, n28, r_Rx_Data;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n6896, n6895, n44700, n27_adj_4381, n30704, n17189, n11_adj_4382, 
        n26, n35915;
    wire [2:0]r_SM_Main_adj_5046;   // verilog/uart_tx.v(31[16:25])
    wire [2:0]r_SM_Main_2__N_3320;
    
    wire n25_adj_4385, n30869, n30868, n24_adj_4386, n14536, n30867, 
        n30866, n18898, n18897, n30703, n30702;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n44579;
    wire [1:0]reg_B_adj_5057;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n23_adj_4389, n22_adj_4390, n21_adj_4391, n20_adj_4392, n19_adj_4393, 
        n18_adj_4394, n17_adj_4395, n16_adj_4396, n15_adj_4397, n14_adj_4398, 
        n13_adj_4399, n12_adj_4400, n11_adj_4401, n10_adj_4402, n9_adj_4403, 
        n8_adj_4404, n7_adj_4405, n6_adj_4406, n5_adj_4407, n4_adj_4408, 
        n3_adj_4409, n44685, n44678, n30865, n30701, n17_adj_4410, 
        n17302, n16_adj_4411, n17308, n1250, n4_adj_4412, n1251, 
        n1283, n44587, n1256, n1255, n8_adj_4413, n9_adj_4414, n10_adj_4415, 
        n11_adj_4416, n12_adj_4417, n13_adj_4418, n14_adj_4419, n15_adj_4420, 
        n16_adj_4421, n17_adj_4422, n18_adj_4423, n19_adj_4424, n20_adj_4425, 
        n21_adj_4426, n22_adj_4427, n23_adj_4428, n24_adj_4429, n25_adj_4430, 
        n6_adj_4431, n7_adj_4432, n986, n510, n17284, n17287, n533, 
        n534, n558, n17290, n18896, n35917, n30700, n44658, n35937, 
        n44654, n45127, n30560, n958, n957, n956, n955, n954, 
        n953, n648, n649, n671, n672, n44576, n44650, n44648, 
        n44966, n783, n784, n785, n44644, n12168, n12167, n12166, 
        n12165, n806, n807, n30449, n914, n915, n916, n917, 
        n918, n938, n939, n27453, n30559, n855, n852, n6900, 
        n6901, n6911, n6922, n43406, n1043, n1044, n1045, n1046, 
        n1047, n1048, n30864, n30448, n1067, n1068, n30558, n30699, 
        n10_adj_4433, n6904, n6905, n6906, n6907, n6908, n6909, 
        n6910, n1169, n1170, n1171, n1172, n1173, n1174, n1175, 
        n1193, n1194, n6962, n6948, n6934, n6892, n6891, n6890, 
        n6889, n6888, n6887, n6914, n6915, n6916, n6917, n6918, 
        n6919, n6920, n6921, n45146, n44634, n1292, n1293, n1294, 
        n1295, n1296, n1297, n1298, n1299, n45149, n45152, n45155, 
        n45158, n3459, n3458, n3457, n3456, n3455, n3454, n3453, 
        n3452, n1316, n1317, n30557, n46559, n749, n748, n746, 
        n2_adj_4434, n6925, n6926, n6927, n6928, n6929, n6930, 
        n6931, n6932, n6933, n30698, n1412, n1413, n1414, n1415, 
        n1416, n1417, n1418, n1419, n1420, n1436, n1437, n43390, 
        n30863, n30862, n12_adj_4435, n30697, n11_adj_4436, n6938, 
        n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, 
        n6947, n44583, n6965, n6966, n44627, n1529, n1530, n1531, 
        n1532, n1533, n1534, n1535, n1536, n1537, n1538, n6993, 
        n6992, n6991, n6990, n6989, n6988, n6987, n6986, n6985, 
        n6984, n6983, n6982, n6981, n6980, n1553, n1554, n3358, 
        n3357, n3356, n3355, n3354, n3353, n3351, n8_adj_4437, 
        n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, 
        n6959, n6960, n6961, n3337, n3340, n3342, n3344, n3346, 
        n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, 
        n1651, n1652, n1653, n3330, n3325, n3324, n1667, n1668, 
        n43384, n3322, n3321, n3320, n3319, n3318, n3317, n3316, 
        n3315, n3314, n3313, n3312, n3311, n30447, n6967, n6968, 
        n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, 
        n6977, n3300, n3301, n3302, n3303, n3304, n3305, n3306, 
        n3307, n3308, n3309, n3310, n30861, n1754, n1755, n1756, 
        n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, 
        n1765, n3299, n3298, n7013, n30446, n1778, n1779, n7039, 
        n7038, n7037, n7036, n7035, n7034, n7033, n7032, n7031, 
        n7062, n7061, n7051, n7052, n7053, n7054, n7055, n7056, 
        n7057, n7058, n7059, n7060, n1862, n1863, n1864, n1865, 
        n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, 
        n1874, n7050, n3263, n3258, n3257, n3256, n3255, n3254, 
        n1886, n1887, n3252, n3251, n3250, n3249, n3248, n3247, 
        n3246, n3245, n3244, n3243, n6997, n6998, n6999, n7000, 
        n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, 
        n7009, n7010, n3234, n3235, n3236, n3237, n3238, n3239, 
        n3240, n3241, n3242, n11305, n1967, n1968, n1969, n1970, 
        n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, 
        n1979, n1980, n3233, n3232, n3231, n3230, n3225, n3224, 
        n1991, n1992, n3222, n3221, n3220, n3219, n3218, n3217, 
        n3216, n3215, n3214, n7014, n7015, n7016, n7017, n7018, 
        n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, 
        n7027, n7028, n3206, n3207, n3208, n3209, n3210, n3211, 
        n3212, n3213, n2069, n2070, n2071, n2072, n2073, n2074, 
        n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, 
        n2083, n3205, n3204, n3203, n3202, n3201, n3200, n3199, 
        n7137, n2093, n2094, n7041, n7042, n7043, n7044, n7045, 
        n7046, n7047, n11304, n2168, n2169, n2170, n2171, n2172, 
        n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, 
        n2181, n2182, n2183, n2192, n2193, n30860, n3164, n7063, 
        n7064, n7065, n7066, n7067, n11303, n7088, n11302, n7110, 
        n11301, n7133, n11300, n7182, n3158, n43777, n2264, n2265, 
        n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, 
        n2274, n2275, n2276, n2277, n2278, n2279, n2280, n3157, 
        n3156, n3155, n3154, n3153, n3152, n3151, n2288, n2289, 
        n32338, n3149, n3148, n3147, n3146, n3145, n3144, n7070, 
        n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, 
        n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, 
        n7087, n3139, n3140, n3141, n3142, n3143, n2357, n2358, 
        n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, 
        n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, 
        n3138, n3137, n3136, n3135, n3134, n3133, n2381, n2382, 
        n6_adj_4438, n32337, n32336, n3131, n32335, n30859, n7091, 
        n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, 
        n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, 
        n7108, n7109, n3123, n3124, n3125, n2447, n2448, n2449, 
        n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, 
        n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, 
        n3122, n3121, n3120, n3119, n3118, n2471, n2472, n30445, 
        n32334, n30858, n3116, n3115, n3114, n3113, n7113, n7114, 
        n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, 
        n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, 
        n7131, n7132, n3110, n3111, n3112, n2534, n2535, n2536, 
        n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, 
        n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, 
        n2553, n3109, n3108, n3107, n3106, n2558, n2559, n3104, 
        n3103, n3102, n32333, n7138, n7139, n7140, n7141, n7142, 
        n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, 
        n7151, n7152, n7153, n7154, n7155, n7156, n7157, n32332, 
        n3100, n3101, n2618, n2619, n2620, n2621, n2622, n2623, 
        n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, 
        n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2642, 
        n2643, n7160, n7161, n7162, n7163, n7164, n7165, n7166, 
        n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, 
        n7175, n7176, n7177, n7178, n7179, n7180, n7181, n32331, 
        n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, 
        n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, 
        n2715, n2716, n2717, n2718, n2719, n2720, n2723, n2724, 
        n2777, n2798, n2799, n2801, n2802, n32330, n32329, n30696, 
        n30857, n18886, n32328, n18885, n18884, n18883, n18882, 
        n18881, n32327, n18880, n30856, n18879, n30855, n18878, 
        n18877, n18876, n18875, n18874, n18873, n18872, n18871, 
        n32326, n18870, n30854, n18869, n18868, n18867, n18866, 
        n18865, n18864, n32325, n18863, n18862, n18861, n32324, 
        n3065, n32323, n18860, n31448, n31447, n3058, n31446, 
        n31445, n3057, n3056, n31444, n3055, n3054, n3053, n3052, 
        n31443, n31442, n3051, n3050, n31441, n3049, n3048, n3047, 
        n38273, n31440, n31439, n31438, n31437, n31436, n31435, 
        n31434, n31433, n31432, n31431, n31430, n31429, n3046, 
        n3045, n3044, n3043, n3042, n3041, n3040, n3039, n31428, 
        n3038, n3037, n3036, n3035, n3034, n31427, n3033, n3032, 
        n31426, n31425, n31424, n31423, n31422, n31421, n31420, 
        n31419, n31418, n31417, n19450, n19449, n19448, n19447, 
        n19446, n19445, n19444, n19443, n19442, n19441, n31416, 
        n3025, n3024, n31415, n3023, n3022, n3021, n3020, n31414, 
        n3019, n31413, n3018, n3017, n31412, n3016, n31411, n3015, 
        n3014, n19440, n19439, n19438, n19437, n19436, n19435, 
        n19434, n19433, n19432, n19431, n19430, n19429, n19428, 
        n19427, n19426, n19425, n19424, n19423, n19422, n19421, 
        n19420, n19419, n31410, n35909, n19414, n35911, n63_adj_4439, 
        n3013, n3012, n35913, n3011, n3010, n3009, n3008, n19406, 
        n3007, n31409, n3006, n3005, n3004, n3003, n19401, n3002, 
        n19400, n3001, n19399, n19398, n19397, n19396, n19395, 
        n19394, n31408, n19393, n19392, n19391, n19390, n19389, 
        n19388, n31407, n19387, n19386, n19385, n19384, n19383, 
        n19382, n19381, n18859, n5_adj_4440, n19380, n19379, n19377, 
        n1184, n19376, n19375, n19374, n19373, n19372, n19371, 
        n19370, n19369, n19368, n2966, n19367, n31406, n19366, 
        n44353, n19365, n19364, n31405, n19363, n19362, n31404, 
        n19361, n31403, n19360, n2958, n19359, n2957, n19358, 
        n2956, n19357, n2955, n19356, n2954, n19355, n2953, n2952, 
        n2951, n2950, n2949, n2948, n17211, n2947, n2946, n2945, 
        n2944, n2943, n2942, n31402, n2941, n2940, n2939, n2938, 
        n2937, n2936, n2935, n2934, n2933, n31401, n2925, n2924, 
        n2923, n2922, n2921, n2920, n2919, n2918, n2917, n2916, 
        n2915, n2914, n31400, n2913, n2912, n2911, n2910, n38338, 
        n2909, n2908, n2907, n2906, n2905, n2904, n2903, n2902, 
        n43334, n18858, n18857, n18856, n18855, n2867_adj_4441, 
        n31399, n2858, n2857_adj_4442, n2856, n2855, n2854, n2853, 
        n2852, n2851, n2850, n2849, n2848, n18467, n31398, n31397, 
        n44676, n31396, n44671, n44970, n31395, n44859, n35925, 
        n43327, n32322, n31394, n35927, n18830, n32321, n18829, 
        n31393, n35931, n18816, n32320, n18815, n31392, n18814, 
        n35933, n32319, n31391, n18810, n35935, n32318, n18806, 
        n18805, n18804, n18802, n32317, n31390, n18798, n18793, 
        n35943, n32316, n31389, n18786, n32315, n18785, n31388, 
        n18784, n18783, n18782, n18781, n18780, n18777, n30853, 
        n32314, n30852, n31387, n30851, n30850, n18767, n32313, 
        n18765, n31386, n18764, n32312, n18762, n31385, n18761, 
        n18759, n18758, n18756, n18755, n44369, n18753, n18752, 
        n32311, n18750, n31384, n18749, n32310, n18747, n31383, 
        n18746, n18744, n36985, n36987, n36989, n31382, n31381, 
        n31380, n31379, n31378, n31377, n30556, n32309, n4_adj_4443, 
        n32308, n13_adj_4444, n11_adj_4445, n31376, n32307, n31375, 
        n32306, n32305, n31374, n31373, n31372, n27365, n31371, 
        n30695, n18435, n31370, n32304, n30849, n6119, n43307, 
        n2847, n2846, n2845, n2844, n2843, n2842, n2841, n2840, 
        n38326, n2839_adj_4446, n2838_adj_4447, n2837_adj_4448, n2836_adj_4449, 
        n2835_adj_4450, n2834_adj_4451, n2825_adj_4452, n2824_adj_4453, 
        n18416, n2823_adj_4454, n2822_adj_4455, n2821_adj_4456, n2820_adj_4457, 
        n2819_adj_4458, n2818_adj_4459, n2817_adj_4460, n2816_adj_4461, 
        n2815, n2814, n2813, n2812, n2811, n2810, n2809, n2808, 
        n2807, n2806, n30848, n2805, n2804, n30847, n2803, n30846, 
        n18402, n30555, n30694, n30845, n30844, n2768, n31369, 
        n44593, n2758, n31368, n2757, n2756, n2755, n2754, n2753, 
        n2752, n2751, n2750, n2749, n2748, n2747, n2746, n2745, 
        n38243, n2744, n2743, n2742, n2741, n2740, n2739, n2738, 
        n2737, n2736, n2735, n2725, n2724_adj_4462, n2723_adj_4463, 
        n2722, n35949, n2721, n2720_adj_4464, n2719_adj_4465, n2718_adj_4466, 
        n2717_adj_4467, n2716_adj_4468, n2715_adj_4469, n2714_adj_4470, 
        n2713_adj_4471, n2712_adj_4472, n2711_adj_4473, n2710_adj_4474, 
        n2709_adj_4475, n2708_adj_4476, n2707_adj_4477, n2706_adj_4478, 
        n2705_adj_4479, n2704_adj_4480, n31367, n31366, n32303, n31365, 
        n31364, n31363, n1646_adj_4481, n1647_adj_4482, n1648_adj_4483, 
        n1649_adj_4484, n1650_adj_4485, n1651_adj_4486, n1652_adj_4487, 
        n1653_adj_4488, n1654, n1655, n1656, n1657, n1658, n31362, 
        n31361, n31360, n31359, n1679, n37376, n1714, n1715, n1716, 
        n1717, n1718, n1719, n1720, n31358, n1721, n1722, n1723, 
        n1724, n1725, n31357, n134, n135, n136, n137, n138, 
        n139, n140, n141, n142, n143, n144, n145, n146, n147, 
        n148, n149, n150, n151, n152, n153, n154, n155, n156, 
        n157, n158, n159, n160, n161, n162, n163, n164, n165, 
        n44371, n1615, n1616, n1617, n1618, n1619, n1620, n1621, 
        n1622, n1623, n1624, n1625, n31356, n31355, n31354, n1580, 
        n30693, n30692, n30691, n2669, n31353, n2658, n2657, n2656, 
        n2655, n2654, n2653, n2652, n2651, n2650, n2649, n2648, 
        n2647, n2646, n2645, n38287, n2644, n2643_adj_4489, n2642_adj_4490, 
        n2641, n2640, n2639, n2638_adj_4491, n2637_adj_4492, n31352, 
        n1481, n1547, n1516, n1548, n1517, n1549, n1518, n1550, 
        n1519, n1551, n1520, n1552, n1521, n1553_adj_4493, n1522, 
        n1554_adj_4494, n1523, n1555, n1524, n1556, n1525, n1557, 
        n1558, n2636_adj_4495, n1448, n1449, n1450, n1451, n1452, 
        n1453, n1454, n1455, n1456, n1457, n1458, n30554, n30690, 
        n31351, n1417_adj_4496, n1418_adj_4497, n1419_adj_4498, n1420_adj_4499, 
        n1421, n1422, n1423, n1424, n1425, n31350, n30444, n38397, 
        n31349, n30689, n31348, n31347, n31346, n35939, n35941, 
        n18663, n35951, n35953, n35955, n35957, n17255, n30843, 
        n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
        n1357, n1358, n30688, n30687, n2625_adj_4500, n31345, n38371, 
        n31344, n31343, n30842, n30686, n31342, n38313, n31341, 
        n1382, n31340, n1158, n1157, n1318, n1319, n1320, n1321, 
        n1322, n1323, n1324, n1325, n31339, n31338, n2624_adj_4501, 
        n35959, n35961, n35963, n35965, n35967, n35969, n35971, 
        n35973, n2620_adj_4502, n2623_adj_4503, n2621_adj_4504, n2622_adj_4505, 
        n35975, n2619_adj_4506, n2615, n2618_adj_4507, n2616, n2617, 
        n35977, n1156, n2614, n2613, n2612, n2611, n2610, n2609, 
        n2608, n2607, n2606, n2605, n2570, n31337, n30841, n2558_adj_4508, 
        n2557, n2556, n2555, n2554, n2553_adj_4509, n2552_adj_4510, 
        n2551_adj_4511, n2550_adj_4512, n2549_adj_4513, n2548_adj_4514, 
        n2547_adj_4515, n30685, n2546_adj_4516, n2545_adj_4517, n31336, 
        n2544_adj_4518, n2543_adj_4519, n2542_adj_4520, n2_adj_4521, 
        n3_adj_4522, n4_adj_4523, n5_adj_4524, n6_adj_4525, n7_adj_4526, 
        n8_adj_4527, n9_adj_4528, n10_adj_4529, n11_adj_4530, n12_adj_4531, 
        n13_adj_4532, n14_adj_4533, n15_adj_4534, n16_adj_4535, n17_adj_4536, 
        n18_adj_4537, n19_adj_4538, n20_adj_4539, n21_adj_4540, n22_adj_4541, 
        n23_adj_4542, n24_adj_4543, n25_adj_4544, n2_adj_4545, n3_adj_4546, 
        n4_adj_4547, n5_adj_4548, n6_adj_4549, n7_adj_4550, n8_adj_4551, 
        n9_adj_4552, n10_adj_4553, n11_adj_4554, n12_adj_4555, n13_adj_4556, 
        n14_adj_4557, n15_adj_4558, n16_adj_4559, n17_adj_4560, n18_adj_4561, 
        n19_adj_4562, n20_adj_4563, n21_adj_4564, n22_adj_4565, n23_adj_4566, 
        n24_adj_4567, n25_adj_4568, n2541_adj_4569, n2540_adj_4570, 
        n2539_adj_4571, n2538_adj_4572, n2537_adj_4573, n31335, n31334, 
        n2525, n2524, n2523, n2522, n2521, n2520, n2519, n2518, 
        n2517, n2516, n2515, n2514, n2513, n2512, n2511, n2510, 
        n2509, n2508, n2507, n2506, n31333, n31332, n31331, n30443, 
        n2471_adj_4574, n31330, n2458_adj_4575, n2457_adj_4576, n2456_adj_4577, 
        n2455_adj_4578, n2454_adj_4579, n2453_adj_4580, n2452_adj_4581, 
        n2451_adj_4582, n2450_adj_4583, n2449_adj_4584, n2448_adj_4585, 
        n2447_adj_4586, n2446, n2445, n2444, n2443, n2442, n2441, 
        n2440, n2439, n2438, n30684, n31329, n30840, n2425, n2424, 
        n2423, n2422, n2421, n2420, n2419, n2418, n2417, n2416, 
        n2415, n2414, n2413, n2412, n2411, n2410, n2409, n2408, 
        n31328, n2407, n2372_adj_4587, n31327, n31326, n46, n2358_adj_4588, 
        n2357_adj_4589, n2356, n2355, n2354, n2353, n2352, n2351, 
        n2350, n2349, n2348, n2347, n2346, n2345, n2344, n2343, 
        n2342, n2341, n2340, n2339, n44255, n12_adj_4590, n2325, 
        n2324, n2323, n2322, n2321, n2320, n2319, n2318, n2317, 
        n2316, n2315, n2314, n2313, n2312, n2311, n2310, n2309, 
        n2308, n31325, n44, n43291, n2273_adj_4591, n31324, n2258, 
        n2257, n2256, n2255, n2254, n2253, n2252, n2251, n2250, 
        n2249, n2248, n31323, n42_adj_4592, n44969, n2247, n2246, 
        n2245, n2244, n2243, n2242, n2241, n2240, n30683, n31322, 
        n2225, n2224, n2223, n2222, n2221, n2220, n2219, n2218, 
        n2217, n2216, n2215, n2214, n2213, n2212, n2211, n2210, 
        n2209, n31321, n40_adj_4593, n42_adj_4594, n44_adj_4595, n45, 
        n34_adj_4596, n2174_adj_4597, n31320, n2158, n2157, n2156, 
        n2155, n2154, n2153, n2152, n2151, n2150, n2149, n2148, 
        n2147, n2146, n2145, n2144, n2143, n2142, n31319, n38_adj_4598, 
        n40_adj_4599, n42_adj_4600, n43, n44633, n2141, n2_adj_4601, 
        n30839, n30682, n30681, n44383, n2125, n2124, n2123, n2122, 
        n2121, n2120, n2119, n2118, n2117, n2116, n2115, n2114, 
        n2113, n2112, n2111, n2110, n31_adj_4602, n31318, n30_adj_4603, 
        n36_adj_4604, n38_adj_4605, n40_adj_4606, n41_adj_4607, n45035, 
        n44858, n28_adj_4608, n2075_adj_4609, n31317, n44241, n30680, 
        n30553, n31316, n2058, n2057, n2056, n2055, n2054, n2053, 
        n2052, n2051, n2050, n2049, n2048, n31315, n34_adj_4610, 
        n36_adj_4611, n38_adj_4612, n39_adj_4613, n41_adj_4614, n43_adj_4615, 
        n44_adj_4616, n45_adj_4617, n44395, n2047, n2046, n2045, 
        n2044, n2043, n2042, n30442, n43289, n30552, n22_adj_4618, 
        n21_adj_4619, n44393, n2025, n2024, n2023, n2022, n2021, 
        n2020, n2019, n2018, n2017, n2016, n2015, n2014, n2013, 
        n2012, n2011, n31314, n32_adj_4620, n34_adj_4621, n37_adj_4622, 
        n39_adj_4623, n41_adj_4624, n44856, n43_adj_4625, n44397, 
        n44968, n6_adj_4626, n1976_adj_4627, n31313, n31312, n30_adj_4628, 
        n31_adj_4629, n32_adj_4630, n33_adj_4631, n34_adj_4632, n35_adj_4633, 
        n37_adj_4634, n39_adj_4635, n44649, n41_adj_4636, n42_adj_4637, 
        n43_adj_4638, n45_adj_4639, n43277, n1958, n1957, n1956, 
        n1955, n1954, n1953, n3362, n1952, n1951, n1950, n1949, 
        n1948, n1947, n1946, n1945, n1944, n1943, n30551, n30550, 
        n31311, n28_adj_4640, n29_adj_4641, n30_adj_4642, n31_adj_4643, 
        n32_adj_4644, n33_adj_4645, n35_adj_4646, n37_adj_4647, n44846, 
        n39_adj_4648, n40_adj_4649, n41_adj_4650, n43_adj_4651, n44972, 
        n45002, n31310, n1925, n1924, n1923, n1922, n1921, n1920, 
        n1919, n1918, n3323, n1917, n1916, n1915, n1914, n1913, 
        n1912, n31309, n26_adj_4652, n27_adj_4653, n28_adj_4654, n29_adj_4655, 
        n30_adj_4656, n31_adj_4657, n33_adj_4658, n35_adj_4659, n44974, 
        n37_adj_4660, n38_adj_4661, n39_adj_4662, n41_adj_4663, n45037, 
        n30441, n7040, n1877, n31308, n31307, n24_adj_4664, n25_adj_4665, 
        n26_adj_4666, n27_adj_4667, n28_adj_4668, n29_adj_4669, n30_adj_4670, 
        n31_adj_4671, n32_adj_4672, n33_adj_4673, n35_adj_4674, n36_adj_4675, 
        n37_adj_4676, n39_adj_4677, n41_adj_4678, n44854, n43_adj_4679, 
        n45_adj_4680, n44663, n1858, n1857, n1856, n3253, n1855, 
        n1854, n1853, n1852, n1851, n1850, n1849, n1848, n1847, 
        n1846, n1845, n1844, n30838, n31306, n22_adj_4681, n22_adj_4682, 
        n23_adj_4683, n24_adj_4684, n25_adj_4685, n26_adj_4686, n27_adj_4687, 
        n28_adj_4688, n29_adj_4689, n30_adj_4690, n31_adj_4691, n33_adj_4692, 
        n34_adj_4693, n35_adj_4694, n37_adj_4695, n39_adj_4696, n44850, 
        n41_adj_4697, n43_adj_4698, n43260, n3223, n1825, n1824, 
        n1823, n1822, n1821, n1820, n1819, n1818, n1817, n1816, 
        n1815, n19_adj_4699, n20_adj_4700, n21_adj_4701, n22_adj_4702, 
        n23_adj_4703, n24_adj_4704, n25_adj_4705, n26_adj_4706, n27_adj_4707, 
        n28_adj_4708, n29_adj_4709, n31_adj_4710, n32_adj_4711, n33_adj_4712, 
        n35_adj_4713, n37_adj_4714, n44844, n39_adj_4715, n41_adj_4716, 
        n1814, n1813, n7136, n18_adj_4717, n31305, n18_adj_4718, 
        n19_adj_4719, n20_adj_4720, n21_adj_4721, n22_adj_4722, n23_adj_4723, 
        n24_adj_4724, n25_adj_4725, n26_adj_4726, n27_adj_4727, n29_adj_4728, 
        n30_adj_4729, n31_adj_4730, n33_adj_4731, n35_adj_4732, n44824, 
        n37_adj_4733, n39_adj_4734, n41_adj_4735, n43_adj_4736, n45_adj_4737, 
        n44673, n1778_adj_4738, n31304, n31303, n16_adj_4739, n16_adj_4740, 
        n17_adj_4741, n18_adj_4742, n19_adj_4743, n20_adj_4744, n21_adj_4745, 
        n22_adj_4746, n23_adj_4747, n25_adj_4748, n27_adj_4749, n28_adj_4750, 
        n29_adj_4751, n31_adj_4752, n33_adj_4753, n35_adj_4754, n44597, 
        n37_adj_4755, n39_adj_4756, n41_adj_4757, n43_adj_4758, n45053, 
        n30549, n31302, n3150, n31301, n31300, n14_adj_4759, n16_adj_4760, 
        n17_adj_4761, n18_adj_4762, n19_adj_4763, n20_adj_4764, n21_adj_4765, 
        n22_adj_4766, n23_adj_4767, n25_adj_4768, n26_adj_4769, n27_adj_4770, 
        n29_adj_4771, n31_adj_4772, n44806, n33_adj_4773, n35_adj_4774, 
        n37_adj_4775, n39_adj_4776, n40_adj_4777, n41_adj_4778, n43_adj_4779, 
        n45_adj_4780, n45004, n1758_adj_4781, n1757_adj_4782, n1756_adj_4783, 
        n1755_adj_4784, n3132, n1754_adj_4785, n1753, n1752, n1751, 
        n1750, n1749, n1748, n12_adj_4786, n14_adj_4787, n15_adj_4788, 
        n16_adj_4789, n17_adj_4790, n18_adj_4791, n19_adj_4792, n20_adj_4793, 
        n21_adj_4794, n23_adj_4795, n24_adj_4796, n25_adj_4797, n27_adj_4798, 
        n29_adj_4799, n31_adj_4800, n44588, n33_adj_4801, n35_adj_4802, 
        n37_adj_4803, n38_adj_4804, n39_adj_4805, n41_adj_4806, n43_adj_4807, 
        n44828, n1747, n1746, n1745, n3117, n30679, n31299, n10_adj_4808, 
        n12_adj_4809, n13_adj_4810, n14_adj_4811, n15_adj_4812, n16_adj_4813, 
        n17_adj_4814, n18_adj_4815, n19_adj_4816, n21_adj_4817, n22_adj_4818, 
        n23_adj_4819, n25_adj_4820, n27_adj_4821, n29_adj_4822, n45039, 
        n31_adj_4823, n33_adj_4824, n44980, n35_adj_4825, n36_adj_4826, 
        n37_adj_4827, n39_adj_4828, n41_adj_4829, n44691, n44882, 
        n45124, n3105, n31298, n8_adj_4830, n10_adj_4831, n11_adj_4832, 
        n12_adj_4833, n13_adj_4834, n14_adj_4835, n15_adj_4836, n16_adj_4837, 
        n17_adj_4838, n19_adj_4839, n20_adj_4840, n21_adj_4841, n23_adj_4842, 
        n25_adj_4843, n27_adj_4844, n29_adj_4845, n31_adj_4846, n44818, 
        n33_adj_4847, n34_adj_4848, n35_adj_4849, n37_adj_4850, n39_adj_4851, 
        n44694, n41_adj_4852, n43_adj_4853, n44_adj_4854, n45_adj_4855, 
        n44696, n31297, n6_adj_4856, n8_adj_4857, n9_adj_4858, n10_adj_4859, 
        n11_adj_4860, n12_adj_4861, n13_adj_4862, n14_adj_4863, n15_adj_4864, 
        n17_adj_4865, n19_adj_4866, n21_adj_4867, n23_adj_4868, n24_adj_4869, 
        n25_adj_4870, n27_adj_4871, n29_adj_4872, n30_adj_4873, n31_adj_4874, 
        n32_adj_4875, n33_adj_4876, n35_adj_4877, n37_adj_4878, n44978, 
        n45125, n44584, n31296, n4_adj_4879, n6_adj_4880, n7_adj_4881, 
        n8_adj_4882, n9_adj_4883, n10_adj_4884, n11_adj_4885, n12_adj_4886, 
        n13_adj_4887, n15_adj_4888, n16_adj_4889, n17_adj_4890, n19_adj_4891, 
        n21_adj_4892, n23_adj_4893, n24_adj_4894, n25_adj_4895, n27_adj_4896, 
        n29_adj_4897, n30_adj_4898, n31_adj_4899, n33_adj_4900, n35_adj_4901, 
        n37_adj_4902, n39_adj_4903, n41_adj_4904, n43_adj_4905, n44706, 
        n45_adj_4906, n45010, n31295, n30678, n30548, n30837, n2_adj_4907, 
        n30836, n31294, n30835, n30834, n45041, n31293, n31292, 
        n31291, n43224, n35947, n31290, n30_adj_4908, n29_adj_4909, 
        n35923, n19_adj_4910, n31289, n11_adj_4911, n38070, n35907, 
        n44661, n28_adj_4912, n27_adj_4913, n18_adj_4914, n31288, 
        n43205, n31287, n43203, n31286, n38299, n44151, n5_adj_4915, 
        n44149, n31285, n8_adj_4916, n46050, n44689, n45008, n31284, 
        n31283, n8_adj_4917, n7_adj_4918, n31282, n45121, n31281, 
        n31280, n43186, n43184, n43178, n16_adj_4919, n11_adj_4920, 
        n10_adj_4921, n44417, n31279, n43176, n31278, n31277, n31276, 
        n31275, n44107, n43172, n43164, n31274, n31273, n45935, 
        n31272, n31271, n6_adj_4922, n44091, n31270, n38358, n30833, 
        n30440, n31269, n30832, n30677, n44421, n30676, n43128, 
        n30831, n30830, n30439, n30829, n30828, n31268, n31267, 
        n30827, n30675, n27445, n31266, n30674, n38343, n31265, 
        n31264, n31263, n31262, n30438, n31261, n31260, n31259, 
        n31258, n30826, n38405, n30673, n31257, n31256, n30672, 
        n31255, n30671, n31254, n31253, n30437, n44039, n31252, 
        n43101, n31251, n28_adj_4923, n40693, n26_adj_4924, n40689, 
        n24_adj_4925, n31250, n31249, n19_adj_4926, n43092, n44010, 
        n16_adj_4927, n44004, n40673, n44002, n31248, n30670, n31247, 
        n30436, n31246, n30825, n31245, n43079, n31244, n30669, 
        n44813, n30668, n43986, n43984, n43980, n43074, n43978, 
        n43070, n43970, n43068, n43968, n43964, n43962, n45038, 
        n43066, n43056, n44445, n43948, n31243, n31242, n43944, 
        n31241, n31240, n38353, n31239, n31238, n43940, n31237, 
        n31236, n39_adj_4928, n31235, n43048, n30824, n31234, n37_adj_4929, 
        n44811, n36_adj_4930, n43044, n34_adj_4931, n33_adj_4932, 
        n43925, n44447, n44809, n24672, n45126, n27_adj_4933, n43034, 
        n31233, n43028, n22_adj_4934, n43024, n43022, n31232, n44808, 
        n30667, n31231, n37348, n31230, n19208, n19207, n31229, 
        n31228, n30823, n30822, n43012, n31227, n43010, n31226, 
        n31225, n31224, n19206, n19203, n31223, n31222, n31221, 
        n43004, n43002, n44805, n43000, n42993, n44803, n45034, 
        n44113, n20_adj_4935, n18_adj_4936, n16_adj_4937, n31220, 
        n31219, n31218, n31217, n30435, n31216, n31215, n45033, 
        n31214, n6996, n31213, n31212, n31211, n31210, n30666, 
        n31209, n31208, n44748, n39307, n43684, n43678, n42970, 
        n44918, n43727, n42968, n43664, n42966, n43680, n43676, 
        n42965, n19205, n42964, n42963, n42962, n42961, n42960, 
        n42959, n43718, n42958, n42957, n42956, n42955, n42954, 
        n42953, n2_adj_4938, n3_adj_4939, n4_adj_4940, n5_adj_4941, 
        n6_adj_4942, n7_adj_4943, n8_adj_4944, n9_adj_4945, n10_adj_4946, 
        n11_adj_4947, n12_adj_4948, n13_adj_4949, n14_adj_4950, n15_adj_4951, 
        n16_adj_4952, n17_adj_4953, n18_adj_4954, n19_adj_4955, n20_adj_4956, 
        n21_adj_4957, n22_adj_4958, n23_adj_4959, n24_adj_4960, n25_adj_4961, 
        n26_adj_4962, n27_adj_4963, n28_adj_4964, n29_adj_4965, n30_adj_4966, 
        n31_adj_4967, n32_adj_4968, n33_adj_4969, n42952, n44796, 
        n42951, n19204, n19202, n42950, n42949, n30821, n30665, 
        n30664, n42948, n38389, n42947, n30820, n30434, n42946, 
        n44754, n42945, n30663, n40501, n42944, n42943, n42942, 
        n42941, n42940, n30662, n42939, n30819, n30661, n45020, 
        n45123, n30818, n42936, n31143, n31142, n31141, n30817, 
        n42935, n42934, n42933, n31140, n31139, n30660, n31138, 
        n30433, n30816, n31137, n31136, n31135, n30815, n31134, 
        n31133, n30659, n31132, n31131, n30658, n31130, n31129, 
        n31128, n30657, n31127, n31126, n31125, n31124, n31123, 
        n31122, n31121, n31120, n31119, n31118, n31117, n31116, 
        n31115, n42920, n42919, n31114, n36695, n31113, n31112, 
        n31111, n31110, n30656, n30655, n30654, n30814, n30813, 
        n31109, n31108, n30812, n30811, n30653, n30652, n30651, 
        n30810, n31107, n30650, n30809, n31106, n30808, n31105, 
        n31104, n31103, n31102, n31101, n30649, n30807, n30806, 
        n30648, n31100, n31099, n30647, n30646, n31098, n31097, 
        n30645, n17281, n31096, n31095, n30805, n30804, n17278, 
        n31094, n30644, n31093, n30803, n31092, n31091, n30802, 
        n31090, n30801, n30800, n31089, n31088, n31087, n31086, 
        n17275, n30799, n30643, n30642, n30798, n31085, n43815, 
        n31084, n31083, n31082, n31081, n31080, n30797, n30641, 
        n30796, n40433, n31079, n31078, n31077, n38251, n44515, 
        n31076, n31075, n31074, n31073, n30640, n31072, n30795, 
        n31071, n31070, n30639, n31069, n31068, n30794, n30638, 
        n31067, n30793, n30637, n30792, n31066, n31065, n31064, 
        n31063, n31062, n31061, n31060, n31059, n31058, n30791, 
        n36_adj_4970, n31057, n31056, n31055, n31054, n31053, n35_adj_4971, 
        n45029, n31052, n31051, n31050, n31049, n31048, n31047, 
        n31046, n34_adj_4972, n30790, n33_adj_4973, n30636, n31045, 
        n30635, n31044, n31043, n31042, n31041, n31040, n31039, 
        n31038, n31037, n31036, n31035, n31034, n31033, n31032, 
        n31031, n31030, n30634, n31029, n31028, n31027, n31026, 
        n31025, n31024, n31023, n31022, n31021, n31020, n31019, 
        n31018, n30633, n31017, n31016, n31015, n31014, n31013, 
        n31012, n31011, n31010, n31009, n31008, n31007, n31_adj_4974, 
        n30789, n31006, n31005, n31004, n31003, n31002, n31001, 
        n31000, n30999, n30998, n30632, n30997, n30996, n30995, 
        n40407, n30994, n30631, n30993, n30992, n30991, n30630, 
        n17296, n40403, n24_adj_4975, n40397, n30990, n30989, n30988, 
        n30987, n30986, n30985, n30984, n30983, n30982, n30788, 
        n30981, n30980, n30629, n30979, n30978, n40389, n38410, 
        n38239, n40387, n30977, n30976, n47, n40385, n30975, n30628, 
        n30974, n30627, n40383, n46_adj_4976, n30973, n30626, n30972, 
        n43_adj_4977, n30625, n42_adj_4978, n30971, n30970, n30969, 
        n40381, n40_adj_4979, n30968, n30967, n30966, n30624, n30965, 
        n30964, n30623, n30622, n30963, n30962, n39036, n40379, 
        n30961, n30960, n30959, n30787, n39_adj_4980, n30958, n38_adj_4981, 
        n30957, n30956, n30955, n30954, n30953, n30621, n30952, 
        n40377, n30951, n30950, n30949, n30620, n30948, n30947, 
        n30946, n30945, n45142, n32_adj_4982, n45028, n26_adj_4983, 
        n24_adj_4984, n22_adj_4985, n18_adj_4986, n44764, n38306, 
        n43835, n45026, n36597, n43753, n37214, n41_adj_4987, n40_adj_4988, 
        n42871, n45865, n40311, n44600, n40309, n40303, n40301, 
        n40299, n43839, n40287, n40281, n40253, n40249, n38192, 
        n40805, n44599, n5_adj_4989, n37216, n16_adj_4990, n40223, 
        n44770, n36743, n43847, n38098, n38094, n44594, n45118, 
        n45862, n44_adj_4991, n43_adj_4992, n42_adj_4993, n41_adj_4994, 
        n40_adj_4995, n38_adj_4996, n30_adj_4997, n38026, n26_adj_4998, 
        n38024, n36919, n37218, n44553, n38022, n39906, n36983, 
        n37215, n37220, n37219, n37217, n28_adj_4999, n27_adj_5000, 
        n26_adj_5001, n25_adj_5002, n47_adj_5003, n46_adj_5004, n39886, 
        n28_adj_5005, n40021, n40019, n45119, n38376, n39863, n40712;
    
    VCC i2 (.Y(VCC_net));
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[0]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF h2_46 (.Q(PIN_21_c), .C(clk32MHz), .D(hall2));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_80[0]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_IO hall2_input (.PACKAGE_PIN(PIN_4), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(PIN_5), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(PIN_12), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), 
          .D_OUT_1(GND_net), .D_OUT_0(tx_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_6_pad (.PACKAGE_PIN(PIN_6), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_6_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_6_pad.PIN_TYPE = 6'b000001;
    defparam PIN_6_pad.PULLUP = 1'b0;
    defparam PIN_6_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_DFF h3_47 (.Q(PIN_22_c), .C(clk32MHz), .D(hall3));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF dir_51 (.Q(PIN_23_c), .C(clk32MHz), .D(duty[23]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_LUT4 rem_4_i1668_3_lut (.I0(n2451_adj_4582), .I1(n2518), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2550_adj_4512));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_IO ID0_input (.PACKAGE_PIN(PIN_9), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), .D_OUT_1(GND_net), 
          .D_OUT_0(GND_net), .D_IN_0(ID0)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ID0_input.PIN_TYPE = 6'b000001;
    defparam ID0_input.PULLUP = 1'b1;
    defparam ID0_input.NEG_TRIGGER = 1'b0;
    defparam ID0_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO ID1_input (.PACKAGE_PIN(PIN_10), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(ID1)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ID1_input.PIN_TYPE = 6'b000001;
    defparam ID1_input.PULLUP = 1'b1;
    defparam ID1_input.NEG_TRIGGER = 1'b0;
    defparam ID1_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO ID2_input (.PACKAGE_PIN(PIN_11), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(ID2)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ID2_input.PIN_TYPE = 6'b000001;
    defparam ID2_input.PULLUP = 1'b1;
    defparam ID2_input.NEG_TRIGGER = 1'b0;
    defparam ID2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall1_input (.PACKAGE_PIN(PIN_3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 rem_4_i1666_3_lut (.I0(n2449_adj_4584), .I1(n2516), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2548_adj_4514));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(n37220), .I1(r_Clock_Count[6]), .I2(n16_adj_4990), 
            .I3(GND_net), .O(n36743));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut.LUT_INIT = 16'heaea;
    neopixel nx (.timer({timer}), .GND_net(GND_net), .\neo_pixel_transmitter.done (\neo_pixel_transmitter.done ), 
            .clk32MHz(clk32MHz), .n42947(n42947), .bit_ctr({bit_ctr}), 
            .n19(n19_adj_4910), .n42956(n42956), .n35971(n35971), .n35973(n35973), 
            .n35975(n35975), .n35967(n35967), .n35969(n35969), .n35963(n35963), 
            .n35965(n35965), .n35959(n35959), .n35961(n35961), .n35955(n35955), 
            .n35957(n35957), .n35951(n35951), .n35953(n35953), .n35947(n35947), 
            .n35949(n35949), .n35933(n35933), .n35935(n35935), .n35937(n35937), 
            .n35939(n35939), .n35941(n35941), .n35943(n35943), .n35931(n35931), 
            .n35925(n35925), .n35907(n35907), .VCC_net(VCC_net), .n35927(n35927), 
            .n35909(n35909), .n35911(n35911), .n35929(n35929), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .\one_wire_N_513[11] (one_wire_N_513[11]), .n42943(n42943), 
            .n10(n10_adj_4350), .n42966(n42966), .\one_wire_N_513[7] (one_wire_N_513[7]), 
            .n8(n8_adj_4437), .n42955(n42955), .\one_wire_N_513[5] (one_wire_N_513[5]), 
            .n42965(n42965), .n42964(n42964), .n42954(n42954), .n38094(n38094), 
            .\state[1] (state[1]), .n42963(n42963), .start(start), .n42968(n42968), 
            .n42962(n42962), .n35923(n35923), .n42953(n42953), .n42961(n42961), 
            .\state_3__N_362[1] (state_3__N_362[1]), .n27365(n27365), .n17195(n17195), 
            .n38070(n38070), .n35913(n35913), .n35917(n35917), .n35915(n35915), 
            .n18886(n18886), .n18885(n18885), .n18884(n18884), .n18883(n18883), 
            .n18882(n18882), .n18881(n18881), .n18880(n18880), .n18879(n18879), 
            .n18878(n18878), .n18877(n18877), .n18876(n18876), .n18875(n18875), 
            .n18874(n18874), .n18873(n18873), .n18872(n18872), .n18871(n18871), 
            .n18870(n18870), .n18869(n18869), .n18868(n18868), .n18867(n18867), 
            .n18866(n18866), .n18865(n18865), .n18864(n18864), .n18863(n18863), 
            .n18862(n18862), .n18861(n18861), .n18860(n18860), .n18859(n18859), 
            .n18858(n18858), .n18857(n18857), .n18856(n18856), .n18855(n18855), 
            .\state[0] (state[0]), .n38192(n38192), .n42960(n42960), .n42952(n42952), 
            .n18416(n18416), .n18584(n18584), .n42959(n42959), .n42951(n42951), 
            .n42950(n42950), .n35977(n35977), .n42946(n42946), .n42945(n42945), 
            .PIN_8_c(PIN_8_c), .n42939(n42939), .n11(n11_adj_4911), .n42940(n42940), 
            .n42958(n42958), .n42936(n42936), .n42935(n42935), .n18663(n18663), 
            .n42934(n42934), .n42957(n42957), .n42933(n42933), .n42944(n42944), 
            .n42942(n42942), .n42941(n42941), .n42949(n42949), .n42948(n42948), 
            .n1105(n1105), .n4754(n4754), .n27453(n27453), .n39307(n39307), 
            .\color[20] (color[20]), .\color[21] (color[21]), .\color[17] (color[17])) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(64[10] 70[2])
    SB_LUT4 rem_4_i1662_3_lut (.I0(n2445), .I1(n2512), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2544_adj_4518));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1050_10_lut (.I0(GND_net), .I1(n1551), .I2(VCC_net), 
            .I3(n31393), .O(n1618)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1671_3_lut (.I0(n2454_adj_4579), .I1(n2521), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2553_adj_4509));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1050_10 (.CI(n31393), .I0(n1551), .I1(VCC_net), 
            .CO(n31394));
    SB_LUT4 rem_4_i1663_3_lut (.I0(n2446), .I1(n2513), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2545_adj_4517));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1772_3_lut_3_lut (.I0(n2642), .I1(n7154), .I2(n2636), 
            .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1772_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1659_3_lut (.I0(n2442), .I1(n2509), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2541_adj_4569));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1754_3_lut_3_lut (.I0(n2642), .I1(n7136), .I2(n2618), 
            .I3(GND_net), .O(n2699));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1754_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1657_3_lut (.I0(n2440), .I1(n2507), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2539_adj_4571));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14397_3_lut (.I0(setpoint[3]), .I1(n4662), .I2(n39863), .I3(GND_net), 
            .O(n19429));   // verilog/coms.v(126[12] 289[6])
    defparam i14397_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1673_3_lut (.I0(n2456_adj_4577), .I1(n2523), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2555));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1661_3_lut (.I0(n2444), .I1(n2511), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2543_adj_4519));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1050_9_lut (.I0(GND_net), .I1(n1552), .I2(VCC_net), 
            .I3(n31392), .O(n1619)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_9 (.CI(n31392), .I0(n1552), .I1(VCC_net), 
            .CO(n31393));
    SB_LUT4 rem_4_add_1050_8_lut (.I0(GND_net), .I1(n1553_adj_4493), .I2(VCC_net), 
            .I3(n31391), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_8 (.CI(n31391), .I0(n1553_adj_4493), .I1(VCC_net), 
            .CO(n31392));
    SB_LUT4 rem_4_add_1050_7_lut (.I0(GND_net), .I1(n1554_adj_4494), .I2(GND_net), 
            .I3(n31390), .O(n1621)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_7 (.CI(n31390), .I0(n1554_adj_4494), .I1(GND_net), 
            .CO(n31391));
    SB_LUT4 rem_4_add_1050_6_lut (.I0(GND_net), .I1(n1555), .I2(GND_net), 
            .I3(n31389), .O(n1622)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_6 (.CI(n31389), .I0(n1555), .I1(GND_net), 
            .CO(n31390));
    SB_LUT4 rem_4_add_1050_5_lut (.I0(GND_net), .I1(n1556), .I2(VCC_net), 
            .I3(n31388), .O(n1623)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i1755_3_lut_3_lut (.I0(n2642), .I1(n7137), .I2(n2619), 
            .I3(GND_net), .O(n2700));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1755_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1672_3_lut (.I0(n2455_adj_4578), .I1(n2522), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2554));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1050_5 (.CI(n31388), .I0(n1556), .I1(VCC_net), 
            .CO(n31389));
    SB_LUT4 rem_4_add_1050_4_lut (.I0(GND_net), .I1(n1557), .I2(VCC_net), 
            .I3(n31387), .O(n1624)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_4 (.CI(n31387), .I0(n1557), .I1(VCC_net), 
            .CO(n31388));
    SB_LUT4 rem_4_add_1050_3_lut (.I0(GND_net), .I1(n1558), .I2(GND_net), 
            .I3(n31386), .O(n1625)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_3 (.CI(n31386), .I0(n1558), .I1(GND_net), 
            .CO(n31387));
    SB_CARRY rem_4_add_1050_2 (.CI(VCC_net), .I0(n1658), .I1(VCC_net), 
            .CO(n31386));
    SB_LUT4 rem_4_add_1117_15_lut (.I0(n1679), .I1(n1646_adj_4481), .I2(VCC_net), 
            .I3(n31385), .O(n1745)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1117_14_lut (.I0(GND_net), .I1(n1647_adj_4482), .I2(VCC_net), 
            .I3(n31384), .O(n1714)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_14 (.CI(n31384), .I0(n1647_adj_4482), .I1(VCC_net), 
            .CO(n31385));
    SB_LUT4 rem_4_i1665_3_lut (.I0(n2448_adj_4585), .I1(n2515), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2547_adj_4515));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1117_13_lut (.I0(GND_net), .I1(n1648_adj_4483), .I2(VCC_net), 
            .I3(n31383), .O(n1715)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_13 (.CI(n31383), .I0(n1648_adj_4483), .I1(VCC_net), 
            .CO(n31384));
    SB_LUT4 rem_4_add_1117_12_lut (.I0(GND_net), .I1(n1649_adj_4484), .I2(VCC_net), 
            .I3(n31382), .O(n1716)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1664_3_lut (.I0(n2447_adj_4586), .I1(n2514), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2546_adj_4516));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1117_12 (.CI(n31382), .I0(n1649_adj_4484), .I1(VCC_net), 
            .CO(n31383));
    SB_LUT4 div_36_i1758_3_lut_3_lut (.I0(n2642), .I1(n7140), .I2(n2622), 
            .I3(GND_net), .O(n2703));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1758_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1670_3_lut (.I0(n2453_adj_4580), .I1(n2520), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2552_adj_4510));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1667_3_lut (.I0(n2450_adj_4583), .I1(n2517), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2549_adj_4513));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1756_3_lut_3_lut (.I0(n2642), .I1(n7138), .I2(n2620), 
            .I3(GND_net), .O(n2701));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1756_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1660_3_lut (.I0(n2443), .I1(n2510), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2542_adj_4520));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1658_3_lut (.I0(n2441), .I1(n2508), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2540_adj_4570));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1117_11_lut (.I0(GND_net), .I1(n1650_adj_4485), .I2(VCC_net), 
            .I3(n31381), .O(n1717)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1656_3_lut (.I0(n2439), .I1(n2506), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2538_adj_4572));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1675_3_lut (.I0(n2458_adj_4575), .I1(n2525), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2557));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1757_3_lut_3_lut (.I0(n2642), .I1(n7139), .I2(n2621), 
            .I3(GND_net), .O(n2702));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1757_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1674_3_lut (.I0(n2457_adj_4576), .I1(n2524), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2556));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1610 (.I0(n2556), .I1(n2557), .I2(n2558_adj_4508), 
            .I3(GND_net), .O(n38313));
    defparam i1_3_lut_adj_1610.LUT_INIT = 16'hfefe;
    SB_LUT4 div_36_i1761_3_lut_3_lut (.I0(n2642), .I1(n7143), .I2(n2625), 
            .I3(GND_net), .O(n2706));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1761_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10_4_lut (.I0(n2538_adj_4572), .I1(n2540_adj_4570), .I2(n2537_adj_4573), 
            .I3(n2542_adj_4520), .O(n28_adj_4608));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(n2549_adj_4513), .I1(n2552_adj_4510), .I2(n2546_adj_4516), 
            .I3(n2547_adj_4515), .O(n31_adj_4602));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1611 (.I0(n37217), .I1(r_Clock_Count[5]), .I2(n16_adj_4990), 
            .I3(GND_net), .O(n36919));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_1611.LUT_INIT = 16'heaea;
    SB_LUT4 i1_3_lut_adj_1612 (.I0(n37216), .I1(r_Clock_Count[4]), .I2(n16_adj_4990), 
            .I3(GND_net), .O(n36989));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_1612.LUT_INIT = 16'heaea;
    SB_LUT4 i1_3_lut_adj_1613 (.I0(n37218), .I1(r_Clock_Count[3]), .I2(n16_adj_4990), 
            .I3(GND_net), .O(n36987));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_1613.LUT_INIT = 16'heaea;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n95), 
            .I3(r_Rx_Data), .O(n16_adj_4990));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_4_lut.LUT_INIT = 16'hbaaa;
    SB_LUT4 i4_4_lut (.I0(n2554), .I1(n2543_adj_4519), .I2(n38313), .I3(n2555), 
            .O(n22_adj_4618));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i4_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i12_4_lut (.I0(n2545_adj_4517), .I1(n2553_adj_4509), .I2(n2544_adj_4518), 
            .I3(n2548_adj_4514), .O(n30_adj_4603));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_36_i1762_3_lut_3_lut (.I0(n2642), .I1(n7144), .I2(n2626), 
            .I3(GND_net), .O(n2707));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1762_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i16_4_lut (.I0(n31_adj_4602), .I1(n2550_adj_4512), .I2(n28_adj_4608), 
            .I3(n2551_adj_4511), .O(n34_adj_4596));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_36_i1759_3_lut_3_lut (.I0(n2642), .I1(n7141), .I2(n2623), 
            .I3(GND_net), .O(n2704));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1759_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1760_3_lut_3_lut (.I0(n2642), .I1(n7142), .I2(n2624), 
            .I3(GND_net), .O(n2705));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1760_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i3_2_lut (.I0(n2539_adj_4571), .I1(n2541_adj_4569), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4619));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i17_4_lut (.I0(n21_adj_4619), .I1(n34_adj_4596), .I2(n30_adj_4603), 
            .I3(n22_adj_4618), .O(n2570));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_36_i1775_3_lut_3_lut (.I0(n2642), .I1(n7157), .I2(n389), 
            .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1775_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1764_3_lut_3_lut (.I0(n2642), .I1(n7146), .I2(n2628), 
            .I3(GND_net), .O(n2709));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1764_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1765_3_lut_3_lut (.I0(n2642), .I1(n7147), .I2(n2629), 
            .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1765_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4418));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_i1766_3_lut_3_lut (.I0(n2642), .I1(n7148), .I2(n2630), 
            .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1766_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1767_3_lut_3_lut (.I0(n2642), .I1(n7149), .I2(n2631), 
            .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1767_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13949_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18981));   // verilog/coms.v(126[12] 289[6])
    defparam i13949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13950_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18982));   // verilog/coms.v(126[12] 289[6])
    defparam i13950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14011_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position[1]), 
            .I2(n14536), .I3(GND_net), .O(n19043));   // verilog/coms.v(126[12] 289[6])
    defparam i14011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13951_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18983));   // verilog/coms.v(126[12] 289[6])
    defparam i13951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13952_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18984));   // verilog/coms.v(126[12] 289[6])
    defparam i13952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13953_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18985));   // verilog/coms.v(126[12] 289[6])
    defparam i13953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14012_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position[2]), 
            .I2(n14536), .I3(GND_net), .O(n19044));   // verilog/coms.v(126[12] 289[6])
    defparam i14012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14013_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position[3]), 
            .I2(n14536), .I3(GND_net), .O(n19045));   // verilog/coms.v(126[12] 289[6])
    defparam i14013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14014_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position[4]), 
            .I2(n14536), .I3(GND_net), .O(n19046));   // verilog/coms.v(126[12] 289[6])
    defparam i14014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14015_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position[5]), 
            .I2(n14536), .I3(GND_net), .O(n19047));   // verilog/coms.v(126[12] 289[6])
    defparam i14015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13954_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18986));   // verilog/coms.v(126[12] 289[6])
    defparam i13954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14016_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position[6]), 
            .I2(n14536), .I3(GND_net), .O(n19048));   // verilog/coms.v(126[12] 289[6])
    defparam i14016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1773_3_lut_3_lut (.I0(n2642), .I1(n7155), .I2(n2637), 
            .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1773_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14017_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position[7]), 
            .I2(n14536), .I3(GND_net), .O(n19049));   // verilog/coms.v(126[12] 289[6])
    defparam i14017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14018_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n14536), .I3(GND_net), .O(n19050));   // verilog/coms.v(126[12] 289[6])
    defparam i14018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14019_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n14536), .I3(GND_net), .O(n19051));   // verilog/coms.v(126[12] 289[6])
    defparam i14019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1774_3_lut_3_lut (.I0(n2642), .I1(n7156), .I2(n2638), 
            .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1774_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14020_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n14536), .I3(GND_net), .O(n19052));   // verilog/coms.v(126[12] 289[6])
    defparam i14020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14021_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n14536), .I3(GND_net), .O(n19053));   // verilog/coms.v(126[12] 289[6])
    defparam i14021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14022_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n14536), .I3(GND_net), .O(n19054));   // verilog/coms.v(126[12] 289[6])
    defparam i14022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1768_3_lut_3_lut (.I0(n2642), .I1(n7150), .I2(n2632), 
            .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1768_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14023_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n14536), .I3(GND_net), .O(n19055));   // verilog/coms.v(126[12] 289[6])
    defparam i14023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14024_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n14536), .I3(GND_net), .O(n19056));   // verilog/coms.v(126[12] 289[6])
    defparam i14024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14025_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n14536), .I3(GND_net), .O(n19057));   // verilog/coms.v(126[12] 289[6])
    defparam i14025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13955_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18987));   // verilog/coms.v(126[12] 289[6])
    defparam i13955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1770_3_lut_3_lut (.I0(n2642), .I1(n7152), .I2(n2634), 
            .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1770_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14026_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n14536), .I3(GND_net), .O(n19058));   // verilog/coms.v(126[12] 289[6])
    defparam i14026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14027_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n14536), .I3(GND_net), .O(n19059));   // verilog/coms.v(126[12] 289[6])
    defparam i14027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13956_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18988));   // verilog/coms.v(126[12] 289[6])
    defparam i13956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1769_3_lut_3_lut (.I0(n2642), .I1(n7151), .I2(n2633), 
            .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1769_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1763_3_lut_3_lut (.I0(n2642), .I1(n7145), .I2(n2627), 
            .I3(GND_net), .O(n2708));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1763_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4417));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_i1771_3_lut_3_lut (.I0(n2642), .I1(n7153), .I2(n2635), 
            .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1771_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13957_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18989));   // verilog/coms.v(126[12] 289[6])
    defparam i13957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i28_1_lut (.I0(communication_counter[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4942));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14028_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n14536), .I3(GND_net), .O(n19060));   // verilog/coms.v(126[12] 289[6])
    defparam i14028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13958_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18990));   // verilog/coms.v(126[12] 289[6])
    defparam i13958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14029_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n14536), .I3(GND_net), .O(n19061));   // verilog/coms.v(126[12] 289[6])
    defparam i14029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14030_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n14536), .I3(GND_net), .O(n19062));   // verilog/coms.v(126[12] 289[6])
    defparam i14030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14031_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n14536), .I3(GND_net), .O(n19063));   // verilog/coms.v(126[12] 289[6])
    defparam i14031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14236_3_lut (.I0(\data_in_frame[15] [3]), .I1(rx_data[3]), 
            .I2(n37348), .I3(GND_net), .O(n19268));   // verilog/coms.v(126[12] 289[6])
    defparam i14236_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14032_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n14536), .I3(GND_net), .O(n19064));   // verilog/coms.v(126[12] 289[6])
    defparam i14032_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1117_11 (.CI(n31381), .I0(n1650_adj_4485), .I1(VCC_net), 
            .CO(n31382));
    SB_LUT4 i14237_3_lut (.I0(\data_in_frame[15] [4]), .I1(rx_data[4]), 
            .I2(n37348), .I3(GND_net), .O(n19269));   // verilog/coms.v(126[12] 289[6])
    defparam i14237_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14033_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n14536), .I3(GND_net), .O(n19065));   // verilog/coms.v(126[12] 289[6])
    defparam i14033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14034_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n14536), .I3(GND_net), .O(n19066));   // verilog/coms.v(126[12] 289[6])
    defparam i14034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14035_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n14536), .I3(GND_net), .O(n19067));   // verilog/coms.v(126[12] 289[6])
    defparam i14035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14036_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n14536), .I3(GND_net), .O(n19068));   // verilog/coms.v(126[12] 289[6])
    defparam i14036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13959_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18991));   // verilog/coms.v(126[12] 289[6])
    defparam i13959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i29_1_lut (.I0(communication_counter[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4941));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14037_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n14536), .I3(GND_net), .O(n19069));   // verilog/coms.v(126[12] 289[6])
    defparam i14037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14038_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n14536), .I3(GND_net), .O(n19070));   // verilog/coms.v(126[12] 289[6])
    defparam i14038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14039_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n14536), .I3(GND_net), .O(n19071));   // verilog/coms.v(126[12] 289[6])
    defparam i14039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14040_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n14536), .I3(GND_net), .O(n19072));   // verilog/coms.v(126[12] 289[6])
    defparam i14040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14041_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n14536), .I3(GND_net), .O(n19073));   // verilog/coms.v(126[12] 289[6])
    defparam i14041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14042_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n14536), .I3(GND_net), .O(n19074));   // verilog/coms.v(126[12] 289[6])
    defparam i14042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14043_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n14536), .I3(GND_net), .O(n19075));   // verilog/coms.v(126[12] 289[6])
    defparam i14043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14044_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n14536), .I3(GND_net), .O(n19076));   // verilog/coms.v(126[12] 289[6])
    defparam i14044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i30_1_lut (.I0(communication_counter[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4940));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13960_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18992));   // verilog/coms.v(126[12] 289[6])
    defparam i13960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13961_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18993));   // verilog/coms.v(126[12] 289[6])
    defparam i13961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4416));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14045_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n14536), .I3(GND_net), .O(n19077));   // verilog/coms.v(126[12] 289[6])
    defparam i14045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14046_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n14536), .I3(GND_net), .O(n19078));   // verilog/coms.v(126[12] 289[6])
    defparam i14046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13962_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18994));   // verilog/coms.v(126[12] 289[6])
    defparam i13962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i31_1_lut (.I0(communication_counter[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4939));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14047_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n14536), .I3(GND_net), .O(n19079));   // verilog/coms.v(126[12] 289[6])
    defparam i14047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i11_3_lut (.I0(communication_counter[10]), .I1(n23_adj_4389), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2558_adj_4508));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_add_2_25_lut (.I0(GND_net), .I1(displacement_23__N_229[23]), 
            .I2(n3_adj_4371), .I3(n30570), .O(displacement_23__N_80[23])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i32_1_lut (.I0(communication_counter[31]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4938));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4415));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14048_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n14536), .I3(GND_net), .O(n19080));   // verilog/coms.v(126[12] 289[6])
    defparam i14048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4414));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_1653_23_lut (.I0(n2471_adj_4574), .I1(n2438), .I2(VCC_net), 
            .I3(n31143), .O(n2537_adj_4573)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1653_22_lut (.I0(GND_net), .I1(n2439), .I2(VCC_net), 
            .I3(n31142), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13797_3_lut (.I0(setpoint[0]), .I1(n4659), .I2(n39863), .I3(GND_net), 
            .O(n18829));   // verilog/coms.v(126[12] 289[6])
    defparam i13797_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1653_22 (.CI(n31142), .I0(n2439), .I1(VCC_net), 
            .CO(n31143));
    SB_LUT4 i13963_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18995));   // verilog/coms.v(126[12] 289[6])
    defparam i13963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1653_21_lut (.I0(GND_net), .I1(n2440), .I2(VCC_net), 
            .I3(n31141), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_21 (.CI(n31141), .I0(n2440), .I1(VCC_net), 
            .CO(n31142));
    SB_LUT4 rem_4_add_1653_20_lut (.I0(GND_net), .I1(n2441), .I2(VCC_net), 
            .I3(n31140), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14049_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n14536), .I3(GND_net), .O(n19081));   // verilog/coms.v(126[12] 289[6])
    defparam i14049_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1653_20 (.CI(n31140), .I0(n2441), .I1(VCC_net), 
            .CO(n31141));
    SB_LUT4 rem_4_add_1653_19_lut (.I0(GND_net), .I1(n2442), .I2(VCC_net), 
            .I3(n31139), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14050_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n14536), .I3(GND_net), .O(n19082));   // verilog/coms.v(126[12] 289[6])
    defparam i14050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14051_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n14536), .I3(GND_net), .O(n19083));   // verilog/coms.v(126[12] 289[6])
    defparam i14051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14052_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n14536), .I3(GND_net), .O(n19084));   // verilog/coms.v(126[12] 289[6])
    defparam i14052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13964_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18996));   // verilog/coms.v(126[12] 289[6])
    defparam i13964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13965_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18997));   // verilog/coms.v(126[12] 289[6])
    defparam i13965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13798_3_lut (.I0(quadB_debounced_adj_4373), .I1(reg_B_adj_5057[0]), 
            .I2(n39886), .I3(GND_net), .O(n18830));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13798_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14053_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n14536), .I3(GND_net), .O(n19085));   // verilog/coms.v(126[12] 289[6])
    defparam i14053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1117_10_lut (.I0(GND_net), .I1(n1651_adj_4486), .I2(VCC_net), 
            .I3(n31380), .O(n1718)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14054_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n14536), .I3(GND_net), .O(n19086));   // verilog/coms.v(126[12] 289[6])
    defparam i14054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14055_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n14536), .I3(GND_net), .O(n19087));   // verilog/coms.v(126[12] 289[6])
    defparam i14055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14396_3_lut (.I0(setpoint[2]), .I1(n4661), .I2(n39863), .I3(GND_net), 
            .O(n19428));   // verilog/coms.v(126[12] 289[6])
    defparam i14396_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14056_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n14536), .I3(GND_net), .O(n19088));   // verilog/coms.v(126[12] 289[6])
    defparam i14056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14057_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n14536), .I3(GND_net), .O(n19089));   // verilog/coms.v(126[12] 289[6])
    defparam i14057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14058_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n14536), .I3(GND_net), .O(n19090));   // verilog/coms.v(126[12] 289[6])
    defparam i14058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14059_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n14536), .I3(GND_net), .O(n19091));   // verilog/coms.v(126[12] 289[6])
    defparam i14059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14060_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n14536), .I3(GND_net), .O(n19092));   // verilog/coms.v(126[12] 289[6])
    defparam i14060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1716_3_lut_3_lut (.I0(n2558), .I1(n7130), .I2(n2551), 
            .I3(GND_net), .O(n2635));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1716_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13966_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18998));   // verilog/coms.v(126[12] 289[6])
    defparam i13966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1699_3_lut_3_lut (.I0(n2558), .I1(n7113), .I2(n2534), 
            .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1699_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut (.I0(control_mode[0]), .I1(n17189), .I2(control_mode[1]), 
            .I3(GND_net), .O(n15_adj_4368));   // verilog/TinyFPGA_B.v(221[5:22])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i14061_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n14536), .I3(GND_net), .O(n19093));   // verilog/coms.v(126[12] 289[6])
    defparam i14061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_add_2_24_lut (.I0(GND_net), .I1(displacement_23__N_229[22]), 
            .I2(n3_adj_4371), .I3(n30569), .O(displacement_23__N_80[22])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_19 (.CI(n31139), .I0(n2442), .I1(VCC_net), 
            .CO(n31140));
    SB_LUT4 rem_4_add_1653_18_lut (.I0(GND_net), .I1(n2443), .I2(VCC_net), 
            .I3(n31138), .O(n2510)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_18 (.CI(n31138), .I0(n2443), .I1(VCC_net), 
            .CO(n31139));
    SB_LUT4 rem_4_add_1653_17_lut (.I0(GND_net), .I1(n2444), .I2(VCC_net), 
            .I3(n31137), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_17 (.CI(n31137), .I0(n2444), .I1(VCC_net), 
            .CO(n31138));
    SB_LUT4 rem_4_add_1653_16_lut (.I0(GND_net), .I1(n2445), .I2(VCC_net), 
            .I3(n31136), .O(n2512)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13967_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18999));   // verilog/coms.v(126[12] 289[6])
    defparam i13967_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1653_16 (.CI(n31136), .I0(n2445), .I1(VCC_net), 
            .CO(n31137));
    SB_LUT4 i14062_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n14536), .I3(GND_net), .O(n19094));   // verilog/coms.v(126[12] 289[6])
    defparam i14062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1653_15_lut (.I0(GND_net), .I1(n2446), .I2(VCC_net), 
            .I3(n31135), .O(n2513)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4413));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1117_10 (.CI(n31380), .I0(n1651_adj_4486), .I1(VCC_net), 
            .CO(n31381));
    SB_LUT4 rem_4_add_1117_9_lut (.I0(GND_net), .I1(n1652_adj_4487), .I2(VCC_net), 
            .I3(n31379), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_9 (.CI(n31379), .I0(n1652_adj_4487), .I1(VCC_net), 
            .CO(n31380));
    SB_CARRY displacement_23__I_0_add_2_24 (.CI(n30569), .I0(displacement_23__N_229[22]), 
            .I1(n3_adj_4371), .CO(n30570));
    SB_LUT4 displacement_23__I_0_add_2_23_lut (.I0(GND_net), .I1(displacement_23__N_229[21]), 
            .I2(n3_adj_4371), .I3(n30568), .O(displacement_23__N_80[21])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_3_lut_adj_1614 (.I0(control_mode[0]), .I1(n17189), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15_adj_4361));   // verilog/TinyFPGA_B.v(221[5:22])
    defparam i1_2_lut_3_lut_adj_1614.LUT_INIT = 16'hefef;
    SB_LUT4 rem_4_add_1117_8_lut (.I0(GND_net), .I1(n1653_adj_4488), .I2(VCC_net), 
            .I3(n31378), .O(n1720)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_8 (.CI(n31378), .I0(n1653_adj_4488), .I1(VCC_net), 
            .CO(n31379));
    SB_LUT4 i13968_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19000));   // verilog/coms.v(126[12] 289[6])
    defparam i13968_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1653_15 (.CI(n31135), .I0(n2446), .I1(VCC_net), 
            .CO(n31136));
    SB_LUT4 div_36_i1700_3_lut_3_lut (.I0(n2558), .I1(n7114), .I2(n2535), 
            .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1700_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1702_3_lut_3_lut (.I0(n2558), .I1(n7116), .I2(n2537), 
            .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1702_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1875_3_lut (.I0(n2754), .I1(n2821_adj_4456), .I2(n2768), 
            .I3(GND_net), .O(n2853));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14063_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n14536), .I3(GND_net), .O(n19095));   // verilog/coms.v(126[12] 289[6])
    defparam i14063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1868_3_lut (.I0(n2747), .I1(n2814), .I2(n2768), .I3(GND_net), 
            .O(n2846));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1868_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY displacement_23__I_0_add_2_23 (.CI(n30568), .I0(displacement_23__N_229[21]), 
            .I1(n3_adj_4371), .CO(n30569));
    SB_LUT4 rem_4_add_1653_14_lut (.I0(GND_net), .I1(n2447_adj_4586), .I2(VCC_net), 
            .I3(n31134), .O(n2514)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_14 (.CI(n31134), .I0(n2447_adj_4586), .I1(VCC_net), 
            .CO(n31135));
    SB_LUT4 rem_4_add_1653_13_lut (.I0(GND_net), .I1(n2448_adj_4585), .I2(VCC_net), 
            .I3(n31133), .O(n2515)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i1701_3_lut_3_lut (.I0(n2558), .I1(n7115), .I2(n2536), 
            .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1701_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1871_3_lut (.I0(n2750), .I1(n2817_adj_4460), .I2(n2768), 
            .I3(GND_net), .O(n2849));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1869_3_lut (.I0(n2748), .I1(n2815), .I2(n2768), .I3(GND_net), 
            .O(n2847));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1869_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1870_3_lut (.I0(n2749), .I1(n2816_adj_4461), .I2(n2768), 
            .I3(GND_net), .O(n2848));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1861_3_lut (.I0(n2740), .I1(n2807), .I2(n2768), .I3(GND_net), 
            .O(n2839_adj_4446));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1859_3_lut (.I0(n2738), .I1(n2805), .I2(n2768), .I3(GND_net), 
            .O(n2837_adj_4448));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1860_3_lut (.I0(n2739), .I1(n2806), .I2(n2768), .I3(GND_net), 
            .O(n2838_adj_4447));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1858_3_lut (.I0(n2737), .I1(n2804), .I2(n2768), .I3(GND_net), 
            .O(n2836_adj_4449));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14064_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n14536), .I3(GND_net), .O(n19096));   // verilog/coms.v(126[12] 289[6])
    defparam i14064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1865_3_lut (.I0(n2744), .I1(n2811), .I2(n2768), .I3(GND_net), 
            .O(n2843));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1865_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1863_3_lut (.I0(n2742), .I1(n2809), .I2(n2768), .I3(GND_net), 
            .O(n2841));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1117_7_lut (.I0(GND_net), .I1(n1654), .I2(GND_net), 
            .I3(n31377), .O(n1721)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_13 (.CI(n31133), .I0(n2448_adj_4585), .I1(VCC_net), 
            .CO(n31134));
    SB_CARRY rem_4_add_1117_7 (.CI(n31377), .I0(n1654), .I1(GND_net), 
            .CO(n31378));
    SB_LUT4 rem_4_add_1653_12_lut (.I0(GND_net), .I1(n2449_adj_4584), .I2(VCC_net), 
            .I3(n31132), .O(n2516)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1117_6_lut (.I0(GND_net), .I1(n1655), .I2(GND_net), 
            .I3(n31376), .O(n1722)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_6 (.CI(n31376), .I0(n1655), .I1(GND_net), 
            .CO(n31377));
    SB_CARRY rem_4_add_1653_12 (.CI(n31132), .I0(n2449_adj_4584), .I1(VCC_net), 
            .CO(n31133));
    SB_LUT4 rem_4_add_1117_5_lut (.I0(GND_net), .I1(n1656), .I2(VCC_net), 
            .I3(n31375), .O(n1723)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4345));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1864_3_lut (.I0(n2743), .I1(n2810), .I2(n2768), .I3(GND_net), 
            .O(n2842));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1862_3_lut (.I0(n2741), .I1(n2808), .I2(n2768), .I3(GND_net), 
            .O(n2840));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1877_3_lut (.I0(n2756), .I1(n2823_adj_4454), .I2(n2768), 
            .I3(GND_net), .O(n2855));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1866_3_lut (.I0(n2745), .I1(n2812), .I2(n2768), .I3(GND_net), 
            .O(n2844));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1866_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1876_3_lut (.I0(n2755), .I1(n2822_adj_4455), .I2(n2768), 
            .I3(GND_net), .O(n2854));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1874_3_lut (.I0(n2753), .I1(n2820_adj_4457), .I2(n2768), 
            .I3(GND_net), .O(n2852));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1874_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1873_3_lut (.I0(n2752), .I1(n2819_adj_4458), .I2(n2768), 
            .I3(GND_net), .O(n2851));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1873_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1653_11_lut (.I0(GND_net), .I1(n2450_adj_4583), .I2(VCC_net), 
            .I3(n31131), .O(n2517)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1872_3_lut (.I0(n2751), .I1(n2818_adj_4459), .I2(n2768), 
            .I3(GND_net), .O(n2850));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1872_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1653_11 (.CI(n31131), .I0(n2450_adj_4583), .I1(VCC_net), 
            .CO(n31132));
    SB_LUT4 rem_4_i1867_3_lut (.I0(n2746), .I1(n2813), .I2(n2768), .I3(GND_net), 
            .O(n2845));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1653_10_lut (.I0(GND_net), .I1(n2451_adj_4582), .I2(VCC_net), 
            .I3(n31130), .O(n2518)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_5 (.CI(n31375), .I0(n1656), .I1(VCC_net), 
            .CO(n31376));
    SB_LUT4 rem_4_i1879_3_lut (.I0(n2758), .I1(n2825_adj_4452), .I2(n2768), 
            .I3(GND_net), .O(n2857_adj_4442));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1878_3_lut (.I0(n2757), .I1(n2824_adj_4453), .I2(n2768), 
            .I3(GND_net), .O(n2856));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1117_4_lut (.I0(GND_net), .I1(n1657), .I2(VCC_net), 
            .I3(n31374), .O(n1724)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1857_3_lut (.I0(n2736), .I1(n2803), .I2(n2768), .I3(GND_net), 
            .O(n2835_adj_4450));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(n2835_adj_4450), .I1(n2834_adj_4451), .I2(GND_net), 
            .I3(GND_net), .O(n22_adj_4934));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 displacement_23__I_0_add_2_22_lut (.I0(GND_net), .I1(displacement_23__N_229[20]), 
            .I2(n3_adj_4371), .I3(n30567), .O(displacement_23__N_80[20])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_4 (.CI(n31374), .I0(n1657), .I1(VCC_net), 
            .CO(n31375));
    SB_LUT4 i14065_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n14536), .I3(GND_net), .O(n19097));   // verilog/coms.v(126[12] 289[6])
    defparam i14065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14066_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n14536), 
            .I3(GND_net), .O(n19098));   // verilog/coms.v(126[12] 289[6])
    defparam i14066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14067_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n14536), 
            .I3(GND_net), .O(n19099));   // verilog/coms.v(126[12] 289[6])
    defparam i14067_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY displacement_23__I_0_add_2_22 (.CI(n30567), .I0(displacement_23__N_229[20]), 
            .I1(n3_adj_4371), .CO(n30568));
    SB_LUT4 i1_3_lut_adj_1615 (.I0(n2856), .I1(n2857_adj_4442), .I2(n2858), 
            .I3(GND_net), .O(n38397));
    defparam i1_3_lut_adj_1615.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_add_1117_3_lut (.I0(GND_net), .I1(n1658), .I2(GND_net), 
            .I3(n31373), .O(n1725)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_21_lut (.I0(GND_net), .I1(displacement_23__N_229[19]), 
            .I2(n6_adj_4345), .I3(n30566), .O(displacement_23__N_80[19])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_10 (.CI(n31130), .I0(n2451_adj_4582), .I1(VCC_net), 
            .CO(n31131));
    SB_CARRY displacement_23__I_0_add_2_21 (.CI(n30566), .I0(displacement_23__N_229[19]), 
            .I1(n6_adj_4345), .CO(n30567));
    SB_CARRY rem_4_add_1117_3 (.CI(n31373), .I0(n1658), .I1(GND_net), 
            .CO(n31374));
    SB_LUT4 displacement_23__I_0_add_2_20_lut (.I0(GND_net), .I1(displacement_23__N_229[18]), 
            .I2(n7), .I3(n30565), .O(displacement_23__N_80[18])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_20 (.CI(n30565), .I0(displacement_23__N_229[18]), 
            .I1(n7), .CO(n30566));
    SB_LUT4 i15_4_lut (.I0(n2845), .I1(n2850), .I2(n2851), .I3(n2852), 
            .O(n36_adj_4930));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(n2854), .I1(n2844), .I2(n38397), .I3(n2855), 
            .O(n27_adj_4933));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i6_4_lut.LUT_INIT = 16'heccc;
    SB_CARRY rem_4_add_1117_2 (.CI(VCC_net), .I0(n1758_adj_4781), .I1(VCC_net), 
            .CO(n31373));
    SB_IO PIN_2_pad (.PACKAGE_PIN(PIN_2), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_2_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_2_pad.PIN_TYPE = 6'b000001;
    defparam PIN_2_pad.PULLUP = 1'b0;
    defparam PIN_2_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_2_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i13_4_lut_adj_1616 (.I0(n2840), .I1(n2842), .I2(n2841), .I3(n2843), 
            .O(n34_adj_4931));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i13_4_lut_adj_1616.LUT_INIT = 16'hfffe;
    SB_LUT4 displacement_23__I_0_add_2_19_lut (.I0(GND_net), .I1(displacement_23__N_229[17]), 
            .I2(n8_adj_4413), .I3(n30564), .O(displacement_23__N_80[17])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_16_lut (.I0(n1778_adj_4738), .I1(n1745), .I2(VCC_net), 
            .I3(n31372), .O(n1844)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i12_4_lut_adj_1617 (.I0(n2836_adj_4449), .I1(n2838_adj_4447), 
            .I2(n2837_adj_4448), .I3(n2839_adj_4446), .O(n33_adj_4932));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i12_4_lut_adj_1617.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1618 (.I0(n2849), .I1(n2846), .I2(n2853), .I3(n22_adj_4934), 
            .O(n37_adj_4929));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i16_4_lut_adj_1618.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(n27_adj_4933), .I1(n36_adj_4930), .I2(n2848), 
            .I3(n2847), .O(n39_adj_4928));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut (.I0(n39_adj_4928), .I1(n37_adj_4929), .I2(n33_adj_4932), 
            .I3(n34_adj_4931), .O(n2867_adj_4441));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i8_3_lut (.I0(communication_counter[7]), .I1(n26), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2858));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1719_3_lut_3_lut (.I0(n2558), .I1(n7133), .I2(n388), 
            .I3(GND_net), .O(n2638));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1705_3_lut_3_lut (.I0(n2558), .I1(n7119), .I2(n2540), 
            .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1705_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1184_15_lut (.I0(GND_net), .I1(n1746), .I2(VCC_net), 
            .I3(n31371), .O(n1813)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_9_lut (.I0(GND_net), .I1(n2452_adj_4581), .I2(VCC_net), 
            .I3(n31129), .O(n2519)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_15 (.CI(n31371), .I0(n1746), .I1(VCC_net), 
            .CO(n31372));
    SB_CARRY displacement_23__I_0_add_2_19 (.CI(n30564), .I0(displacement_23__N_229[17]), 
            .I1(n8_adj_4413), .CO(n30565));
    SB_LUT4 rem_4_add_1184_14_lut (.I0(GND_net), .I1(n1747), .I2(VCC_net), 
            .I3(n31370), .O(n1814)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_14 (.CI(n31370), .I0(n1747), .I1(VCC_net), 
            .CO(n31371));
    SB_CARRY rem_4_add_1653_9 (.CI(n31129), .I0(n2452_adj_4581), .I1(VCC_net), 
            .CO(n31130));
    SB_LUT4 rem_4_add_1653_8_lut (.I0(GND_net), .I1(n2453_adj_4580), .I2(VCC_net), 
            .I3(n31128), .O(n2520)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_8 (.CI(n31128), .I0(n2453_adj_4580), .I1(VCC_net), 
            .CO(n31129));
    SB_LUT4 rem_4_add_1184_13_lut (.I0(GND_net), .I1(n1748), .I2(VCC_net), 
            .I3(n31369), .O(n1815)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14068_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n14536), 
            .I3(GND_net), .O(n19100));   // verilog/coms.v(126[12] 289[6])
    defparam i14068_3_lut.LUT_INIT = 16'hcaca;
    SB_IO PIN_1_pad (.PACKAGE_PIN(PIN_1), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_1_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_1_pad.PIN_TYPE = 6'b000001;
    defparam PIN_1_pad.PULLUP = 1'b0;
    defparam PIN_1_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_24_pad (.PACKAGE_PIN(PIN_24), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_24_pad.PIN_TYPE = 6'b011001;
    defparam PIN_24_pad.PULLUP = 1'b0;
    defparam PIN_24_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_23_pad (.PACKAGE_PIN(PIN_23), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_23_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_23_pad.PIN_TYPE = 6'b011001;
    defparam PIN_23_pad.PULLUP = 1'b0;
    defparam PIN_23_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_7_pad (.PACKAGE_PIN(PIN_7), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_7_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_7_pad.PIN_TYPE = 6'b000001;
    defparam PIN_7_pad.PULLUP = 1'b0;
    defparam PIN_7_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_36_i1706_3_lut_3_lut (.I0(n2558), .I1(n7120), .I2(n2541), 
            .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1706_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1184_13 (.CI(n31369), .I0(n1748), .I1(VCC_net), 
            .CO(n31370));
    SB_LUT4 rem_4_add_1653_7_lut (.I0(GND_net), .I1(n2454_adj_4579), .I2(GND_net), 
            .I3(n31127), .O(n2521)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_7 (.CI(n31127), .I0(n2454_adj_4579), .I1(GND_net), 
            .CO(n31128));
    SB_LUT4 rem_4_add_1184_12_lut (.I0(GND_net), .I1(n1749), .I2(VCC_net), 
            .I3(n31368), .O(n1816)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_12 (.CI(n31368), .I0(n1749), .I1(VCC_net), 
            .CO(n31369));
    SB_LUT4 rem_4_add_1184_11_lut (.I0(GND_net), .I1(n1750), .I2(VCC_net), 
            .I3(n31367), .O(n1817)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14238_3_lut (.I0(\data_in_frame[15] [5]), .I1(rx_data[5]), 
            .I2(n37348), .I3(GND_net), .O(n19270));   // verilog/coms.v(126[12] 289[6])
    defparam i14238_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1184_11 (.CI(n31367), .I0(n1750), .I1(VCC_net), 
            .CO(n31368));
    SB_LUT4 rem_4_add_1653_6_lut (.I0(GND_net), .I1(n2455_adj_4578), .I2(GND_net), 
            .I3(n31126), .O(n2522)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_6 (.CI(n31126), .I0(n2455_adj_4578), .I1(GND_net), 
            .CO(n31127));
    SB_LUT4 rem_4_add_1653_5_lut (.I0(GND_net), .I1(n2456_adj_4577), .I2(VCC_net), 
            .I3(n31125), .O(n2523)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_10_lut (.I0(GND_net), .I1(n1751), .I2(VCC_net), 
            .I3(n31366), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_10 (.CI(n31366), .I0(n1751), .I1(VCC_net), 
            .CO(n31367));
    SB_LUT4 rem_4_add_1184_9_lut (.I0(GND_net), .I1(n1752), .I2(VCC_net), 
            .I3(n31365), .O(n1819)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_9 (.CI(n31365), .I0(n1752), .I1(VCC_net), 
            .CO(n31366));
    SB_LUT4 rem_4_add_1184_8_lut (.I0(GND_net), .I1(n1753), .I2(VCC_net), 
            .I3(n31364), .O(n1820)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i1708_3_lut_3_lut (.I0(n2558), .I1(n7122), .I2(n2543), 
            .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1708_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_3_lut_adj_1619 (.I0(n37219), .I1(r_Clock_Count[2]), .I2(n16_adj_4990), 
            .I3(GND_net), .O(n36985));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_1619.LUT_INIT = 16'heaea;
    SB_LUT4 div_36_i1709_3_lut_3_lut (.I0(n2558), .I1(n7123), .I2(n2544), 
            .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1709_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_add_2_18_lut (.I0(GND_net), .I1(displacement_23__N_229[16]), 
            .I2(n9_adj_4414), .I3(n30563), .O(displacement_23__N_80[16])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_8 (.CI(n31364), .I0(n1753), .I1(VCC_net), 
            .CO(n31365));
    SB_CARRY displacement_23__I_0_add_2_18 (.CI(n30563), .I0(displacement_23__N_229[16]), 
            .I1(n9_adj_4414), .CO(n30564));
    SB_LUT4 rem_4_add_1184_7_lut (.I0(GND_net), .I1(n1754_adj_4785), .I2(GND_net), 
            .I3(n31363), .O(n1821)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_7 (.CI(n31363), .I0(n1754_adj_4785), .I1(GND_net), 
            .CO(n31364));
    SB_LUT4 displacement_23__I_0_add_2_17_lut (.I0(GND_net), .I1(displacement_23__N_229[15]), 
            .I2(n10_adj_4415), .I3(n30562), .O(displacement_23__N_80[15])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_5 (.CI(n31125), .I0(n2456_adj_4577), .I1(VCC_net), 
            .CO(n31126));
    SB_CARRY displacement_23__I_0_add_2_17 (.CI(n30562), .I0(displacement_23__N_229[15]), 
            .I1(n10_adj_4415), .CO(n30563));
    SB_LUT4 rem_4_add_1653_4_lut (.I0(GND_net), .I1(n2457_adj_4576), .I2(VCC_net), 
            .I3(n31124), .O(n2524)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_4 (.CI(n31124), .I0(n2457_adj_4576), .I1(VCC_net), 
            .CO(n31125));
    SB_LUT4 rem_4_add_1184_6_lut (.I0(GND_net), .I1(n1755_adj_4784), .I2(GND_net), 
            .I3(n31362), .O(n1822)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_3_lut (.I0(GND_net), .I1(n2458_adj_4575), .I2(GND_net), 
            .I3(n31123), .O(n2525)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_3 (.CI(n31123), .I0(n2458_adj_4575), .I1(GND_net), 
            .CO(n31124));
    SB_CARRY rem_4_add_1653_2 (.CI(VCC_net), .I0(n2558_adj_4508), .I1(VCC_net), 
            .CO(n31123));
    SB_LUT4 communication_counter_1146_add_4_33_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[31]), .I3(n31122), .O(n134)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_6 (.CI(n31362), .I0(n1755_adj_4784), .I1(GND_net), 
            .CO(n31363));
    SB_LUT4 rem_4_add_1184_5_lut (.I0(GND_net), .I1(n1756_adj_4783), .I2(VCC_net), 
            .I3(n31361), .O(n1823)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1146_add_4_32_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[30]), .I3(n31121), .O(n135)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13969_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19001));   // verilog/coms.v(126[12] 289[6])
    defparam i13969_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1146_add_4_32 (.CI(n31121), .I0(GND_net), 
            .I1(communication_counter[30]), .CO(n31122));
    SB_LUT4 communication_counter_1146_add_4_31_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[29]), .I3(n31120), .O(n136)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i1710_3_lut_3_lut (.I0(n2558), .I1(n7124), .I2(n2545), 
            .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1710_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i33753_1_lut (.I0(n40223), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n40287));
    defparam i33753_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY communication_counter_1146_add_4_31 (.CI(n31120), .I0(GND_net), 
            .I1(communication_counter[29]), .CO(n31121));
    SB_LUT4 i14239_3_lut (.I0(\data_in_frame[15] [6]), .I1(rx_data[6]), 
            .I2(n37348), .I3(GND_net), .O(n19271));   // verilog/coms.v(126[12] 289[6])
    defparam i14239_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1184_5 (.CI(n31361), .I0(n1756_adj_4783), .I1(VCC_net), 
            .CO(n31362));
    SB_LUT4 displacement_23__I_0_add_2_16_lut (.I0(GND_net), .I1(displacement_23__N_229[14]), 
            .I2(n11_adj_4416), .I3(n30561), .O(displacement_23__N_80[14])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_4_lut (.I0(GND_net), .I1(n1757_adj_4782), .I2(VCC_net), 
            .I3(n31360), .O(n1824)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1146_add_4_30_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[28]), .I3(n31119), .O(n137)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1146_add_4_30 (.CI(n31119), .I0(GND_net), 
            .I1(communication_counter[28]), .CO(n31120));
    SB_LUT4 communication_counter_1146_add_4_29_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[27]), .I3(n31118), .O(n138)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_4 (.CI(n31360), .I0(n1757_adj_4782), .I1(VCC_net), 
            .CO(n31361));
    SB_CARRY communication_counter_1146_add_4_29 (.CI(n31118), .I0(GND_net), 
            .I1(communication_counter[27]), .CO(n31119));
    SB_LUT4 communication_counter_1146_add_4_28_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[26]), .I3(n31117), .O(n139)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1146_add_4_28 (.CI(n31117), .I0(GND_net), 
            .I1(communication_counter[26]), .CO(n31118));
    SB_LUT4 rem_4_add_1184_3_lut (.I0(GND_net), .I1(n1758_adj_4781), .I2(GND_net), 
            .I3(n31359), .O(n1825)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1146_add_4_27_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[25]), .I3(n31116), .O(n140)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_3 (.CI(n31359), .I0(n1758_adj_4781), .I1(GND_net), 
            .CO(n31360));
    SB_CARRY communication_counter_1146_add_4_27 (.CI(n31116), .I0(GND_net), 
            .I1(communication_counter[25]), .CO(n31117));
    SB_LUT4 communication_counter_1146_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[24]), .I3(n31115), .O(n141)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 PIN_13_I_0_1_lut (.I0(PIN_13_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(PIN_13_N_105));   // verilog/TinyFPGA_B.v(200[10:15])
    defparam PIN_13_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY communication_counter_1146_add_4_26 (.CI(n31115), .I0(GND_net), 
            .I1(communication_counter[24]), .CO(n31116));
    SB_CARRY rem_4_add_1184_2 (.CI(VCC_net), .I0(n1858), .I1(VCC_net), 
            .CO(n31359));
    SB_LUT4 communication_counter_1146_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[23]), .I3(n31114), .O(n142)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1146_add_4_25 (.CI(n31114), .I0(GND_net), 
            .I1(communication_counter[23]), .CO(n31115));
    SB_LUT4 communication_counter_1146_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[22]), .I3(n31113), .O(n143)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_17_lut (.I0(n1877), .I1(n1844), .I2(VCC_net), 
            .I3(n31358), .O(n1943)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY communication_counter_1146_add_4_24 (.CI(n31113), .I0(GND_net), 
            .I1(communication_counter[22]), .CO(n31114));
    SB_LUT4 i13970_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19002));   // verilog/coms.v(126[12] 289[6])
    defparam i13970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1146_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[21]), .I3(n31112), .O(n144)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_16 (.CI(n30561), .I0(displacement_23__N_229[14]), 
            .I1(n11_adj_4416), .CO(n30562));
    SB_CARRY communication_counter_1146_add_4_23 (.CI(n31112), .I0(GND_net), 
            .I1(communication_counter[21]), .CO(n31113));
    SB_LUT4 communication_counter_1146_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[20]), .I3(n31111), .O(n145)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1146_add_4_22 (.CI(n31111), .I0(GND_net), 
            .I1(communication_counter[20]), .CO(n31112));
    SB_LUT4 rem_4_add_1251_16_lut (.I0(GND_net), .I1(n1845), .I2(VCC_net), 
            .I3(n31357), .O(n1912)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_16 (.CI(n31357), .I0(n1845), .I1(VCC_net), 
            .CO(n31358));
    SB_LUT4 rem_4_add_1251_15_lut (.I0(GND_net), .I1(n1846), .I2(VCC_net), 
            .I3(n31356), .O(n1913)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1146_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[19]), .I3(n31110), .O(n146)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_15 (.CI(n31356), .I0(n1846), .I1(VCC_net), 
            .CO(n31357));
    SB_LUT4 i14240_3_lut (.I0(\data_in_frame[15] [7]), .I1(rx_data[7]), 
            .I2(n37348), .I3(GND_net), .O(n19272));   // verilog/coms.v(126[12] 289[6])
    defparam i14240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1251_14_lut (.I0(GND_net), .I1(n1847), .I2(VCC_net), 
            .I3(n31355), .O(n1914)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1146_add_4_21 (.CI(n31110), .I0(GND_net), 
            .I1(communication_counter[19]), .CO(n31111));
    SB_CARRY rem_4_add_1251_14 (.CI(n31355), .I0(n1847), .I1(VCC_net), 
            .CO(n31356));
    SB_LUT4 i13971_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19003));   // verilog/coms.v(126[12] 289[6])
    defparam i13971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1251_13_lut (.I0(GND_net), .I1(n1848), .I2(VCC_net), 
            .I3(n31354), .O(n1915)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1146_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[18]), .I3(n31109), .O(n147)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_13 (.CI(n31354), .I0(n1848), .I1(VCC_net), 
            .CO(n31355));
    SB_CARRY communication_counter_1146_add_4_20 (.CI(n31109), .I0(GND_net), 
            .I1(communication_counter[18]), .CO(n31110));
    SB_LUT4 rem_4_add_1251_12_lut (.I0(GND_net), .I1(n1849), .I2(VCC_net), 
            .I3(n31353), .O(n1916)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_12_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_21_pad (.PACKAGE_PIN(PIN_21), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_21_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_21_pad.PIN_TYPE = 6'b011001;
    defparam PIN_21_pad.PULLUP = 1'b0;
    defparam PIN_21_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY rem_4_add_1251_12 (.CI(n31353), .I0(n1849), .I1(VCC_net), 
            .CO(n31354));
    SB_LUT4 rem_4_add_1251_11_lut (.I0(GND_net), .I1(n1850), .I2(VCC_net), 
            .I3(n31352), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1146_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[17]), .I3(n31108), .O(n148)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_20_pad (.PACKAGE_PIN(PIN_20), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_20_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_20_pad.PIN_TYPE = 6'b011001;
    defparam PIN_20_pad.PULLUP = 1'b0;
    defparam PIN_20_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY communication_counter_1146_add_4_19 (.CI(n31108), .I0(GND_net), 
            .I1(communication_counter[17]), .CO(n31109));
    SB_LUT4 communication_counter_1146_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[16]), .I3(n31107), .O(n149)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1146_add_4_18 (.CI(n31107), .I0(GND_net), 
            .I1(communication_counter[16]), .CO(n31108));
    SB_LUT4 communication_counter_1146_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[15]), .I3(n31106), .O(n150)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i1711_3_lut_3_lut (.I0(n2558), .I1(n7125), .I2(n2546), 
            .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1711_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1251_11 (.CI(n31352), .I0(n1850), .I1(VCC_net), 
            .CO(n31353));
    SB_CARRY communication_counter_1146_add_4_17 (.CI(n31106), .I0(GND_net), 
            .I1(communication_counter[15]), .CO(n31107));
    SB_LUT4 communication_counter_1146_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[14]), .I3(n31105), .O(n151)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_10_lut (.I0(GND_net), .I1(n1851), .I2(VCC_net), 
            .I3(n31351), .O(n1918)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_10 (.CI(n31351), .I0(n1851), .I1(VCC_net), 
            .CO(n31352));
    SB_CARRY communication_counter_1146_add_4_16 (.CI(n31105), .I0(GND_net), 
            .I1(communication_counter[14]), .CO(n31106));
    SB_LUT4 displacement_23__I_0_add_2_15_lut (.I0(GND_net), .I1(displacement_23__N_229[13]), 
            .I2(n12_adj_4417), .I3(n30560), .O(displacement_23__N_80[13])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_9_lut (.I0(GND_net), .I1(n1852), .I2(VCC_net), 
            .I3(n31350), .O(n1919)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_9 (.CI(n31350), .I0(n1852), .I1(VCC_net), 
            .CO(n31351));
    SB_LUT4 communication_counter_1146_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[13]), .I3(n31104), .O(n152)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1146_add_4_15 (.CI(n31104), .I0(GND_net), 
            .I1(communication_counter[13]), .CO(n31105));
    SB_LUT4 i13972_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19004));   // verilog/coms.v(126[12] 289[6])
    defparam i13972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1146_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[12]), .I3(n31103), .O(n153)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_8_lut (.I0(GND_net), .I1(n1853), .I2(VCC_net), 
            .I3(n31349), .O(n1920)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_8 (.CI(n31349), .I0(n1853), .I1(VCC_net), 
            .CO(n31350));
    SB_LUT4 rem_4_add_1251_7_lut (.I0(GND_net), .I1(n1854), .I2(GND_net), 
            .I3(n31348), .O(n1921)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_7 (.CI(n31348), .I0(n1854), .I1(GND_net), 
            .CO(n31349));
    SB_CARRY communication_counter_1146_add_4_14 (.CI(n31103), .I0(GND_net), 
            .I1(communication_counter[12]), .CO(n31104));
    SB_LUT4 communication_counter_1146_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[11]), .I3(n31102), .O(n154)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_6_lut (.I0(GND_net), .I1(n1855), .I2(GND_net), 
            .I3(n31347), .O(n1922)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_6 (.CI(n31347), .I0(n1855), .I1(GND_net), 
            .CO(n31348));
    SB_LUT4 rem_4_add_1251_5_lut (.I0(GND_net), .I1(n1856), .I2(VCC_net), 
            .I3(n31346), .O(n1923)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_5 (.CI(n31346), .I0(n1856), .I1(VCC_net), 
            .CO(n31347));
    SB_LUT4 i14069_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n14536), 
            .I3(GND_net), .O(n19101));   // verilog/coms.v(126[12] 289[6])
    defparam i14069_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1146_add_4_13 (.CI(n31102), .I0(GND_net), 
            .I1(communication_counter[11]), .CO(n31103));
    SB_LUT4 communication_counter_1146_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[10]), .I3(n31101), .O(n155)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1146_add_4_12 (.CI(n31101), .I0(GND_net), 
            .I1(communication_counter[10]), .CO(n31102));
    SB_LUT4 communication_counter_1146_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[9]), .I3(n31100), .O(n156)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1146_add_4_11 (.CI(n31100), .I0(GND_net), 
            .I1(communication_counter[9]), .CO(n31101));
    SB_LUT4 communication_counter_1146_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[8]), .I3(n31099), .O(n157)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_4_lut (.I0(GND_net), .I1(n1857), .I2(VCC_net), 
            .I3(n31345), .O(n1924)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_4 (.CI(n31345), .I0(n1857), .I1(VCC_net), 
            .CO(n31346));
    SB_LUT4 rem_4_add_1251_3_lut (.I0(GND_net), .I1(n1858), .I2(GND_net), 
            .I3(n31344), .O(n1925)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1146_add_4_10 (.CI(n31099), .I0(GND_net), 
            .I1(communication_counter[8]), .CO(n31100));
    SB_LUT4 communication_counter_1146_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[7]), .I3(n31098), .O(n158)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1146_add_4_9 (.CI(n31098), .I0(GND_net), 
            .I1(communication_counter[7]), .CO(n31099));
    SB_LUT4 communication_counter_1146_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[6]), .I3(n31097), .O(n159)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_3 (.CI(n31344), .I0(n1858), .I1(GND_net), 
            .CO(n31345));
    SB_CARRY communication_counter_1146_add_4_8 (.CI(n31097), .I0(GND_net), 
            .I1(communication_counter[6]), .CO(n31098));
    SB_LUT4 communication_counter_1146_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[5]), .I3(n31096), .O(n160)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1146_add_4_7 (.CI(n31096), .I0(GND_net), 
            .I1(communication_counter[5]), .CO(n31097));
    SB_LUT4 communication_counter_1146_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[4]), .I3(n31095), .O(n161)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1146_add_4_6 (.CI(n31095), .I0(GND_net), 
            .I1(communication_counter[4]), .CO(n31096));
    SB_LUT4 communication_counter_1146_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[3]), .I3(n31094), .O(n162)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1146_add_4_5 (.CI(n31094), .I0(GND_net), 
            .I1(communication_counter[3]), .CO(n31095));
    SB_LUT4 div_36_i1717_3_lut_3_lut (.I0(n2558), .I1(n7131), .I2(n2552), 
            .I3(GND_net), .O(n2636));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1717_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1251_2 (.CI(VCC_net), .I0(n1958), .I1(VCC_net), 
            .CO(n31344));
    SB_CARRY displacement_23__I_0_add_2_15 (.CI(n30560), .I0(displacement_23__N_229[13]), 
            .I1(n12_adj_4417), .CO(n30561));
    SB_LUT4 i13973_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19005));   // verilog/coms.v(126[12] 289[6])
    defparam i13973_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF h1_45 (.Q(PIN_20_c), .C(clk32MHz), .D(hall1));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_LUT4 i13974_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19006));   // verilog/coms.v(126[12] 289[6])
    defparam i13974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_add_2_14_lut (.I0(GND_net), .I1(displacement_23__N_229[12]), 
            .I2(n13_adj_4418), .I3(n30559), .O(displacement_23__N_80[12])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1146_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[2]), .I3(n31093), .O(n163)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1146_add_4_4 (.CI(n31093), .I0(GND_net), 
            .I1(communication_counter[2]), .CO(n31094));
    SB_LUT4 rem_4_add_1318_18_lut (.I0(n1976_adj_4627), .I1(n1943), .I2(VCC_net), 
            .I3(n31343), .O(n2042)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 communication_counter_1146_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[1]), .I3(n31092), .O(n164)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1318_17_lut (.I0(GND_net), .I1(n1944), .I2(VCC_net), 
            .I3(n31342), .O(n2011)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1146_add_4_3 (.CI(n31092), .I0(GND_net), 
            .I1(communication_counter[1]), .CO(n31093));
    SB_LUT4 i13975_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19007));   // verilog/coms.v(126[12] 289[6])
    defparam i13975_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1318_17 (.CI(n31342), .I0(n1944), .I1(VCC_net), 
            .CO(n31343));
    SB_LUT4 i13976_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19008));   // verilog/coms.v(126[12] 289[6])
    defparam i13976_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY displacement_23__I_0_add_2_14 (.CI(n30559), .I0(displacement_23__N_229[12]), 
            .I1(n13_adj_4418), .CO(n30560));
    SB_LUT4 communication_counter_1146_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[0]), .I3(VCC_net), .O(n165)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1146_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1146_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(communication_counter[0]), .CO(n31092));
    SB_LUT4 rem_4_add_1720_24_lut (.I0(n2570), .I1(n2537_adj_4573), .I2(VCC_net), 
            .I3(n31091), .O(n2636_adj_4495)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1720_23_lut (.I0(GND_net), .I1(n2538_adj_4572), .I2(VCC_net), 
            .I3(n31090), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_23 (.CI(n31090), .I0(n2538_adj_4572), .I1(VCC_net), 
            .CO(n31091));
    SB_LUT4 displacement_23__I_0_add_2_13_lut (.I0(GND_net), .I1(displacement_23__N_229[11]), 
            .I2(n14_adj_4419), .I3(n30558), .O(displacement_23__N_80[11])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_22_lut (.I0(GND_net), .I1(n2539_adj_4571), .I2(VCC_net), 
            .I3(n31089), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_22 (.CI(n31089), .I0(n2539_adj_4571), .I1(VCC_net), 
            .CO(n31090));
    SB_LUT4 rem_4_add_1318_16_lut (.I0(GND_net), .I1(n1945), .I2(VCC_net), 
            .I3(n31341), .O(n2012)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_16_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_80[23]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_LUT4 rem_4_add_1720_21_lut (.I0(GND_net), .I1(n2540_adj_4570), .I2(VCC_net), 
            .I3(n31088), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_16 (.CI(n31341), .I0(n1945), .I1(VCC_net), 
            .CO(n31342));
    SB_LUT4 rem_4_add_1318_15_lut (.I0(GND_net), .I1(n1946), .I2(VCC_net), 
            .I3(n31340), .O(n2013)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_13 (.CI(n30558), .I0(displacement_23__N_229[11]), 
            .I1(n14_adj_4419), .CO(n30559));
    SB_CARRY rem_4_add_1318_15 (.CI(n31340), .I0(n1946), .I1(VCC_net), 
            .CO(n31341));
    SB_LUT4 rem_4_add_1318_14_lut (.I0(GND_net), .I1(n1947), .I2(VCC_net), 
            .I3(n31339), .O(n2014)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_21 (.CI(n31088), .I0(n2540_adj_4570), .I1(VCC_net), 
            .CO(n31089));
    SB_LUT4 rem_4_add_1720_20_lut (.I0(GND_net), .I1(n2541_adj_4569), .I2(VCC_net), 
            .I3(n31087), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_12_lut (.I0(GND_net), .I1(displacement_23__N_229[10]), 
            .I2(n15_adj_4420), .I3(n30557), .O(displacement_23__N_80[10])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_14 (.CI(n31339), .I0(n1947), .I1(VCC_net), 
            .CO(n31340));
    SB_CARRY rem_4_add_1720_20 (.CI(n31087), .I0(n2541_adj_4569), .I1(VCC_net), 
            .CO(n31088));
    SB_LUT4 rem_4_add_1720_19_lut (.I0(GND_net), .I1(n2542_adj_4520), .I2(VCC_net), 
            .I3(n31086), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1318_13_lut (.I0(GND_net), .I1(n1948), .I2(VCC_net), 
            .I3(n31338), .O(n2015)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_19 (.CI(n31086), .I0(n2542_adj_4520), .I1(VCC_net), 
            .CO(n31087));
    SB_LUT4 rem_4_add_1720_18_lut (.I0(GND_net), .I1(n2543_adj_4519), .I2(VCC_net), 
            .I3(n31085), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_18 (.CI(n31085), .I0(n2543_adj_4519), .I1(VCC_net), 
            .CO(n31086));
    SB_LUT4 rem_4_add_1720_17_lut (.I0(GND_net), .I1(n2544_adj_4518), .I2(VCC_net), 
            .I3(n31084), .O(n2611)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_13 (.CI(n31338), .I0(n1948), .I1(VCC_net), 
            .CO(n31339));
    SB_CARRY rem_4_add_1720_17 (.CI(n31084), .I0(n2544_adj_4518), .I1(VCC_net), 
            .CO(n31085));
    SB_LUT4 rem_4_add_1720_16_lut (.I0(GND_net), .I1(n2545_adj_4517), .I2(VCC_net), 
            .I3(n31083), .O(n2612)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_16 (.CI(n31083), .I0(n2545_adj_4517), .I1(VCC_net), 
            .CO(n31084));
    SB_LUT4 rem_4_add_1720_15_lut (.I0(GND_net), .I1(n2546_adj_4516), .I2(VCC_net), 
            .I3(n31082), .O(n2613)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1318_12_lut (.I0(GND_net), .I1(n1949), .I2(VCC_net), 
            .I3(n31337), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13977_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19009));   // verilog/coms.v(126[12] 289[6])
    defparam i13977_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY displacement_23__I_0_add_2_12 (.CI(n30557), .I0(displacement_23__N_229[10]), 
            .I1(n15_adj_4420), .CO(n30558));
    SB_CARRY rem_4_add_1318_12 (.CI(n31337), .I0(n1949), .I1(VCC_net), 
            .CO(n31338));
    SB_LUT4 displacement_23__I_0_add_2_11_lut (.I0(GND_net), .I1(displacement_23__N_229[9]), 
            .I2(n16_adj_4421), .I3(n30556), .O(displacement_23__N_80[9])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_15 (.CI(n31082), .I0(n2546_adj_4516), .I1(VCC_net), 
            .CO(n31083));
    SB_LUT4 div_36_i1718_3_lut_3_lut (.I0(n2558), .I1(n7132), .I2(n2553), 
            .I3(GND_net), .O(n2637));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1718_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1318_11_lut (.I0(GND_net), .I1(n1950), .I2(VCC_net), 
            .I3(n31336), .O(n2017)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_14_lut (.I0(GND_net), .I1(n2547_adj_4515), .I2(VCC_net), 
            .I3(n31081), .O(n2614)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_14 (.CI(n31081), .I0(n2547_adj_4515), .I1(VCC_net), 
            .CO(n31082));
    SB_LUT4 i13978_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19010));   // verilog/coms.v(126[12] 289[6])
    defparam i13978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1720_13_lut (.I0(GND_net), .I1(n2548_adj_4514), .I2(VCC_net), 
            .I3(n31080), .O(n2615)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_13 (.CI(n31080), .I0(n2548_adj_4514), .I1(VCC_net), 
            .CO(n31081));
    SB_CARRY rem_4_add_1318_11 (.CI(n31336), .I0(n1950), .I1(VCC_net), 
            .CO(n31337));
    SB_LUT4 rem_4_add_1720_12_lut (.I0(GND_net), .I1(n2549_adj_4513), .I2(VCC_net), 
            .I3(n31079), .O(n2616)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1318_10_lut (.I0(GND_net), .I1(n1951), .I2(VCC_net), 
            .I3(n31335), .O(n2018)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_10 (.CI(n31335), .I0(n1951), .I1(VCC_net), 
            .CO(n31336));
    SB_LUT4 rem_4_add_1318_9_lut (.I0(GND_net), .I1(n1952), .I2(VCC_net), 
            .I3(n31334), .O(n2019)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13979_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n19011));   // verilog/coms.v(126[12] 289[6])
    defparam i13979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13980_3_lut (.I0(\data_out_frame[0] [3]), .I1(n6119), .I2(n18435), 
            .I3(GND_net), .O(n19012));   // verilog/coms.v(126[12] 289[6])
    defparam i13980_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1720_12 (.CI(n31079), .I0(n2549_adj_4513), .I1(VCC_net), 
            .CO(n31080));
    SB_CARRY rem_4_add_1318_9 (.CI(n31334), .I0(n1952), .I1(VCC_net), 
            .CO(n31335));
    SB_LUT4 rem_4_add_1720_11_lut (.I0(GND_net), .I1(n2550_adj_4512), .I2(VCC_net), 
            .I3(n31078), .O(n2617)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_11 (.CI(n30556), .I0(displacement_23__N_229[9]), 
            .I1(n16_adj_4421), .CO(n30557));
    SB_LUT4 rem_4_add_1318_8_lut (.I0(GND_net), .I1(n1953), .I2(VCC_net), 
            .I3(n31333), .O(n2020)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_8 (.CI(n31333), .I0(n1953), .I1(VCC_net), 
            .CO(n31334));
    SB_LUT4 div_36_i1712_3_lut_3_lut (.I0(n2558), .I1(n7126), .I2(n2547), 
            .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1712_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4568));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_1318_7_lut (.I0(GND_net), .I1(n1954), .I2(GND_net), 
            .I3(n31332), .O(n2021)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_11 (.CI(n31078), .I0(n2550_adj_4512), .I1(VCC_net), 
            .CO(n31079));
    SB_LUT4 rem_4_add_1720_10_lut (.I0(GND_net), .I1(n2551_adj_4511), .I2(VCC_net), 
            .I3(n31077), .O(n2618_adj_4507)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_7 (.CI(n31332), .I0(n1954), .I1(GND_net), 
            .CO(n31333));
    SB_LUT4 i13981_3_lut (.I0(\data_out_frame[0] [4]), .I1(n6119), .I2(n18435), 
            .I3(GND_net), .O(n19013));   // verilog/coms.v(126[12] 289[6])
    defparam i13981_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1720_10 (.CI(n31077), .I0(n2551_adj_4511), .I1(VCC_net), 
            .CO(n31078));
    SB_LUT4 rem_4_add_1318_6_lut (.I0(GND_net), .I1(n1955), .I2(GND_net), 
            .I3(n31331), .O(n2022)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_6 (.CI(n31331), .I0(n1955), .I1(GND_net), 
            .CO(n31332));
    SB_LUT4 displacement_23__I_0_add_2_10_lut (.I0(GND_net), .I1(displacement_23__N_229[8]), 
            .I2(n17_adj_4422), .I3(n30555), .O(displacement_23__N_80[8])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_10 (.CI(n30555), .I0(displacement_23__N_229[8]), 
            .I1(n17_adj_4422), .CO(n30556));
    SB_LUT4 rem_4_add_1720_9_lut (.I0(GND_net), .I1(n2552_adj_4510), .I2(VCC_net), 
            .I3(n31076), .O(n2619_adj_4506)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_1665_i41_2_lut (.I0(n2537), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4829));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_i1714_3_lut_3_lut (.I0(n2558), .I1(n7128), .I2(n2549), 
            .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1714_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1720_9 (.CI(n31076), .I0(n2552_adj_4510), .I1(VCC_net), 
            .CO(n31077));
    SB_LUT4 div_36_mux_3_i4_3_lut (.I0(encoder0_position[3]), .I1(n22), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n388));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1318_5_lut (.I0(GND_net), .I1(n1956), .I2(VCC_net), 
            .I3(n31330), .O(n2023)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_5 (.CI(n31330), .I0(n1956), .I1(VCC_net), 
            .CO(n31331));
    SB_LUT4 rem_4_add_1720_8_lut (.I0(GND_net), .I1(n2553_adj_4509), .I2(VCC_net), 
            .I3(n31075), .O(n2620_adj_4502)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13982_3_lut (.I0(\data_out_frame[4] [0]), .I1(ID0), .I2(n14536), 
            .I3(GND_net), .O(n19014));   // verilog/coms.v(126[12] 289[6])
    defparam i13982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1318_4_lut (.I0(GND_net), .I1(n1957), .I2(VCC_net), 
            .I3(n31329), .O(n2024)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_4 (.CI(n31329), .I0(n1957), .I1(VCC_net), 
            .CO(n31330));
    SB_CARRY rem_4_add_1720_8 (.CI(n31075), .I0(n2553_adj_4509), .I1(VCC_net), 
            .CO(n31076));
    SB_LUT4 rem_4_add_1720_7_lut (.I0(GND_net), .I1(n2554), .I2(GND_net), 
            .I3(n31074), .O(n2621_adj_4504)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_7 (.CI(n31074), .I0(n2554), .I1(GND_net), 
            .CO(n31075));
    SB_LUT4 rem_4_add_1318_3_lut (.I0(GND_net), .I1(n1958), .I2(GND_net), 
            .I3(n31328), .O(n2025)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_6_lut (.I0(GND_net), .I1(n2555), .I2(GND_net), 
            .I3(n31073), .O(n2622_adj_4505)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_9_lut (.I0(GND_net), .I1(displacement_23__N_229[7]), 
            .I2(n18_adj_4423), .I3(n30554), .O(displacement_23__N_80[7])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_6 (.CI(n31073), .I0(n2555), .I1(GND_net), 
            .CO(n31074));
    SB_LUT4 div_36_LessThan_1665_i29_2_lut (.I0(n2543), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4822));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1665_i31_2_lut (.I0(n2542), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4823));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1720_5_lut (.I0(GND_net), .I1(n2556), .I2(VCC_net), 
            .I3(n31072), .O(n2623_adj_4503)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_9 (.CI(n30554), .I0(displacement_23__N_229[7]), 
            .I1(n18_adj_4423), .CO(n30555));
    SB_CARRY rem_4_add_1318_3 (.CI(n31328), .I0(n1958), .I1(GND_net), 
            .CO(n31329));
    SB_CARRY rem_4_add_1318_2 (.CI(VCC_net), .I0(n2058), .I1(VCC_net), 
            .CO(n31328));
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_80[22]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_LUT4 rem_4_add_1385_19_lut (.I0(n2075_adj_4609), .I1(n2042), .I2(VCC_net), 
            .I3(n31327), .O(n2141)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i22_3_lut (.I0(bit_ctr[20]), .I1(n42941), .I2(n4754), .I3(GND_net), 
            .O(n35923));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY rem_4_add_1720_5 (.CI(n31072), .I0(n2556), .I1(VCC_net), 
            .CO(n31073));
    SB_LUT4 rem_4_add_1720_4_lut (.I0(GND_net), .I1(n2557), .I2(VCC_net), 
            .I3(n31071), .O(n2624_adj_4501)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_18_lut (.I0(GND_net), .I1(n2043), .I2(VCC_net), 
            .I3(n31326), .O(n2110)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_1665_i23_2_lut (.I0(n2546), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4819));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i23_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1720_4 (.CI(n31071), .I0(n2557), .I1(VCC_net), 
            .CO(n31072));
    SB_LUT4 div_36_LessThan_1665_i25_2_lut (.I0(n2545), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4820));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1720_3_lut (.I0(GND_net), .I1(n2558_adj_4508), .I2(GND_net), 
            .I3(n31070), .O(n2625_adj_4500)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_3 (.CI(n31070), .I0(n2558_adj_4508), .I1(GND_net), 
            .CO(n31071));
    SB_CARRY rem_4_add_1385_18 (.CI(n31326), .I0(n2043), .I1(VCC_net), 
            .CO(n31327));
    SB_LUT4 div_36_LessThan_1665_i27_2_lut (.I0(n2544), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4821));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i27_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1720_2 (.CI(VCC_net), .I0(n2658), .I1(VCC_net), 
            .CO(n31070));
    SB_LUT4 rem_4_add_1787_25_lut (.I0(n2669), .I1(n2636_adj_4495), .I2(VCC_net), 
            .I3(n31069), .O(n2735)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1787_24_lut (.I0(GND_net), .I1(n2637_adj_4492), .I2(VCC_net), 
            .I3(n31068), .O(n2704_adj_4480)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_24 (.CI(n31068), .I0(n2637_adj_4492), .I1(VCC_net), 
            .CO(n31069));
    SB_LUT4 displacement_23__I_0_add_2_8_lut (.I0(GND_net), .I1(displacement_23__N_229[6]), 
            .I2(n19_adj_4424), .I3(n30553), .O(displacement_23__N_80[6])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_23_lut (.I0(GND_net), .I1(n2638_adj_4491), .I2(VCC_net), 
            .I3(n31067), .O(n2705_adj_4479)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_23 (.CI(n31067), .I0(n2638_adj_4491), .I1(VCC_net), 
            .CO(n31068));
    SB_LUT4 rem_4_add_1787_22_lut (.I0(GND_net), .I1(n2639), .I2(VCC_net), 
            .I3(n31066), .O(n2706_adj_4478)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_22 (.CI(n31066), .I0(n2639), .I1(VCC_net), 
            .CO(n31067));
    SB_LUT4 rem_4_add_1385_17_lut (.I0(GND_net), .I1(n2044), .I2(VCC_net), 
            .I3(n31325), .O(n2111)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_17 (.CI(n31325), .I0(n2044), .I1(VCC_net), 
            .CO(n31326));
    SB_LUT4 div_36_LessThan_1665_i13_2_lut (.I0(n2551), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4810));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1787_21_lut (.I0(GND_net), .I1(n2640), .I2(VCC_net), 
            .I3(n31065), .O(n2707_adj_4477)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_21_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_80[21]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_80[20]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_80[19]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_80[18]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_80[17]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_CARRY rem_4_add_1787_21 (.CI(n31065), .I0(n2640), .I1(VCC_net), 
            .CO(n31066));
    SB_LUT4 div_36_LessThan_1665_i15_2_lut (.I0(n2550), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4812));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1385_16_lut (.I0(GND_net), .I1(n2045), .I2(VCC_net), 
            .I3(n31324), .O(n2112)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_20_lut (.I0(GND_net), .I1(n2641), .I2(VCC_net), 
            .I3(n31064), .O(n2708_adj_4476)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13985_3_lut (.I0(\data_out_frame[4] [2]), .I1(ID2), .I2(n14536), 
            .I3(GND_net), .O(n19017));   // verilog/coms.v(126[12] 289[6])
    defparam i13985_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_80[16]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_80[15]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_80[14]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_80[13]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_80[12]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_80[11]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_80[10]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_80[9]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_80[8]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_80[7]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_80[6]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_80[5]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_80[4]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_80[3]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_80[2]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_80[1]));   // verilog/TinyFPGA_B.v(242[10] 244[6])
    SB_CARRY rem_4_add_1787_20 (.CI(n31064), .I0(n2641), .I1(VCC_net), 
            .CO(n31065));
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[22]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[21]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[20]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[19]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[18]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[17]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[16]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[15]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[14]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[13]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[12]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[11]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[10]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[9]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[8]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[7]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[6]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_LUT4 rem_4_add_1787_19_lut (.I0(GND_net), .I1(n2642_adj_4490), .I2(VCC_net), 
            .I3(n31063), .O(n2709_adj_4475)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_1665_i17_2_lut (.I0(n2549), .I1(n95_adj_4360), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4814));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i17_2_lut.LUT_INIT = 16'h9999;
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[5]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[4]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[3]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[2]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[1]));   // verilog/TinyFPGA_B.v(127[10] 140[6])
    SB_DFF communication_counter_1146__i0 (.Q(communication_counter[0]), .C(LED_c), 
           .D(n165));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_CARRY rem_4_add_1385_16 (.CI(n31324), .I0(n2045), .I1(VCC_net), 
            .CO(n31325));
    SB_LUT4 div_36_LessThan_1665_i19_2_lut (.I0(n2548), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4816));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i19_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY displacement_23__I_0_add_2_8 (.CI(n30553), .I0(displacement_23__N_229[6]), 
            .I1(n19_adj_4424), .CO(n30554));
    SB_LUT4 i13986_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n14536), .I3(GND_net), .O(n19018));   // verilog/coms.v(126[12] 289[6])
    defparam i13986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1665_i21_2_lut (.I0(n2547), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4817));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1665_i33_2_lut (.I0(n2541), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4824));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1385_15_lut (.I0(GND_net), .I1(n2046), .I2(VCC_net), 
            .I3(n31323), .O(n2113)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_15 (.CI(n31323), .I0(n2046), .I1(VCC_net), 
            .CO(n31324));
    SB_CARRY rem_4_add_1787_19 (.CI(n31063), .I0(n2642_adj_4490), .I1(VCC_net), 
            .CO(n31064));
    SB_LUT4 i14070_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n14536), 
            .I3(GND_net), .O(n19102));   // verilog/coms.v(126[12] 289[6])
    defparam i14070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_add_2_7_lut (.I0(GND_net), .I1(displacement_23__N_229[5]), 
            .I2(n20_adj_4425), .I3(n30552), .O(displacement_23__N_80[5])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_18_lut (.I0(GND_net), .I1(n2643_adj_4489), .I2(VCC_net), 
            .I3(n31062), .O(n2710_adj_4474)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_14_lut (.I0(GND_net), .I1(n2047), .I2(VCC_net), 
            .I3(n31322), .O(n2114)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_14 (.CI(n31322), .I0(n2047), .I1(VCC_net), 
            .CO(n31323));
    SB_LUT4 div_36_LessThan_1665_i35_2_lut (.I0(n2540), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4825));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1385_13_lut (.I0(GND_net), .I1(n2048), .I2(VCC_net), 
            .I3(n31321), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14071_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n14536), 
            .I3(GND_net), .O(n19103));   // verilog/coms.v(126[12] 289[6])
    defparam i14071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14395_3_lut (.I0(setpoint[1]), .I1(n4660), .I2(n39863), .I3(GND_net), 
            .O(n19427));   // verilog/coms.v(126[12] 289[6])
    defparam i14395_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_LessThan_1665_i37_2_lut (.I0(n2539), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4827));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i37_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1385_13 (.CI(n31321), .I0(n2048), .I1(VCC_net), 
            .CO(n31322));
    SB_LUT4 div_36_LessThan_1665_i39_2_lut (.I0(n2538), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4828));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i39_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1787_18 (.CI(n31062), .I0(n2643_adj_4489), .I1(VCC_net), 
            .CO(n31063));
    SB_LUT4 rem_4_add_1385_12_lut (.I0(GND_net), .I1(n2049), .I2(VCC_net), 
            .I3(n31320), .O(n2116)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i1667_1_lut (.I0(n2558), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2559));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1667_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY displacement_23__I_0_add_2_7 (.CI(n30552), .I0(displacement_23__N_229[5]), 
            .I1(n20_adj_4425), .CO(n30553));
    SB_CARRY rem_4_add_1385_12 (.CI(n31320), .I0(n2049), .I1(VCC_net), 
            .CO(n31321));
    SB_LUT4 rem_4_add_1385_11_lut (.I0(GND_net), .I1(n2050), .I2(VCC_net), 
            .I3(n31319), .O(n2117)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_17_lut (.I0(GND_net), .I1(n2644), .I2(VCC_net), 
            .I3(n31061), .O(n2711_adj_4473)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_17 (.CI(n31061), .I0(n2644), .I1(VCC_net), 
            .CO(n31062));
    SB_LUT4 i36060_4_lut (.I0(n33_adj_4824), .I1(n21_adj_4817), .I2(n19_adj_4816), 
            .I3(n17_adj_4814), .O(n43184));
    defparam i36060_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY rem_4_add_1385_11 (.CI(n31319), .I0(n2050), .I1(VCC_net), 
            .CO(n31320));
    SB_LUT4 displacement_23__I_0_add_2_6_lut (.I0(GND_net), .I1(displacement_23__N_229[4]), 
            .I2(n21_adj_4426), .I3(n30551), .O(displacement_23__N_80[4])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36800_4_lut (.I0(n15_adj_4812), .I1(n13_adj_4810), .I2(n2552), 
            .I3(n98), .O(n43925));
    defparam i36800_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i37246_4_lut (.I0(n21_adj_4817), .I1(n19_adj_4816), .I2(n17_adj_4814), 
            .I3(n43925), .O(n44371));
    defparam i37246_4_lut.LUT_INIT = 16'hfeff;
    SB_CARRY displacement_23__I_0_add_2_6 (.CI(n30551), .I0(displacement_23__N_229[4]), 
            .I1(n21_adj_4426), .CO(n30552));
    SB_LUT4 rem_4_add_1385_10_lut (.I0(GND_net), .I1(n2051), .I2(VCC_net), 
            .I3(n31318), .O(n2118)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37244_4_lut (.I0(n27_adj_4821), .I1(n25_adj_4820), .I2(n23_adj_4819), 
            .I3(n44371), .O(n44369));
    defparam i37244_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i36062_4_lut (.I0(n33_adj_4824), .I1(n31_adj_4823), .I2(n29_adj_4822), 
            .I3(n44369), .O(n43186));
    defparam i36062_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_36_LessThan_1665_i10_4_lut (.I0(n388), .I1(n99), .I2(n2553), 
            .I3(n558), .O(n10_adj_4808));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i10_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i37699_3_lut (.I0(n10_adj_4808), .I1(n87), .I2(n33_adj_4824), 
            .I3(GND_net), .O(n44824));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37699_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37700_3_lut (.I0(n44824), .I1(n86), .I2(n35_adj_4825), .I3(GND_net), 
            .O(n44825));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37700_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_36_LessThan_1665_i36_3_lut (.I0(n18_adj_4815), .I1(n83), 
            .I2(n41_adj_4829), .I3(GND_net), .O(n36_adj_4826));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36052_4_lut (.I0(n39_adj_4828), .I1(n37_adj_4827), .I2(n35_adj_4825), 
            .I3(n43184), .O(n43176));
    defparam i36052_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37914_4_lut (.I0(n36_adj_4826), .I1(n16_adj_4813), .I2(n41_adj_4829), 
            .I3(n43172), .O(n45039));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37914_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i37560_3_lut (.I0(n44825), .I1(n85), .I2(n37_adj_4827), .I3(GND_net), 
            .O(n44685));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37560_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_36_LessThan_1665_i22_3_lut (.I0(n14_adj_4811), .I1(n91), 
            .I2(n25_adj_4820), .I3(GND_net), .O(n22_adj_4818));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i22_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37912_4_lut (.I0(n22_adj_4818), .I1(n12_adj_4809), .I2(n25_adj_4820), 
            .I3(n43205), .O(n45037));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37912_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i14072_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n14536), 
            .I3(GND_net), .O(n19104));   // verilog/coms.v(126[12] 289[6])
    defparam i14072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14073_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n14536), 
            .I3(GND_net), .O(n19105));   // verilog/coms.v(126[12] 289[6])
    defparam i14073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14074_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n14536), 
            .I3(GND_net), .O(n19106));   // verilog/coms.v(126[12] 289[6])
    defparam i14074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14075_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n14536), 
            .I3(GND_net), .O(n19107));   // verilog/coms.v(126[12] 289[6])
    defparam i14075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1801_3_lut (.I0(n2648), .I1(n2715_adj_4469), .I2(n2669), 
            .I3(GND_net), .O(n2747));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37913_3_lut (.I0(n45037), .I1(n90), .I2(n27_adj_4821), .I3(GND_net), 
            .O(n45038));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37913_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37830_3_lut (.I0(n45038), .I1(n89), .I2(n29_adj_4822), .I3(GND_net), 
            .O(n44955));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37830_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37472_4_lut (.I0(n39_adj_4828), .I1(n37_adj_4827), .I2(n35_adj_4825), 
            .I3(n43186), .O(n44597));
    defparam i37472_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i37985_4_lut (.I0(n44685), .I1(n45039), .I2(n41_adj_4829), 
            .I3(n43176), .O(n45110));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37985_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i37754_3_lut (.I0(n44955), .I1(n88), .I2(n31_adj_4823), .I3(GND_net), 
            .O(n44879));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37754_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i38001_4_lut (.I0(n44879), .I1(n45110), .I2(n41_adj_4829), 
            .I3(n44597), .O(n45126));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i38001_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i38002_3_lut (.I0(n45126), .I1(n82), .I2(n2536), .I3(GND_net), 
            .O(n45127));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i38002_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i37998_3_lut (.I0(n45127), .I1(n81), .I2(n2535), .I3(GND_net), 
            .O(n45123));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37998_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 rem_4_i1800_3_lut (.I0(n2647), .I1(n2714_adj_4470), .I2(n2669), 
            .I3(GND_net), .O(n2746));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1800_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1620 (.I0(n45123), .I1(n17241), .I2(n80), .I3(n2534), 
            .O(n2558));
    defparam i1_4_lut_adj_1620.LUT_INIT = 16'hceef;
    SB_CARRY rem_4_add_1385_10 (.CI(n31318), .I0(n2051), .I1(VCC_net), 
            .CO(n31319));
    SB_LUT4 rem_4_add_1385_9_lut (.I0(GND_net), .I1(n2052), .I2(VCC_net), 
            .I3(n31317), .O(n2119)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_9 (.CI(n31317), .I0(n2052), .I1(VCC_net), 
            .CO(n31318));
    SB_LUT4 displacement_23__I_0_add_2_5_lut (.I0(GND_net), .I1(displacement_23__N_229[3]), 
            .I2(n22_adj_4427), .I3(n30550), .O(displacement_23__N_80[3])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_8_lut (.I0(GND_net), .I1(n2053), .I2(VCC_net), 
            .I3(n31316), .O(n2120)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_5 (.CI(n30550), .I0(displacement_23__N_229[3]), 
            .I1(n22_adj_4427), .CO(n30551));
    SB_CARRY rem_4_add_1385_8 (.CI(n31316), .I0(n2053), .I1(VCC_net), 
            .CO(n31317));
    SB_LUT4 displacement_23__I_0_add_2_4_lut (.I0(GND_net), .I1(displacement_23__N_229[2]), 
            .I2(n23_adj_4428), .I3(n30549), .O(displacement_23__N_80[2])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1803_3_lut (.I0(n2650), .I1(n2717_adj_4467), .I2(n2669), 
            .I3(GND_net), .O(n2749));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14076_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n14536), 
            .I3(GND_net), .O(n19108));   // verilog/coms.v(126[12] 289[6])
    defparam i14076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1385_7_lut (.I0(GND_net), .I1(n2054), .I2(GND_net), 
            .I3(n31315), .O(n2121)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_7 (.CI(n31315), .I0(n2054), .I1(GND_net), 
            .CO(n31316));
    SB_LUT4 rem_4_add_1787_16_lut (.I0(GND_net), .I1(n2645), .I2(VCC_net), 
            .I3(n31060), .O(n2712_adj_4472)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_4 (.CI(n30549), .I0(displacement_23__N_229[2]), 
            .I1(n23_adj_4428), .CO(n30550));
    SB_LUT4 rem_4_i1807_3_lut (.I0(n2654), .I1(n2721), .I2(n2669), .I3(GND_net), 
            .O(n2753));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1805_3_lut (.I0(n2652), .I1(n2719_adj_4465), .I2(n2669), 
            .I3(GND_net), .O(n2751));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1804_3_lut (.I0(n2651), .I1(n2718_adj_4466), .I2(n2669), 
            .I3(GND_net), .O(n2750));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1797_3_lut (.I0(n2644), .I1(n2711_adj_4473), .I2(n2669), 
            .I3(GND_net), .O(n2743));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1385_6_lut (.I0(GND_net), .I1(n2055), .I2(GND_net), 
            .I3(n31314), .O(n2122)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14077_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n14536), 
            .I3(GND_net), .O(n19109));   // verilog/coms.v(126[12] 289[6])
    defparam i14077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1593_3_lut (.I0(n2344), .I1(n2411), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2443));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1795_3_lut (.I0(n2642_adj_4490), .I1(n2709_adj_4475), 
            .I2(n2669), .I3(GND_net), .O(n2741));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1799_3_lut (.I0(n2646), .I1(n2713_adj_4471), .I2(n2669), 
            .I3(GND_net), .O(n2745));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1799_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1385_6 (.CI(n31314), .I0(n2055), .I1(GND_net), 
            .CO(n31315));
    SB_LUT4 rem_4_add_1385_5_lut (.I0(GND_net), .I1(n2056), .I2(VCC_net), 
            .I3(n31313), .O(n2123)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_16 (.CI(n31060), .I0(n2645), .I1(VCC_net), 
            .CO(n31061));
    SB_LUT4 rem_4_i1591_3_lut (.I0(n2342), .I1(n2409), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2441));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1592_3_lut (.I0(n2343), .I1(n2410), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2442));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1385_5 (.CI(n31313), .I0(n2056), .I1(VCC_net), 
            .CO(n31314));
    SB_LUT4 rem_4_add_1787_15_lut (.I0(GND_net), .I1(n2646), .I2(VCC_net), 
            .I3(n31059), .O(n2713_adj_4471)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_4_lut (.I0(GND_net), .I1(n2057), .I2(VCC_net), 
            .I3(n31312), .O(n2124)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1590_3_lut (.I0(n2341), .I1(n2408), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2440));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1385_4 (.CI(n31312), .I0(n2057), .I1(VCC_net), 
            .CO(n31313));
    SB_LUT4 i37250_3_lut (.I0(n2252), .I1(n2319), .I2(n2273_adj_4591), 
            .I3(GND_net), .O(n2351));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i37250_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1787_15 (.CI(n31059), .I0(n2646), .I1(VCC_net), 
            .CO(n31060));
    SB_LUT4 i14408_3_lut (.I0(setpoint[14]), .I1(n4673), .I2(n39863), 
            .I3(GND_net), .O(n19440));   // verilog/coms.v(126[12] 289[6])
    defparam i14408_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14407_3_lut (.I0(setpoint[13]), .I1(n4672), .I2(n39863), 
            .I3(GND_net), .O(n19439));   // verilog/coms.v(126[12] 289[6])
    defparam i14407_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14406_3_lut (.I0(setpoint[12]), .I1(n4671), .I2(n39863), 
            .I3(GND_net), .O(n19438));   // verilog/coms.v(126[12] 289[6])
    defparam i14406_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14405_3_lut (.I0(setpoint[11]), .I1(n4670), .I2(n39863), 
            .I3(GND_net), .O(n19437));   // verilog/coms.v(126[12] 289[6])
    defparam i14405_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14404_3_lut (.I0(setpoint[10]), .I1(n4669), .I2(n39863), 
            .I3(GND_net), .O(n19436));   // verilog/coms.v(126[12] 289[6])
    defparam i14404_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14403_3_lut (.I0(setpoint[9]), .I1(n4668), .I2(n39863), .I3(GND_net), 
            .O(n19435));   // verilog/coms.v(126[12] 289[6])
    defparam i14403_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1787_14_lut (.I0(GND_net), .I1(n2647), .I2(VCC_net), 
            .I3(n31058), .O(n2714_adj_4470)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_3_lut (.I0(GND_net), .I1(n2058), .I2(GND_net), 
            .I3(n31311), .O(n2125)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_14 (.CI(n31058), .I0(n2647), .I1(VCC_net), 
            .CO(n31059));
    SB_LUT4 rem_4_add_1787_13_lut (.I0(GND_net), .I1(n2648), .I2(VCC_net), 
            .I3(n31057), .O(n2715_adj_4469)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_3 (.CI(n31311), .I0(n2058), .I1(GND_net), 
            .CO(n31312));
    SB_CARRY rem_4_add_1787_13 (.CI(n31057), .I0(n2648), .I1(VCC_net), 
            .CO(n31058));
    SB_LUT4 rem_4_add_1787_12_lut (.I0(GND_net), .I1(n2649), .I2(VCC_net), 
            .I3(n31056), .O(n2716_adj_4468)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_3_lut (.I0(GND_net), .I1(displacement_23__N_229[1]), 
            .I2(n24_adj_4429), .I3(n30548), .O(displacement_23__N_80[1])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_12 (.CI(n31056), .I0(n2649), .I1(VCC_net), 
            .CO(n31057));
    SB_LUT4 rem_4_add_1787_11_lut (.I0(GND_net), .I1(n2650), .I2(VCC_net), 
            .I3(n31055), .O(n2717_adj_4467)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_2 (.CI(VCC_net), .I0(n2158), .I1(VCC_net), 
            .CO(n31311));
    SB_LUT4 rem_4_add_1452_20_lut (.I0(n2174_adj_4597), .I1(n2141), .I2(VCC_net), 
            .I3(n31310), .O(n2240)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY displacement_23__I_0_add_2_3 (.CI(n30548), .I0(displacement_23__N_229[1]), 
            .I1(n24_adj_4429), .CO(n30549));
    SB_LUT4 rem_4_add_1452_19_lut (.I0(GND_net), .I1(n2142), .I2(VCC_net), 
            .I3(n31309), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_19 (.CI(n31309), .I0(n2142), .I1(VCC_net), 
            .CO(n31310));
    SB_LUT4 rem_4_add_1452_18_lut (.I0(GND_net), .I1(n2143), .I2(VCC_net), 
            .I3(n31308), .O(n2210)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_2_lut (.I0(GND_net), .I1(displacement_23__N_229[0]), 
            .I2(n25_adj_4430), .I3(VCC_net), .O(displacement_23__N_80[0])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_11 (.CI(n31055), .I0(n2650), .I1(VCC_net), 
            .CO(n31056));
    SB_LUT4 rem_4_add_1787_10_lut (.I0(GND_net), .I1(n2651), .I2(VCC_net), 
            .I3(n31054), .O(n2718_adj_4466)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_18 (.CI(n31308), .I0(n2143), .I1(VCC_net), 
            .CO(n31309));
    SB_CARRY rem_4_add_1787_10 (.CI(n31054), .I0(n2651), .I1(VCC_net), 
            .CO(n31055));
    SB_LUT4 rem_4_add_1787_9_lut (.I0(GND_net), .I1(n2652), .I2(VCC_net), 
            .I3(n31053), .O(n2719_adj_4465)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36505_3_lut_3_lut (.I0(n392), .I1(n558), .I2(n369), .I3(GND_net), 
            .O(n510));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36505_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 i37251_3_lut (.I0(n2351), .I1(n2418), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2450_adj_4583));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i37251_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1787_9 (.CI(n31053), .I0(n2652), .I1(VCC_net), 
            .CO(n31054));
    SB_IO PIN_19_pad (.PACKAGE_PIN(PIN_19), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_19_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_19_pad.PIN_TYPE = 6'b011001;
    defparam PIN_19_pad.PULLUP = 1'b0;
    defparam PIN_19_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 rem_4_i1602_3_lut (.I0(n2353), .I1(n2420), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2452_adj_4581));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1056_3_lut (.I0(n1551), .I1(n1618), .I2(n1580), .I3(GND_net), 
            .O(n1650_adj_4485));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1055_3_lut (.I0(n1550), .I1(n1617), .I2(n1580), .I3(GND_net), 
            .O(n1649_adj_4484));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1061_3_lut (.I0(n1556), .I1(n1623), .I2(n1580), .I3(GND_net), 
            .O(n1655));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1060_3_lut (.I0(n1555), .I1(n1622), .I2(n1580), .I3(GND_net), 
            .O(n1654));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1054_3_lut (.I0(n1549), .I1(n1616), .I2(n1580), .I3(GND_net), 
            .O(n1648_adj_4483));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1057_3_lut (.I0(n1552), .I1(n1619), .I2(n1580), .I3(GND_net), 
            .O(n1651_adj_4486));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1059_rep_40_3_lut (.I0(n1554_adj_4494), .I1(n1621), .I2(n1580), 
            .I3(GND_net), .O(n1653_adj_4488));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1059_rep_40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i988_3_lut (.I0(n1451), .I1(n1518), .I2(n1481), .I3(GND_net), 
            .O(n1550));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i987_3_lut (.I0(n1450), .I1(n1517), .I2(n1481), .I3(GND_net), 
            .O(n1549));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i986_3_lut (.I0(n1449), .I1(n1516), .I2(n1481), .I3(GND_net), 
            .O(n1548));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1621 (.I0(n1556), .I1(n1557), .I2(n1558), .I3(GND_net), 
            .O(n38270));
    defparam i1_3_lut_adj_1621.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut (.I0(n1554_adj_4494), .I1(n1551), .I2(n38270), .I3(n1555), 
            .O(n11_adj_4445));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i3_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i5_4_lut (.I0(n1548), .I1(n1549), .I2(n1547), .I3(n1550), 
            .O(n13_adj_4444));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(n13_adj_4444), .I1(n11_adj_4445), .I2(n1553_adj_4493), 
            .I3(n1552), .O(n1580));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1063_3_lut (.I0(n1558), .I1(n1625), .I2(n1580), .I3(GND_net), 
            .O(n1657));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1062_3_lut (.I0(n1557), .I1(n1624), .I2(n1580), .I3(GND_net), 
            .O(n1656));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1787_8_lut (.I0(GND_net), .I1(n2653), .I2(VCC_net), 
            .I3(n31052), .O(n2720_adj_4464)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_8 (.CI(n31052), .I0(n2653), .I1(VCC_net), 
            .CO(n31053));
    SB_LUT4 rem_4_add_1787_7_lut (.I0(GND_net), .I1(n2654), .I2(GND_net), 
            .I3(n31051), .O(n2721)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_7 (.CI(n31051), .I0(n2654), .I1(GND_net), 
            .CO(n31052));
    SB_LUT4 div_36_i274_4_lut_4_lut (.I0(n392), .I1(n99), .I2(n2), .I3(n5_adj_4915), 
            .O(n38022));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i274_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 rem_4_add_1787_6_lut (.I0(GND_net), .I1(n2655), .I2(GND_net), 
            .I3(n31050), .O(n2722)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_6 (.CI(n31050), .I0(n2655), .I1(GND_net), 
            .CO(n31051));
    SB_LUT4 rem_4_add_1787_5_lut (.I0(GND_net), .I1(n2656), .I2(VCC_net), 
            .I3(n31049), .O(n2723_adj_4463)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_5 (.CI(n31049), .I0(n2656), .I1(VCC_net), 
            .CO(n31050));
    SB_LUT4 rem_4_add_1787_4_lut (.I0(GND_net), .I1(n2657), .I2(VCC_net), 
            .I3(n31048), .O(n2724_adj_4462)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1597_3_lut (.I0(n2348), .I1(n2415), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2447_adj_4586));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1597_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1787_4 (.CI(n31048), .I0(n2657), .I1(VCC_net), 
            .CO(n31049));
    SB_LUT4 rem_4_add_1452_17_lut (.I0(GND_net), .I1(n2144), .I2(VCC_net), 
            .I3(n31307), .O(n2211)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1603_3_lut (.I0(n2354), .I1(n2421), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2453_adj_4580));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1596_3_lut (.I0(n2347), .I1(n2414), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2446));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1596_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY displacement_23__I_0_add_2_2 (.CI(VCC_net), .I0(displacement_23__N_229[0]), 
            .I1(n25_adj_4430), .CO(n30548));
    SB_LUT4 rem_4_add_1787_3_lut (.I0(GND_net), .I1(n2658), .I2(GND_net), 
            .I3(n31047), .O(n2725)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_3 (.CI(n31047), .I0(n2658), .I1(GND_net), 
            .CO(n31048));
    SB_LUT4 rem_4_i1798_3_lut (.I0(n2645), .I1(n2712_adj_4472), .I2(n2669), 
            .I3(GND_net), .O(n2744));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1802_3_lut (.I0(n2649), .I1(n2716_adj_4468), .I2(n2669), 
            .I3(GND_net), .O(n2748));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1802_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1787_2 (.CI(VCC_net), .I0(n2758), .I1(VCC_net), 
            .CO(n31047));
    SB_LUT4 rem_4_add_1854_26_lut (.I0(n2768), .I1(n2735), .I2(VCC_net), 
            .I3(n31046), .O(n2834_adj_4451)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_1452_17 (.CI(n31307), .I0(n2144), .I1(VCC_net), 
            .CO(n31308));
    SB_LUT4 rem_4_add_1452_16_lut (.I0(GND_net), .I1(n2145), .I2(VCC_net), 
            .I3(n31306), .O(n2212)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1595_3_lut (.I0(n2346), .I1(n2413), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2445));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1854_25_lut (.I0(GND_net), .I1(n2736), .I2(VCC_net), 
            .I3(n31045), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_25 (.CI(n31045), .I0(n2736), .I1(VCC_net), 
            .CO(n31046));
    SB_LUT4 rem_4_add_1854_24_lut (.I0(GND_net), .I1(n2737), .I2(VCC_net), 
            .I3(n31044), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_24 (.CI(n31044), .I0(n2737), .I1(VCC_net), 
            .CO(n31045));
    SB_LUT4 rem_4_i1594_3_lut (.I0(n2345), .I1(n2412), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2444));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37254_3_lut (.I0(n2250), .I1(n2317), .I2(n2273_adj_4591), 
            .I3(GND_net), .O(n2349));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i37254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1854_23_lut (.I0(GND_net), .I1(n2738), .I2(VCC_net), 
            .I3(n31043), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_23 (.CI(n31043), .I0(n2738), .I1(VCC_net), 
            .CO(n31044));
    SB_LUT4 rem_4_add_1854_22_lut (.I0(GND_net), .I1(n2739), .I2(VCC_net), 
            .I3(n31042), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37255_3_lut (.I0(n2349), .I1(n2416), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2448_adj_4585));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i37255_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1854_22 (.CI(n31042), .I0(n2739), .I1(VCC_net), 
            .CO(n31043));
    SB_LUT4 rem_4_add_1854_21_lut (.I0(GND_net), .I1(n2740), .I2(VCC_net), 
            .I3(n31041), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37248_3_lut (.I0(n2253), .I1(n2320), .I2(n2273_adj_4591), 
            .I3(GND_net), .O(n2352));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i37248_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37249_3_lut (.I0(n2352), .I1(n2419), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2451_adj_4582));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i37249_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37252_3_lut (.I0(n2251), .I1(n2318), .I2(n2273_adj_4591), 
            .I3(GND_net), .O(n2350));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i37252_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1806_3_lut (.I0(n2653), .I1(n2720_adj_4464), .I2(n2669), 
            .I3(GND_net), .O(n2752));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1806_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36502_3_lut_3_lut (.I0(n533), .I1(n558), .I2(n370), .I3(GND_net), 
            .O(n649));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36502_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 i37253_3_lut (.I0(n2350), .I1(n2417), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2449_adj_4584));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i37253_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1854_21 (.CI(n31041), .I0(n2740), .I1(VCC_net), 
            .CO(n31042));
    SB_CARRY rem_4_add_1452_16 (.CI(n31306), .I0(n2145), .I1(VCC_net), 
            .CO(n31307));
    SB_LUT4 rem_4_mux_3_i12_3_lut (.I0(communication_counter[11]), .I1(n22_adj_4390), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2458_adj_4575));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1606_3_lut (.I0(n2357_adj_4589), .I1(n2424), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2456_adj_4577));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1589_3_lut (.I0(n2340), .I1(n2407), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2439));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1053_3_lut (.I0(n1548), .I1(n1615), .I2(n1580), .I3(GND_net), 
            .O(n1647_adj_4482));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i367_4_lut_4_lut (.I0(n533), .I1(n98), .I2(n4_adj_4339), 
            .I3(n38022), .O(n38024));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i367_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 rem_4_i1524_3_lut (.I0(n2243), .I1(n2310), .I2(n2273_adj_4591), 
            .I3(GND_net), .O(n2342));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1523_3_lut (.I0(n2242), .I1(n2309), .I2(n2273_adj_4591), 
            .I3(GND_net), .O(n2341));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i368_4_lut_4_lut (.I0(n533), .I1(n99), .I2(n2_adj_4601), 
            .I3(n510), .O(n648));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i368_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 rem_4_i1796_3_lut (.I0(n2643_adj_4489), .I1(n2710_adj_4474), 
            .I2(n2669), .I3(GND_net), .O(n2742));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1522_3_lut (.I0(n2241), .I1(n2308), .I2(n2273_adj_4591), 
            .I3(GND_net), .O(n2340));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1854_20_lut (.I0(GND_net), .I1(n2741), .I2(VCC_net), 
            .I3(n31040), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1793_3_lut (.I0(n2640), .I1(n2707_adj_4477), .I2(n2669), 
            .I3(GND_net), .O(n2739));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1707_3_lut_3_lut (.I0(n2558), .I1(n7121), .I2(n2542), 
            .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1707_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1529_3_lut (.I0(n2248), .I1(n2315), .I2(n2273_adj_4591), 
            .I3(GND_net), .O(n2347));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1529_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1854_20 (.CI(n31040), .I0(n2741), .I1(VCC_net), 
            .CO(n31041));
    SB_LUT4 rem_4_add_1452_15_lut (.I0(GND_net), .I1(n2146), .I2(VCC_net), 
            .I3(n31305), .O(n2213)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_19_lut (.I0(GND_net), .I1(n2742), .I2(VCC_net), 
            .I3(n31039), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_19 (.CI(n31039), .I0(n2742), .I1(VCC_net), 
            .CO(n31040));
    SB_LUT4 rem_4_add_1854_18_lut (.I0(GND_net), .I1(n2743), .I2(VCC_net), 
            .I3(n31038), .O(n2810)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1528_3_lut (.I0(n2247), .I1(n2314), .I2(n2273_adj_4591), 
            .I3(GND_net), .O(n2346));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1530_3_lut (.I0(n2249), .I1(n2316), .I2(n2273_adj_4591), 
            .I3(GND_net), .O(n2348));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1530_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1854_18 (.CI(n31038), .I0(n2743), .I1(VCC_net), 
            .CO(n31039));
    SB_LUT4 rem_4_i1535_3_lut (.I0(n2254), .I1(n2321), .I2(n2273_adj_4591), 
            .I3(GND_net), .O(n2353));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1854_17_lut (.I0(GND_net), .I1(n2744), .I2(VCC_net), 
            .I3(n31037), .O(n2811)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1526_3_lut (.I0(n2245), .I1(n2312), .I2(n2273_adj_4591), 
            .I3(GND_net), .O(n2344));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1526_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1854_17 (.CI(n31037), .I0(n2744), .I1(VCC_net), 
            .CO(n31038));
    SB_LUT4 rem_4_add_1854_16_lut (.I0(GND_net), .I1(n2745), .I2(VCC_net), 
            .I3(n31036), .O(n2812)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1527_3_lut (.I0(n2246), .I1(n2313), .I2(n2273_adj_4591), 
            .I3(GND_net), .O(n2345));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1527_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1854_16 (.CI(n31036), .I0(n2745), .I1(VCC_net), 
            .CO(n31037));
    SB_LUT4 rem_4_i1792_3_lut (.I0(n2639), .I1(n2706_adj_4478), .I2(n2669), 
            .I3(GND_net), .O(n2738));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1854_15_lut (.I0(GND_net), .I1(n2746), .I2(VCC_net), 
            .I3(n31035), .O(n2813)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_15 (.CI(n31035), .I0(n2746), .I1(VCC_net), 
            .CO(n31036));
    SB_LUT4 rem_4_i1525_3_lut (.I0(n2244), .I1(n2311), .I2(n2273_adj_4591), 
            .I3(GND_net), .O(n2343));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1525_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1538_3_lut (.I0(n2257), .I1(n2324), .I2(n2273_adj_4591), 
            .I3(GND_net), .O(n2356));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1465_rep_32_3_lut (.I0(n2152), .I1(n2219), .I2(n2174_adj_4597), 
            .I3(GND_net), .O(n2251));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1465_rep_32_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1854_14_lut (.I0(GND_net), .I1(n2747), .I2(VCC_net), 
            .I3(n31034), .O(n2814)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_14 (.CI(n31034), .I0(n2747), .I1(VCC_net), 
            .CO(n31035));
    SB_LUT4 rem_4_add_1854_13_lut (.I0(GND_net), .I1(n2748), .I2(VCC_net), 
            .I3(n31033), .O(n2815)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_13 (.CI(n31033), .I0(n2748), .I1(VCC_net), 
            .CO(n31034));
    SB_LUT4 rem_4_i1791_3_lut (.I0(n2638_adj_4491), .I1(n2705_adj_4479), 
            .I2(n2669), .I3(GND_net), .O(n2737));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1464_rep_30_3_lut (.I0(n2151), .I1(n2218), .I2(n2174_adj_4597), 
            .I3(GND_net), .O(n2250));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1464_rep_30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1461_3_lut (.I0(n2148), .I1(n2215), .I2(n2174_adj_4597), 
            .I3(GND_net), .O(n2247));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1461_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1452_15 (.CI(n31305), .I0(n2146), .I1(VCC_net), 
            .CO(n31306));
    SB_LUT4 rem_4_i1790_3_lut (.I0(n2637_adj_4492), .I1(n2704_adj_4480), 
            .I2(n2669), .I3(GND_net), .O(n2736));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1622 (.I0(n1647_adj_4482), .I1(n1646_adj_4481), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4921));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i1_2_lut_adj_1622.LUT_INIT = 16'heeee;
    SB_LUT4 rem_4_i1455_3_lut (.I0(n2142), .I1(n2209), .I2(n2174_adj_4597), 
            .I3(GND_net), .O(n2241));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1459_3_lut (.I0(n2146), .I1(n2213), .I2(n2174_adj_4597), 
            .I3(GND_net), .O(n2245));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1457_3_lut (.I0(n2144), .I1(n2211), .I2(n2174_adj_4597), 
            .I3(GND_net), .O(n2243));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1458_3_lut (.I0(n2145), .I1(n2212), .I2(n2174_adj_4597), 
            .I3(GND_net), .O(n2244));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1854_12_lut (.I0(GND_net), .I1(n2749), .I2(VCC_net), 
            .I3(n31032), .O(n2816_adj_4461)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1809_3_lut (.I0(n2656), .I1(n2723_adj_4463), .I2(n2669), 
            .I3(GND_net), .O(n2755));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1809_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1854_12 (.CI(n31032), .I0(n2749), .I1(VCC_net), 
            .CO(n31033));
    SB_LUT4 rem_4_i1456_3_lut (.I0(n2143), .I1(n2210), .I2(n2174_adj_4597), 
            .I3(GND_net), .O(n2242));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1452_14_lut (.I0(GND_net), .I1(n2147), .I2(VCC_net), 
            .I3(n31304), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_14 (.CI(n31304), .I0(n2147), .I1(VCC_net), 
            .CO(n31305));
    SB_LUT4 rem_4_i1469_3_lut (.I0(n2156), .I1(n2223), .I2(n2174_adj_4597), 
            .I3(GND_net), .O(n2255));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1468_3_lut (.I0(n2155), .I1(n2222), .I2(n2174_adj_4597), 
            .I3(GND_net), .O(n2254));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1460_3_lut (.I0(n2147), .I1(n2214), .I2(n2174_adj_4597), 
            .I3(GND_net), .O(n2246));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1471_3_lut (.I0(n2158), .I1(n2225), .I2(n2174_adj_4597), 
            .I3(GND_net), .O(n2257));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1470_3_lut (.I0(n2157), .I1(n2224), .I2(n2174_adj_4597), 
            .I3(GND_net), .O(n2256));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1391_3_lut (.I0(n2046), .I1(n2113), .I2(n2075_adj_4609), 
            .I3(GND_net), .O(n2145));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1389_3_lut (.I0(n2044), .I1(n2111), .I2(n2075_adj_4609), 
            .I3(GND_net), .O(n2143));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1390_3_lut (.I0(n2045), .I1(n2112), .I2(n2075_adj_4609), 
            .I3(GND_net), .O(n2144));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1623 (.I0(n1656), .I1(n1657), .I2(n1658), .I3(GND_net), 
            .O(n38287));
    defparam i1_3_lut_adj_1623.LUT_INIT = 16'hfefe;
    SB_LUT4 i7_4_lut_adj_1624 (.I0(n1653_adj_4488), .I1(n1652_adj_4487), 
            .I2(n1651_adj_4486), .I3(n10_adj_4921), .O(n16_adj_4919));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i7_4_lut_adj_1624.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(n1648_adj_4483), .I1(n1654), .I2(n38287), .I3(n1655), 
            .O(n11_adj_4920));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i2_4_lut.LUT_INIT = 16'heaaa;
    SB_LUT4 i8_4_lut (.I0(n11_adj_4920), .I1(n16_adj_4919), .I2(n1649_adj_4484), 
            .I3(n1650_adj_4485), .O(n1679));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i20_3_lut (.I0(communication_counter[19]), .I1(n14_adj_4398), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1658));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i21_3_lut (.I0(communication_counter[20]), .I1(n13_adj_4399), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1558));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i995_3_lut (.I0(n1458), .I1(n1525), .I2(n1481), .I3(GND_net), 
            .O(n1557));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1388_3_lut (.I0(n2043), .I1(n2110), .I2(n2075_adj_4609), 
            .I3(GND_net), .O(n2142));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1397_3_lut (.I0(n2052), .I1(n2119), .I2(n2075_adj_4609), 
            .I3(GND_net), .O(n2151));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1399_3_lut (.I0(n2054), .I1(n2121), .I2(n2075_adj_4609), 
            .I3(GND_net), .O(n2153));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1394_3_lut (.I0(n2049), .I1(n2116), .I2(n2075_adj_4609), 
            .I3(GND_net), .O(n2148));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i994_3_lut (.I0(n1457), .I1(n1524), .I2(n1481), .I3(GND_net), 
            .O(n1556));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1395_3_lut (.I0(n2050), .I1(n2117), .I2(n2075_adj_4609), 
            .I3(GND_net), .O(n2149));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1393_3_lut (.I0(n2048), .I1(n2115), .I2(n2075_adj_4609), 
            .I3(GND_net), .O(n2147));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1398_3_lut (.I0(n2053), .I1(n2120), .I2(n2075_adj_4609), 
            .I3(GND_net), .O(n2152));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1392_3_lut (.I0(n2047), .I1(n2114), .I2(n2075_adj_4609), 
            .I3(GND_net), .O(n2146));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1331_3_lut (.I0(n1954), .I1(n2021), .I2(n1976_adj_4627), 
            .I3(GND_net), .O(n2053));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1327_3_lut (.I0(n1950), .I1(n2017), .I2(n1976_adj_4627), 
            .I3(GND_net), .O(n2049));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1323_3_lut (.I0(n1946), .I1(n2013), .I2(n1976_adj_4627), 
            .I3(GND_net), .O(n2045));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1322_3_lut (.I0(n1945), .I1(n2012), .I2(n1976_adj_4627), 
            .I3(GND_net), .O(n2044));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1321_3_lut (.I0(n1944), .I1(n2011), .I2(n1976_adj_4627), 
            .I3(GND_net), .O(n2043));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1328_3_lut (.I0(n1951), .I1(n2018), .I2(n1976_adj_4627), 
            .I3(GND_net), .O(n2050));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1329_3_lut (.I0(n1952), .I1(n2019), .I2(n1976_adj_4627), 
            .I3(GND_net), .O(n2051));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1326_3_lut (.I0(n1949), .I1(n2016), .I2(n1976_adj_4627), 
            .I3(GND_net), .O(n2048));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1330_3_lut (.I0(n1953), .I1(n2020), .I2(n1976_adj_4627), 
            .I3(GND_net), .O(n2052));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1325_3_lut (.I0(n1948), .I1(n2015), .I2(n1976_adj_4627), 
            .I3(GND_net), .O(n2047));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1333_3_lut (.I0(n1956), .I1(n2023), .I2(n1976_adj_4627), 
            .I3(GND_net), .O(n2055));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1332_3_lut (.I0(n1955), .I1(n2022), .I2(n1976_adj_4627), 
            .I3(GND_net), .O(n2054));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1324_3_lut (.I0(n1947), .I1(n2014), .I2(n1976_adj_4627), 
            .I3(GND_net), .O(n2046));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1257_3_lut (.I0(n1848), .I1(n1915), .I2(n1877), .I3(GND_net), 
            .O(n1947));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1258_3_lut (.I0(n1849), .I1(n1916), .I2(n1877), .I3(GND_net), 
            .O(n1948));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1261_3_lut (.I0(n1852), .I1(n1919), .I2(n1877), .I3(GND_net), 
            .O(n1951));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1854_11_lut (.I0(GND_net), .I1(n2750), .I2(VCC_net), 
            .I3(n31031), .O(n2817_adj_4460)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_13_lut (.I0(GND_net), .I1(n2148), .I2(VCC_net), 
            .I3(n31303), .O(n2215)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_11 (.CI(n31031), .I0(n2750), .I1(VCC_net), 
            .CO(n31032));
    SB_CARRY rem_4_add_1452_13 (.CI(n31303), .I0(n2148), .I1(VCC_net), 
            .CO(n31304));
    SB_LUT4 div_36_i1704_3_lut_3_lut (.I0(n2558), .I1(n7118), .I2(n2539), 
            .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1704_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1452_12_lut (.I0(GND_net), .I1(n2149), .I2(VCC_net), 
            .I3(n31302), .O(n2216)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i460_4_lut_4_lut (.I0(n671), .I1(n99), .I2(n2_adj_4907), 
            .I3(n649), .O(n784));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i460_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 rem_4_i1263_3_lut (.I0(n1854), .I1(n1921), .I2(n1877), .I3(GND_net), 
            .O(n1953));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1256_3_lut (.I0(n1847), .I1(n1914), .I2(n1877), .I3(GND_net), 
            .O(n1946));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1854_10_lut (.I0(GND_net), .I1(n2751), .I2(VCC_net), 
            .I3(n31030), .O(n2818_adj_4459)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1808_3_lut (.I0(n2655), .I1(n2722), .I2(n2669), .I3(GND_net), 
            .O(n2754));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1808_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1255_3_lut (.I0(n1846), .I1(n1913), .I2(n1877), .I3(GND_net), 
            .O(n1945));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i458_4_lut_4_lut (.I0(n671), .I1(n97), .I2(n6_adj_4438), 
            .I3(n38024), .O(n38026));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i458_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_CARRY rem_4_add_1854_10 (.CI(n31030), .I0(n2751), .I1(VCC_net), 
            .CO(n31031));
    SB_CARRY rem_4_add_1452_12 (.CI(n31302), .I0(n2149), .I1(VCC_net), 
            .CO(n31303));
    SB_LUT4 rem_4_add_1854_9_lut (.I0(GND_net), .I1(n2752), .I2(VCC_net), 
            .I3(n31029), .O(n2819_adj_4458)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_9 (.CI(n31029), .I0(n2752), .I1(VCC_net), 
            .CO(n31030));
    SB_LUT4 rem_4_i1254_3_lut (.I0(n1845), .I1(n1912), .I2(n1877), .I3(GND_net), 
            .O(n1944));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1254_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1854_8_lut (.I0(GND_net), .I1(n2753), .I2(VCC_net), 
            .I3(n31028), .O(n2820_adj_4457)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_11_lut (.I0(GND_net), .I1(n2150), .I2(VCC_net), 
            .I3(n31301), .O(n2217)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_8 (.CI(n31028), .I0(n2753), .I1(VCC_net), 
            .CO(n31029));
    SB_CARRY rem_4_add_1452_11 (.CI(n31301), .I0(n2150), .I1(VCC_net), 
            .CO(n31302));
    SB_LUT4 rem_4_i1794_3_lut (.I0(n2641), .I1(n2708_adj_4476), .I2(n2669), 
            .I3(GND_net), .O(n2740));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1452_10_lut (.I0(GND_net), .I1(n2151), .I2(VCC_net), 
            .I3(n31300), .O(n2218)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_7_lut (.I0(GND_net), .I1(n2754), .I2(GND_net), 
            .I3(n31027), .O(n2821_adj_4456)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1811_3_lut (.I0(n2658), .I1(n2725), .I2(n2669), .I3(GND_net), 
            .O(n2757));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1811_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1854_7 (.CI(n31027), .I0(n2754), .I1(GND_net), 
            .CO(n31028));
    SB_LUT4 i36499_3_lut_3_lut (.I0(n671), .I1(n558), .I2(n371), .I3(GND_net), 
            .O(n785));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36499_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 rem_4_add_1854_6_lut (.I0(GND_net), .I1(n2755), .I2(GND_net), 
            .I3(n31026), .O(n2822_adj_4455)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1810_3_lut (.I0(n2657), .I1(n2724_adj_4462), .I2(n2669), 
            .I3(GND_net), .O(n2756));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1262_3_lut (.I0(n1853), .I1(n1920), .I2(n1877), .I3(GND_net), 
            .O(n1952));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1262_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1452_10 (.CI(n31300), .I0(n2151), .I1(VCC_net), 
            .CO(n31301));
    SB_LUT4 rem_4_add_1452_9_lut (.I0(GND_net), .I1(n2152), .I2(VCC_net), 
            .I3(n31299), .O(n2219)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_6 (.CI(n31026), .I0(n2755), .I1(GND_net), 
            .CO(n31027));
    SB_CARRY rem_4_add_1452_9 (.CI(n31299), .I0(n2152), .I1(VCC_net), 
            .CO(n31300));
    SB_LUT4 rem_4_add_1854_5_lut (.I0(GND_net), .I1(n2756), .I2(VCC_net), 
            .I3(n31025), .O(n2823_adj_4454)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_5 (.CI(n31025), .I0(n2756), .I1(VCC_net), 
            .CO(n31026));
    SB_LUT4 i1_3_lut_adj_1625 (.I0(n2756), .I1(n2757), .I2(n2758), .I3(GND_net), 
            .O(n38326));
    defparam i1_3_lut_adj_1625.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_add_1854_4_lut (.I0(GND_net), .I1(n2757), .I2(VCC_net), 
            .I3(n31024), .O(n2824_adj_4453)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_8_lut (.I0(GND_net), .I1(n2153), .I2(VCC_net), 
            .I3(n31298), .O(n2220)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_8 (.CI(n31298), .I0(n2153), .I1(VCC_net), 
            .CO(n31299));
    SB_LUT4 rem_4_add_1452_7_lut (.I0(GND_net), .I1(n2154), .I2(GND_net), 
            .I3(n31297), .O(n2221)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_4 (.CI(n31024), .I0(n2757), .I1(VCC_net), 
            .CO(n31025));
    SB_LUT4 rem_4_add_1854_3_lut (.I0(GND_net), .I1(n2758), .I2(GND_net), 
            .I3(n31023), .O(n2825_adj_4452)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_7 (.CI(n31297), .I0(n2154), .I1(GND_net), 
            .CO(n31298));
    SB_LUT4 add_7258_7_lut (.I0(n40287), .I1(n746), .I2(GND_net), .I3(n32338), 
            .O(n39906)) /* synthesis syn_instantiated=1 */ ;
    defparam add_7258_7_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 rem_4_i1259_3_lut (.I0(n1850), .I1(n1917), .I2(n1877), .I3(GND_net), 
            .O(n1949));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1452_6_lut (.I0(GND_net), .I1(n2155), .I2(GND_net), 
            .I3(n31296), .O(n2222)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1267_3_lut (.I0(n1858), .I1(n1925), .I2(n1877), .I3(GND_net), 
            .O(n1957));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_1626 (.I0(n2740), .I1(n2754), .I2(n38326), .I3(n2755), 
            .O(n24_adj_4975));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i4_4_lut_adj_1626.LUT_INIT = 16'heaaa;
    SB_LUT4 i11_4_lut (.I0(n2736), .I1(n2737), .I2(n2735), .I3(n2738), 
            .O(n31_adj_4974));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1627 (.I0(n31_adj_4974), .I1(n2739), .I2(n24_adj_4975), 
            .I3(n2742), .O(n36_adj_4970));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i16_4_lut_adj_1627.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n2752), .I1(n2748), .I2(n2744), .I3(n2745), 
            .O(n34_adj_4972));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1854_3 (.CI(n31023), .I0(n2758), .I1(GND_net), 
            .CO(n31024));
    SB_CARRY rem_4_add_1452_6 (.CI(n31296), .I0(n2155), .I1(GND_net), 
            .CO(n31297));
    SB_CARRY rem_4_add_1854_2 (.CI(VCC_net), .I0(n2858), .I1(VCC_net), 
            .CO(n31023));
    SB_LUT4 rem_4_add_1921_26_lut (.I0(n2867_adj_4441), .I1(n2834_adj_4451), 
            .I2(VCC_net), .I3(n31022), .O(n2933)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1452_5_lut (.I0(GND_net), .I1(n2156), .I2(VCC_net), 
            .I3(n31295), .O(n2223)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1266_rep_57_3_lut (.I0(n1857), .I1(n1924), .I2(n1877), 
            .I3(GND_net), .O(n1956));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1266_rep_57_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1921_25_lut (.I0(GND_net), .I1(n2835_adj_4450), .I2(VCC_net), 
            .I3(n31021), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_25 (.CI(n31021), .I0(n2835_adj_4450), .I1(VCC_net), 
            .CO(n31022));
    SB_LUT4 rem_4_add_1921_24_lut (.I0(GND_net), .I1(n2836_adj_4449), .I2(VCC_net), 
            .I3(n31020), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_24 (.CI(n31020), .I0(n2836_adj_4449), .I1(VCC_net), 
            .CO(n31021));
    SB_LUT4 add_7258_6_lut (.I0(GND_net), .I1(n852), .I2(GND_net), .I3(n32337), 
            .O(n12165)) /* synthesis syn_instantiated=1 */ ;
    defparam add_7258_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_5 (.CI(n31295), .I0(n2156), .I1(VCC_net), 
            .CO(n31296));
    SB_LUT4 rem_4_add_1452_4_lut (.I0(GND_net), .I1(n2157), .I2(VCC_net), 
            .I3(n31294), .O(n2224)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_4 (.CI(n31294), .I0(n2157), .I1(VCC_net), 
            .CO(n31295));
    SB_CARRY add_7258_6 (.CI(n32337), .I0(n852), .I1(GND_net), .CO(n32338));
    SB_LUT4 rem_4_add_1452_3_lut (.I0(GND_net), .I1(n2158), .I2(GND_net), 
            .I3(n31293), .O(n2225)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15_4_lut_adj_1628 (.I0(n2753), .I1(n2749), .I2(n2746), .I3(n2747), 
            .O(n35_adj_4971));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i15_4_lut_adj_1628.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1629 (.I0(n2741), .I1(n2743), .I2(n2750), .I3(n2751), 
            .O(n33_adj_4973));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i13_4_lut_adj_1629.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n33_adj_4973), .I1(n35_adj_4971), .I2(n34_adj_4972), 
            .I3(n36_adj_4970), .O(n2768));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i9_3_lut (.I0(communication_counter[8]), .I1(n25_adj_4385), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2758));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1452_3 (.CI(n31293), .I0(n2158), .I1(GND_net), 
            .CO(n31294));
    SB_LUT4 i37439_3_lut (.I0(n1652_adj_4487), .I1(n1719), .I2(n1679), 
            .I3(GND_net), .O(n1751));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i37439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_7258_5_lut (.I0(GND_net), .I1(n748), .I2(VCC_net), .I3(n32336), 
            .O(n12166)) /* synthesis syn_instantiated=1 */ ;
    defparam add_7258_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_2 (.CI(VCC_net), .I0(n2258), .I1(VCC_net), 
            .CO(n31293));
    SB_CARRY add_7258_5 (.CI(n32336), .I0(n748), .I1(VCC_net), .CO(n32337));
    SB_LUT4 rem_4_add_1519_21_lut (.I0(n2273_adj_4591), .I1(n2240), .I2(VCC_net), 
            .I3(n31292), .O(n2339)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1921_23_lut (.I0(GND_net), .I1(n2837_adj_4448), .I2(VCC_net), 
            .I3(n31019), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_7258_4_lut (.I0(GND_net), .I1(n749), .I2(VCC_net), .I3(n32335), 
            .O(n12167)) /* synthesis syn_instantiated=1 */ ;
    defparam add_7258_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37263_3_lut (.I0(n1751), .I1(n1818), .I2(n1778_adj_4738), 
            .I3(GND_net), .O(n1850));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i37263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1191_3_lut (.I0(n1750), .I1(n1817), .I2(n1778_adj_4738), 
            .I3(GND_net), .O(n1849));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1194_3_lut (.I0(n1753), .I1(n1820), .I2(n1778_adj_4738), 
            .I3(GND_net), .O(n1852));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i459_4_lut_4_lut (.I0(n671), .I1(n98), .I2(n4_adj_4443), 
            .I3(n648), .O(n783));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i459_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 rem_4_i1195_rep_58_3_lut (.I0(n1754_adj_4785), .I1(n1821), .I2(n1778_adj_4738), 
            .I3(GND_net), .O(n1853));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1195_rep_58_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1190_3_lut (.I0(n1749), .I1(n1816), .I2(n1778_adj_4738), 
            .I3(GND_net), .O(n1848));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1189_3_lut (.I0(n1748), .I1(n1815), .I2(n1778_adj_4738), 
            .I3(GND_net), .O(n1847));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1519_20_lut (.I0(GND_net), .I1(n2241), .I2(VCC_net), 
            .I3(n31291), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_23 (.CI(n31019), .I0(n2837_adj_4448), .I1(VCC_net), 
            .CO(n31020));
    SB_CARRY add_7258_4 (.CI(n32335), .I0(n749), .I1(VCC_net), .CO(n32336));
    SB_LUT4 rem_4_i1188_3_lut (.I0(n1747), .I1(n1814), .I2(n1778_adj_4738), 
            .I3(GND_net), .O(n1846));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1188_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1519_20 (.CI(n31291), .I0(n2241), .I1(VCC_net), 
            .CO(n31292));
    SB_LUT4 rem_4_add_1519_19_lut (.I0(GND_net), .I1(n2242), .I2(VCC_net), 
            .I3(n31290), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_7258_3_lut (.I0(GND_net), .I1(n855), .I2(GND_net), .I3(n32334), 
            .O(n12168)) /* synthesis syn_instantiated=1 */ ;
    defparam add_7258_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_19 (.CI(n31290), .I0(n2242), .I1(VCC_net), 
            .CO(n31291));
    SB_CARRY add_7258_3 (.CI(n32334), .I0(n855), .I1(GND_net), .CO(n32335));
    SB_LUT4 rem_4_i1199_3_lut (.I0(n1758_adj_4781), .I1(n1825), .I2(n1778_adj_4738), 
            .I3(GND_net), .O(n1857));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1197_3_lut (.I0(n1756_adj_4783), .I1(n1823), .I2(n1778_adj_4738), 
            .I3(GND_net), .O(n1855));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1197_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_7258_2 (.CI(VCC_net), .I0(n958), .I1(VCC_net), .CO(n32334));
    SB_LUT4 rem_4_unary_minus_2_add_3_33_lut (.I0(communication_counter[31]), 
            .I1(GND_net), .I2(n2_adj_4938), .I3(n32333), .O(n746)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_unary_minus_2_add_3_32_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4939), .I3(n32332), .O(n3_adj_4409)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_18_lut (.I0(GND_net), .I1(n2243), .I2(VCC_net), 
            .I3(n31289), .O(n2310)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_18 (.CI(n31289), .I0(n2243), .I1(VCC_net), 
            .CO(n31290));
    SB_LUT4 rem_4_add_1921_22_lut (.I0(GND_net), .I1(n2838_adj_4447), .I2(VCC_net), 
            .I3(n31018), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_17_lut (.I0(GND_net), .I1(n2244), .I2(VCC_net), 
            .I3(n31288), .O(n2311)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4430));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_i1703_3_lut_3_lut (.I0(n2558), .I1(n7117), .I2(n2538), 
            .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1703_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1196_3_lut (.I0(n1755_adj_4784), .I1(n1822), .I2(n1778_adj_4738), 
            .I3(GND_net), .O(n1854));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i18_3_lut (.I0(communication_counter[17]), .I1(n16_adj_4396), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1858));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_unary_minus_2_add_3_32 (.CI(n32332), .I0(GND_net), .I1(n3_adj_4939), 
            .CO(n32333));
    SB_LUT4 rem_4_i1124_3_lut (.I0(n1651_adj_4486), .I1(n1718), .I2(n1679), 
            .I3(GND_net), .O(n1750));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1124_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1519_17 (.CI(n31288), .I0(n2244), .I1(VCC_net), 
            .CO(n31289));
    SB_LUT4 rem_4_i1126_3_lut (.I0(n1653_adj_4488), .I1(n1720), .I2(n1679), 
            .I3(GND_net), .O(n1752));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1129_3_lut (.I0(n1656), .I1(n1723), .I2(n1679), .I3(GND_net), 
            .O(n1755_adj_4784));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_add_3_31_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4940), .I3(n32331), .O(n4_adj_4408)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1123_3_lut (.I0(n1650_adj_4485), .I1(n1717), .I2(n1679), 
            .I3(GND_net), .O(n1749));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1123_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_22 (.CI(n31018), .I0(n2838_adj_4447), .I1(VCC_net), 
            .CO(n31019));
    SB_LUT4 rem_4_i1128_3_lut (.I0(n1655), .I1(n1722), .I2(n1679), .I3(GND_net), 
            .O(n1754_adj_4785));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37266_3_lut (.I0(n1553_adj_4493), .I1(n1620), .I2(n1580), 
            .I3(GND_net), .O(n1652_adj_4487));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i37266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1127_3_lut (.I0(n1654), .I1(n1721), .I2(n1679), .I3(GND_net), 
            .O(n1753));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1122_3_lut (.I0(n1649_adj_4484), .I1(n1716), .I2(n1679), 
            .I3(GND_net), .O(n1748));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1122_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_unary_minus_2_add_3_31 (.CI(n32331), .I0(GND_net), .I1(n4_adj_4940), 
            .CO(n32332));
    SB_LUT4 rem_4_i1121_3_lut (.I0(n1648_adj_4483), .I1(n1715), .I2(n1679), 
            .I3(GND_net), .O(n1747));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i19_3_lut (.I0(communication_counter[18]), .I1(n15_adj_4397), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1758_adj_4781));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_add_3_30_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4941), .I3(n32330), .O(n5_adj_4407)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i549_4_lut_4_lut (.I0(n806), .I1(n98), .I2(n4_adj_4349), 
            .I3(n784), .O(n916));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i549_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 rem_4_i1131_3_lut (.I0(n1658), .I1(n1725), .I2(n1679), .I3(GND_net), 
            .O(n1757_adj_4782));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13987_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n14536), .I3(GND_net), .O(n19019));   // verilog/coms.v(126[12] 289[6])
    defparam i13987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4429));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_unary_minus_2_add_3_30 (.CI(n32330), .I0(GND_net), .I1(n5_adj_4941), 
            .CO(n32331));
    SB_LUT4 rem_4_unary_minus_2_add_3_29_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4942), .I3(n32329), .O(n6_adj_4406)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1130_3_lut (.I0(n1657), .I1(n1724), .I2(n1679), .I3(GND_net), 
            .O(n1756_adj_4783));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1630 (.I0(n1746), .I1(n1747), .I2(n1745), .I3(n1748), 
            .O(n16));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i6_4_lut_adj_1630.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1631 (.I0(n1756_adj_4783), .I1(n1757_adj_4782), 
            .I2(n1758_adj_4781), .I3(GND_net), .O(n38279));
    defparam i1_3_lut_adj_1631.LUT_INIT = 16'hfefe;
    SB_LUT4 i8_3_lut (.I0(n1753), .I1(n16), .I2(n1751), .I3(GND_net), 
            .O(n18));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i8_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1632 (.I0(n1754_adj_4785), .I1(n1749), .I2(n38279), 
            .I3(n1755_adj_4784), .O(n13));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i3_4_lut_adj_1632.LUT_INIT = 16'heccc;
    SB_LUT4 div_36_i1715_3_lut_3_lut (.I0(n2558), .I1(n7129), .I2(n2550), 
            .I3(GND_net), .O(n2634));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1715_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i550_4_lut_4_lut (.I0(n806), .I1(n99), .I2(n2_adj_4434), 
            .I3(n785), .O(n917));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i550_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i9_4_lut (.I0(n13), .I1(n18), .I2(n1752), .I3(n1750), .O(n1778_adj_4738));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1120_3_lut (.I0(n1647_adj_4482), .I1(n1714), .I2(n1679), 
            .I3(GND_net), .O(n1746));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1120_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_unary_minus_2_add_3_29 (.CI(n32329), .I0(GND_net), .I1(n6_adj_4942), 
            .CO(n32330));
    SB_LUT4 div_36_i547_4_lut_4_lut (.I0(n806), .I1(n96), .I2(n8_adj_4346), 
            .I3(n38026), .O(n914));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i547_4_lut_4_lut.LUT_INIT = 16'h14eb;
    SB_LUT4 rem_4_i1187_3_lut (.I0(n1746), .I1(n1813), .I2(n1778_adj_4738), 
            .I3(GND_net), .O(n1845));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1921_21_lut (.I0(GND_net), .I1(n2839_adj_4446), .I2(VCC_net), 
            .I3(n31017), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37261_3_lut (.I0(n1752), .I1(n1819), .I2(n1778_adj_4738), 
            .I3(GND_net), .O(n1851));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i37261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i548_4_lut_4_lut (.I0(n806), .I1(n97), .I2(n6_adj_4348), 
            .I3(n783), .O(n915));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i548_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i36490_3_lut_3_lut (.I0(n806), .I1(n558), .I2(n372), .I3(GND_net), 
            .O(n918));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36490_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 i1_2_lut_adj_1633 (.I0(n1856), .I1(n1858), .I2(GND_net), .I3(GND_net), 
            .O(n40501));
    defparam i1_2_lut_adj_1633.LUT_INIT = 16'heeee;
    SB_CARRY rem_4_add_1921_21 (.CI(n31017), .I0(n2839_adj_4446), .I1(VCC_net), 
            .CO(n31018));
    SB_LUT4 i1_4_lut_adj_1634 (.I0(n1854), .I1(n40501), .I2(n1855), .I3(n1857), 
            .O(n38306));
    defparam i1_4_lut_adj_1634.LUT_INIT = 16'ha080;
    SB_LUT4 i7_4_lut_adj_1635 (.I0(n1846), .I1(n38306), .I2(n1847), .I3(n1848), 
            .O(n18_adj_4936));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i7_4_lut_adj_1635.LUT_INIT = 16'hfffe;
    SB_LUT4 div_36_i1713_3_lut_3_lut (.I0(n2558), .I1(n7127), .I2(n2548), 
            .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1713_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i637_3_lut_3_lut (.I0(n938), .I1(n6890), .I2(n917), 
            .I3(GND_net), .O(n1046));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i637_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i638_3_lut_3_lut (.I0(n938), .I1(n6891), .I2(n918), 
            .I3(GND_net), .O(n1047));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i638_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i5_2_lut (.I0(n1853), .I1(n1852), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4937));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1636 (.I0(n1851), .I1(n18_adj_4936), .I2(n1845), 
            .I3(n1844), .O(n20_adj_4935));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i9_4_lut_adj_1636.LUT_INIT = 16'hfffe;
    SB_LUT4 i13720_2_lut (.I0(n18897), .I1(n18750), .I2(GND_net), .I3(GND_net), 
            .O(n18752));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13720_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13717_2_lut (.I0(n18897), .I1(n18747), .I2(GND_net), .I3(GND_net), 
            .O(n18749));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13717_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 rem_4_add_1921_20_lut (.I0(GND_net), .I1(n2840), .I2(VCC_net), 
            .I3(n31016), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i993_3_lut (.I0(n1456), .I1(n1523), .I2(n1481), .I3(GND_net), 
            .O(n1555));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i993_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_20 (.CI(n31016), .I0(n2840), .I1(VCC_net), 
            .CO(n31017));
    SB_LUT4 rem_4_add_1519_16_lut (.I0(GND_net), .I1(n2245), .I2(VCC_net), 
            .I3(n31287), .O(n2312)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10_4_lut_adj_1637 (.I0(n1849), .I1(n20_adj_4935), .I2(n16_adj_4937), 
            .I3(n1850), .O(n1877));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i10_4_lut_adj_1637.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_3_lut (.I0(n1105), .I1(n38070), .I2(state[0]), .I3(GND_net), 
            .O(n19_adj_4910));   // verilog/neopixel.v(35[12] 117[6])
    defparam i27_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_36_i639_3_lut_3_lut (.I0(n938), .I1(n6892), .I2(n373), 
            .I3(GND_net), .O(n1048));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i639_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1198_3_lut (.I0(n1757_adj_4782), .I1(n1824), .I2(n1778_adj_4738), 
            .I3(GND_net), .O(n1856));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13988_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n14536), .I3(GND_net), .O(n19020));   // verilog/coms.v(126[12] 289[6])
    defparam i13988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_add_3_28_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4943), .I3(n32328), .O(n7_adj_4405)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1265_3_lut (.I0(n1856), .I1(n1923), .I2(n1877), .I3(GND_net), 
            .O(n1955));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1265_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1260_3_lut (.I0(n1851), .I1(n1918), .I2(n1877), .I3(GND_net), 
            .O(n1950));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1264_3_lut (.I0(n1855), .I1(n1922), .I2(n1877), .I3(GND_net), 
            .O(n1954));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1638 (.I0(n1956), .I1(n1957), .I2(n1958), .I3(GND_net), 
            .O(n38295));
    defparam i1_3_lut_adj_1638.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_1639 (.I0(n1954), .I1(n1950), .I2(n38295), .I3(n1955), 
            .O(n16_adj_4739));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i4_4_lut_adj_1639.LUT_INIT = 16'heccc;
    SB_LUT4 i7_4_lut_adj_1640 (.I0(n1944), .I1(n1945), .I2(n1943), .I3(n1946), 
            .O(n19_adj_4699));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i7_4_lut_adj_1640.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1519_16 (.CI(n31287), .I0(n2245), .I1(VCC_net), 
            .CO(n31288));
    SB_LUT4 i6_2_lut (.I0(n1953), .I1(n1951), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4717));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1641 (.I0(n19_adj_4699), .I1(n1948), .I2(n16_adj_4739), 
            .I3(n1947), .O(n22_adj_4681));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i10_4_lut_adj_1641.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1642 (.I0(n1949), .I1(n22_adj_4681), .I2(n18_adj_4717), 
            .I3(n1952), .O(n1976_adj_4627));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i11_4_lut_adj_1642.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_unary_minus_2_add_3_28 (.CI(n32328), .I0(GND_net), .I1(n7_adj_4943), 
            .CO(n32329));
    SB_LUT4 rem_4_mux_3_i17_3_lut (.I0(communication_counter[16]), .I1(n17_adj_4395), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1958));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_IO PIN_8_pad (.PACKAGE_PIN(PIN_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_8_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_8_pad.PIN_TYPE = 6'b011001;
    defparam PIN_8_pad.PULLUP = 1'b0;
    defparam PIN_8_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_13_pad (.PACKAGE_PIN(PIN_13), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_13_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_13_pad.PIN_TYPE = 6'b000001;
    defparam PIN_13_pad.PULLUP = 1'b0;
    defparam PIN_13_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_36_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4567));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13989_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n14536), .I3(GND_net), .O(n19021));   // verilog/coms.v(126[12] 289[6])
    defparam i13989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1335_3_lut (.I0(n1958), .I1(n2025), .I2(n1976_adj_4627), 
            .I3(GND_net), .O(n2057));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1334_3_lut (.I0(n1957), .I1(n2024), .I2(n1976_adj_4627), 
            .I3(GND_net), .O(n2056));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1643 (.I0(n2056), .I1(n2057), .I2(n2058), .I3(GND_net), 
            .O(n38338));
    defparam i1_3_lut_adj_1643.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1644 (.I0(n2046), .I1(n2054), .I2(n38338), .I3(n2055), 
            .O(n16_adj_4357));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i3_4_lut_adj_1644.LUT_INIT = 16'heaaa;
    SB_LUT4 rem_4_add_1519_15_lut (.I0(GND_net), .I1(n2246), .I2(VCC_net), 
            .I3(n31286), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_15 (.CI(n31286), .I0(n2246), .I1(VCC_net), 
            .CO(n31287));
    SB_LUT4 i9_4_lut_adj_1645 (.I0(n2047), .I1(n2052), .I2(n2048), .I3(n2051), 
            .O(n22_adj_4355));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i9_4_lut_adj_1645.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1519_14_lut (.I0(GND_net), .I1(n2247), .I2(VCC_net), 
            .I3(n31285), .O(n2314)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_19_lut (.I0(GND_net), .I1(n2841), .I2(VCC_net), 
            .I3(n31015), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_3_lut (.I0(n2050), .I1(n2043), .I2(n2042), .I3(GND_net), 
            .O(n20_adj_4356));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1646 (.I0(n2044), .I1(n22_adj_4355), .I2(n16_adj_4357), 
            .I3(n2045), .O(n24_adj_4354));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i11_4_lut_adj_1646.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1647 (.I0(n2049), .I1(n24_adj_4354), .I2(n20_adj_4356), 
            .I3(n2053), .O(n2075_adj_4609));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i12_4_lut_adj_1647.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i16_3_lut (.I0(communication_counter[15]), .I1(n18_adj_4394), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2058));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF color__i19 (.Q(color[21]), .C(LED_c), .D(n18940));   // verilog/TinyFPGA_B.v(48[8] 62[4])
    SB_LUT4 rem_4_i1403_3_lut (.I0(n2058), .I1(n2125), .I2(n2075_adj_4609), 
            .I3(GND_net), .O(n2157));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1403_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_19 (.CI(n31015), .I0(n2841), .I1(VCC_net), 
            .CO(n31016));
    SB_LUT4 div_36_i636_3_lut_3_lut (.I0(n938), .I1(n6889), .I2(n916), 
            .I3(GND_net), .O(n1045));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i636_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4566));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1401_3_lut (.I0(n2056), .I1(n2123), .I2(n2075_adj_4609), 
            .I3(GND_net), .O(n2155));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1400_3_lut (.I0(n2055), .I1(n2122), .I2(n2075_adj_4609), 
            .I3(GND_net), .O(n2154));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i15_3_lut (.I0(communication_counter[14]), .I1(n19_adj_4393), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2158));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1402_3_lut (.I0(n2057), .I1(n2124), .I2(n2075_adj_4609), 
            .I3(GND_net), .O(n2156));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1648 (.I0(n2156), .I1(n2158), .I2(GND_net), .I3(GND_net), 
            .O(n40407));
    defparam i1_2_lut_adj_1648.LUT_INIT = 16'heeee;
    SB_LUT4 div_36_i635_3_lut_3_lut (.I0(n938), .I1(n6888), .I2(n915), 
            .I3(GND_net), .O(n1044));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i635_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_unary_minus_2_add_3_27_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4944), .I3(n32327), .O(n8_adj_4404)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_18_lut (.I0(GND_net), .I1(n2842), .I2(VCC_net), 
            .I3(n31014), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_18 (.CI(n31014), .I0(n2842), .I1(VCC_net), 
            .CO(n31015));
    SB_DFF color__i18 (.Q(color[20]), .C(LED_c), .D(n18939));   // verilog/TinyFPGA_B.v(48[8] 62[4])
    SB_LUT4 i1_4_lut_adj_1649 (.I0(n2154), .I1(n40407), .I2(n2155), .I3(n2157), 
            .O(n38299));
    defparam i1_4_lut_adj_1649.LUT_INIT = 16'ha080;
    SB_LUT4 i4_2_lut (.I0(n2150), .I1(n2146), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4986));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_36_i634_3_lut_3_lut (.I0(n938), .I1(n6887), .I2(n914), 
            .I3(GND_net), .O(n1043));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i634_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1921_17_lut (.I0(GND_net), .I1(n2843), .I2(VCC_net), 
            .I3(n31013), .O(n2910)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4565));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_DFF color__i17 (.Q(color[17]), .C(LED_c), .D(n18938));   // verilog/TinyFPGA_B.v(48[8] 62[4])
    SB_CARRY rem_4_add_1921_17 (.CI(n31013), .I0(n2843), .I1(VCC_net), 
            .CO(n31014));
    SB_LUT4 div_36_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4564));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_570_i42_3_lut_3_lut (.I0(n916), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n42_adj_4594));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_570_i42_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i36100_3_lut_4_lut (.I0(n916), .I1(n97), .I2(n98), .I3(n917), 
            .O(n43224));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36100_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_CARRY rem_4_unary_minus_2_add_3_27 (.CI(n32327), .I0(GND_net), .I1(n8_adj_4944), 
            .CO(n32328));
    SB_LUT4 rem_4_add_1921_16_lut (.I0(GND_net), .I1(n2844), .I2(VCC_net), 
            .I3(n31012), .O(n2911)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10_4_lut_adj_1650 (.I0(n2152), .I1(n2147), .I2(n2149), .I3(n2148), 
            .O(n24_adj_4984));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i10_4_lut_adj_1650.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1651 (.I0(n2142), .I1(n2144), .I2(n2141), .I3(n38299), 
            .O(n22_adj_4985));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i8_4_lut_adj_1651.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_unary_minus_2_add_3_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4945), .I3(n32326), .O(n9_adj_4403)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_14 (.CI(n31285), .I0(n2247), .I1(VCC_net), 
            .CO(n31286));
    SB_CARRY rem_4_add_1921_16 (.CI(n31012), .I0(n2844), .I1(VCC_net), 
            .CO(n31013));
    SB_LUT4 i12_4_lut_adj_1652 (.I0(n2143), .I1(n24_adj_4984), .I2(n18_adj_4986), 
            .I3(n2145), .O(n26_adj_4983));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i12_4_lut_adj_1652.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1653 (.I0(n2153), .I1(n26_adj_4983), .I2(n22_adj_4985), 
            .I3(n2151), .O(n2174_adj_4597));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i13_4_lut_adj_1653.LUT_INIT = 16'hfffe;
    SB_LUT4 div_36_LessThan_1606_i39_2_lut (.I0(n2451), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4805));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i1396_3_lut (.I0(n2051), .I1(n2118), .I2(n2075_adj_4609), 
            .I3(GND_net), .O(n2150));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1463_3_lut (.I0(n2150), .I1(n2217), .I2(n2174_adj_4597), 
            .I3(GND_net), .O(n2249));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1466_rep_28_3_lut (.I0(n2153), .I1(n2220), .I2(n2174_adj_4597), 
            .I3(GND_net), .O(n2252));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1466_rep_28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1606_i37_2_lut (.I0(n2452), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4803));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i1467_rep_26_3_lut (.I0(n2154), .I1(n2221), .I2(n2174_adj_4597), 
            .I3(GND_net), .O(n2253));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1467_rep_26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1462_3_lut (.I0(n2149), .I1(n2216), .I2(n2174_adj_4597), 
            .I3(GND_net), .O(n2248));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1654 (.I0(n2256), .I1(n2257), .I2(n2258), .I3(GND_net), 
            .O(n38371));
    defparam i1_3_lut_adj_1654.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_add_1921_15_lut (.I0(GND_net), .I1(n2845), .I2(VCC_net), 
            .I3(n31011), .O(n2912)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_15 (.CI(n31011), .I0(n2845), .I1(VCC_net), 
            .CO(n31012));
    SB_LUT4 i11_4_lut_adj_1655 (.I0(n2248), .I1(n2253), .I2(n2252), .I3(n2249), 
            .O(n26_adj_4924));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i11_4_lut_adj_1655.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut_adj_1656 (.I0(n2246), .I1(n2254), .I2(n38371), .I3(n2255), 
            .O(n19_adj_4926));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i4_4_lut_adj_1656.LUT_INIT = 16'heaaa;
    SB_LUT4 div_36_LessThan_1606_i43_2_lut (.I0(n2449), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4807));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1606_i41_2_lut (.I0(n2450), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4806));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1657 (.I0(n2241), .I1(n2240), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4927));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i1_2_lut_adj_1657.LUT_INIT = 16'heeee;
    SB_LUT4 rem_4_add_1921_14_lut (.I0(GND_net), .I1(n2846), .I2(VCC_net), 
            .I3(n31010), .O(n2913)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9_4_lut_adj_1658 (.I0(n2242), .I1(n2244), .I2(n2243), .I3(n2245), 
            .O(n24_adj_4925));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i9_4_lut_adj_1658.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_1519_13_lut (.I0(GND_net), .I1(n2248), .I2(VCC_net), 
            .I3(n31284), .O(n2315)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13_4_lut_adj_1659 (.I0(n19_adj_4926), .I1(n26_adj_4924), .I2(n2247), 
            .I3(n2250), .O(n28_adj_4923));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i13_4_lut_adj_1659.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1921_14 (.CI(n31010), .I0(n2846), .I1(VCC_net), 
            .CO(n31011));
    SB_CARRY rem_4_unary_minus_2_add_3_26 (.CI(n32326), .I0(GND_net), .I1(n9_adj_4945), 
            .CO(n32327));
    SB_LUT4 i14_4_lut_adj_1660 (.I0(n2251), .I1(n28_adj_4923), .I2(n24_adj_4925), 
            .I3(n16_adj_4927), .O(n2273_adj_4591));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i14_4_lut_adj_1660.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i14_3_lut (.I0(communication_counter[13]), .I1(n20_adj_4392), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2258));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1606_i25_2_lut (.I0(n2458), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4797));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1921_13_lut (.I0(GND_net), .I1(n2847), .I2(VCC_net), 
            .I3(n31009), .O(n2914)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i992_3_lut (.I0(n1455), .I1(n1522), .I2(n1481), .I3(GND_net), 
            .O(n1554_adj_4494));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1539_3_lut (.I0(n2258), .I1(n2325), .I2(n2273_adj_4591), 
            .I3(GND_net), .O(n2357_adj_4589));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1537_3_lut (.I0(n2256), .I1(n2323), .I2(n2273_adj_4591), 
            .I3(GND_net), .O(n2355));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1606_i27_2_lut (.I0(n2457), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4798));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1606_i29_2_lut (.I0(n2456), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4799));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i1536_3_lut (.I0(n2255), .I1(n2322), .I2(n2273_adj_4591), 
            .I3(GND_net), .O(n2354));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_mux_3_i5_3_lut (.I0(encoder0_position[4]), .I1(n21), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n387));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13990_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n14536), .I3(GND_net), .O(n19022));   // verilog/coms.v(126[12] 289[6])
    defparam i13990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1661 (.I0(n2356), .I1(n2358_adj_4588), .I2(GND_net), 
            .I3(GND_net), .O(n40433));
    defparam i1_2_lut_adj_1661.LUT_INIT = 16'heeee;
    SB_CARRY rem_4_add_1519_13 (.CI(n31284), .I0(n2248), .I1(VCC_net), 
            .CO(n31285));
    SB_LUT4 rem_4_add_1519_12_lut (.I0(GND_net), .I1(n2249), .I2(VCC_net), 
            .I3(n31283), .O(n2316)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_12 (.CI(n31283), .I0(n2249), .I1(VCC_net), 
            .CO(n31284));
    SB_CARRY rem_4_add_1921_13 (.CI(n31009), .I0(n2847), .I1(VCC_net), 
            .CO(n31010));
    SB_LUT4 i1_4_lut_adj_1662 (.I0(n2354), .I1(n40433), .I2(n2355), .I3(n2357_adj_4589), 
            .O(n38308));
    defparam i1_4_lut_adj_1662.LUT_INIT = 16'ha080;
    SB_LUT4 i12_4_lut_adj_1663 (.I0(n2353), .I1(n2350), .I2(n2352), .I3(n2348), 
            .O(n28_adj_4999));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i12_4_lut_adj_1663.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1664 (.I0(n2343), .I1(n2345), .I2(n2344), .I3(n38308), 
            .O(n26_adj_5001));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i10_4_lut_adj_1664.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1665 (.I0(n2346), .I1(n2349), .I2(n2351), .I3(n2347), 
            .O(n27_adj_5000));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i11_4_lut_adj_1665.LUT_INIT = 16'hfffe;
    SB_LUT4 div_36_LessThan_1606_i31_2_lut (.I0(n2455), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4800));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1606_i33_2_lut (.I0(n2454), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4801));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1921_12_lut (.I0(GND_net), .I1(n2848), .I2(VCC_net), 
            .I3(n31008), .O(n2915)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9_4_lut_adj_1666 (.I0(n2340), .I1(n2341), .I2(n2339), .I3(n2342), 
            .O(n25_adj_5002));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i9_4_lut_adj_1666.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1667 (.I0(n25_adj_5002), .I1(n27_adj_5000), .I2(n26_adj_5001), 
            .I3(n28_adj_4999), .O(n2372_adj_4587));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i15_4_lut_adj_1667.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i13_3_lut (.I0(communication_counter[12]), .I1(n21_adj_4391), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2358_adj_4588));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1607_3_lut (.I0(n2358_adj_4588), .I1(n2425), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2457_adj_4576));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_add_3_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4946), .I3(n32325), .O(n10_adj_4402)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_25 (.CI(n32325), .I0(GND_net), .I1(n10_adj_4946), 
            .CO(n32326));
    SB_LUT4 rem_4_unary_minus_2_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4947), .I3(n32324), .O(n11_adj_4401)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_24 (.CI(n32324), .I0(GND_net), .I1(n11_adj_4947), 
            .CO(n32325));
    SB_LUT4 rem_4_i1605_3_lut (.I0(n2356), .I1(n2423), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2455_adj_4578));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1605_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_12 (.CI(n31008), .I0(n2848), .I1(VCC_net), 
            .CO(n31009));
    SB_LUT4 rem_4_add_1921_11_lut (.I0(GND_net), .I1(n2849), .I2(VCC_net), 
            .I3(n31007), .O(n2916)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1604_3_lut (.I0(n2355), .I1(n2422), .I2(n2372_adj_4587), 
            .I3(GND_net), .O(n2454_adj_4579));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1668 (.I0(n2439), .I1(n2438), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4914));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i1_2_lut_adj_1668.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1669 (.I0(n2456_adj_4577), .I1(n2458_adj_4575), 
            .I2(GND_net), .I3(GND_net), .O(n40689));
    defparam i1_2_lut_adj_1669.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1670 (.I0(n2454_adj_4579), .I1(n40689), .I2(n2455_adj_4578), 
            .I3(n2457_adj_4576), .O(n38376));
    defparam i1_4_lut_adj_1670.LUT_INIT = 16'ha080;
    SB_LUT4 div_36_LessThan_1606_i19_2_lut (.I0(n2461), .I1(n95_adj_4360), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4792));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_unary_minus_2_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4948), .I3(n32323), .O(n12_adj_4400)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_23 (.CI(n32323), .I0(GND_net), .I1(n12_adj_4948), 
            .CO(n32324));
    SB_CARRY rem_4_add_1921_11 (.CI(n31007), .I0(n2849), .I1(VCC_net), 
            .CO(n31008));
    SB_LUT4 rem_4_add_1921_10_lut (.I0(GND_net), .I1(n2850), .I2(VCC_net), 
            .I3(n31006), .O(n2917)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13_4_lut_adj_1671 (.I0(n2449_adj_4584), .I1(n2451_adj_4582), 
            .I2(n2448_adj_4585), .I3(n18_adj_4914), .O(n30_adj_4908));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i13_4_lut_adj_1671.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1672 (.I0(n2444), .I1(n38376), .I2(n2445), .I3(n2446), 
            .O(n28_adj_4912));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i11_4_lut_adj_1672.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1673 (.I0(n2453_adj_4580), .I1(n2447_adj_4586), 
            .I2(n2452_adj_4581), .I3(n2450_adj_4583), .O(n29_adj_4909));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i12_4_lut_adj_1673.LUT_INIT = 16'hfffe;
    SB_LUT4 div_36_LessThan_1606_i21_2_lut (.I0(n2460), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4794));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 displacement_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4428));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut_adj_1674 (.I0(n2440), .I1(n2442), .I2(n2441), .I3(n2443), 
            .O(n27_adj_4913));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i10_4_lut_adj_1674.LUT_INIT = 16'hfffe;
    SB_LUT4 div_36_LessThan_1606_i23_2_lut (.I0(n2459), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4795));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13991_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n14536), .I3(GND_net), .O(n19023));   // verilog/coms.v(126[12] 289[6])
    defparam i13991_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_10 (.CI(n31006), .I0(n2850), .I1(VCC_net), 
            .CO(n31007));
    SB_LUT4 i16_4_lut_adj_1675 (.I0(n27_adj_4913), .I1(n29_adj_4909), .I2(n28_adj_4912), 
            .I3(n30_adj_4908), .O(n2471_adj_4574));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i16_4_lut_adj_1675.LUT_INIT = 16'hfffe;
    SB_LUT4 div_36_LessThan_1606_i35_2_lut (.I0(n2453), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4802));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i14078_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n14536), 
            .I3(GND_net), .O(n19110));   // verilog/coms.v(126[12] 289[6])
    defparam i14078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1921_9_lut (.I0(GND_net), .I1(n2851), .I2(VCC_net), 
            .I3(n31005), .O(n2918)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14079_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n14536), 
            .I3(GND_net), .O(n19111));   // verilog/coms.v(126[12] 289[6])
    defparam i14079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14080_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n14536), 
            .I3(GND_net), .O(n19112));   // verilog/coms.v(126[12] 289[6])
    defparam i14080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14081_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n14536), 
            .I3(GND_net), .O(n19113));   // verilog/coms.v(126[12] 289[6])
    defparam i14081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4949), .I3(n32322), .O(n13_adj_4399)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_1606_i15_2_lut (.I0(n2463), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4788));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1606_i17_2_lut (.I0(n2462), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4790));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1519_11_lut (.I0(GND_net), .I1(n2250), .I2(VCC_net), 
            .I3(n31282), .O(n2317)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_9 (.CI(n31005), .I0(n2851), .I1(VCC_net), 
            .CO(n31006));
    SB_CARRY rem_4_unary_minus_2_add_3_22 (.CI(n32322), .I0(GND_net), .I1(n13_adj_4949), 
            .CO(n32323));
    SB_LUT4 rem_4_add_1921_8_lut (.I0(GND_net), .I1(n2852), .I2(VCC_net), 
            .I3(n31004), .O(n2919)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i1608_1_lut (.I0(n2471), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2472));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1608_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1921_8 (.CI(n31004), .I0(n2852), .I1(VCC_net), 
            .CO(n31005));
    SB_LUT4 i14082_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n14536), 
            .I3(GND_net), .O(n19114));   // verilog/coms.v(126[12] 289[6])
    defparam i14082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14083_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n14536), 
            .I3(GND_net), .O(n19115));   // verilog/coms.v(126[12] 289[6])
    defparam i14083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14084_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n14536), 
            .I3(GND_net), .O(n19116));   // verilog/coms.v(126[12] 289[6])
    defparam i14084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14085_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n14536), 
            .I3(GND_net), .O(n19117));   // verilog/coms.v(126[12] 289[6])
    defparam i14085_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14086_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n14536), 
            .I3(GND_net), .O(n19118));   // verilog/coms.v(126[12] 289[6])
    defparam i14086_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1519_11 (.CI(n31282), .I0(n2250), .I1(VCC_net), 
            .CO(n31283));
    SB_LUT4 i36165_4_lut (.I0(n35_adj_4802), .I1(n23_adj_4795), .I2(n21_adj_4794), 
            .I3(n19_adj_4792), .O(n43289));
    defparam i36165_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i14087_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n14536), 
            .I3(GND_net), .O(n19119));   // verilog/coms.v(126[12] 289[6])
    defparam i14087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1921_7_lut (.I0(GND_net), .I1(n2853), .I2(VCC_net), 
            .I3(n31003), .O(n2920)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14088_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n14536), 
            .I3(GND_net), .O(n19120));   // verilog/coms.v(126[12] 289[6])
    defparam i14088_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14089_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n14536), 
            .I3(GND_net), .O(n19121));   // verilog/coms.v(126[12] 289[6])
    defparam i14089_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36914_4_lut (.I0(n17_adj_4790), .I1(n15_adj_4788), .I2(n2464), 
            .I3(n98), .O(n44039));
    defparam i36914_4_lut.LUT_INIT = 16'hfeef;
    SB_CARRY rem_4_add_1921_7 (.CI(n31003), .I0(n2853), .I1(VCC_net), 
            .CO(n31004));
    SB_LUT4 i14090_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n14536), .I3(GND_net), .O(n19122));   // verilog/coms.v(126[12] 289[6])
    defparam i14090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14091_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n14536), .I3(GND_net), .O(n19123));   // verilog/coms.v(126[12] 289[6])
    defparam i14091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4371));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14092_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n14536), .I3(GND_net), .O(n19124));   // verilog/coms.v(126[12] 289[6])
    defparam i14092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37296_4_lut (.I0(n23_adj_4795), .I1(n21_adj_4794), .I2(n19_adj_4792), 
            .I3(n44039), .O(n44421));
    defparam i37296_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i37292_4_lut (.I0(n29_adj_4799), .I1(n27_adj_4798), .I2(n25_adj_4797), 
            .I3(n44421), .O(n44417));
    defparam i37292_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i36167_4_lut (.I0(n35_adj_4802), .I1(n33_adj_4801), .I2(n31_adj_4800), 
            .I3(n44417), .O(n43291));
    defparam i36167_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i14093_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n14536), .I3(GND_net), .O(n19125));   // verilog/coms.v(126[12] 289[6])
    defparam i14093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14094_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n14536), .I3(GND_net), .O(n19126));   // verilog/coms.v(126[12] 289[6])
    defparam i14094_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1606_i12_4_lut (.I0(n387), .I1(n99), .I2(n2465), 
            .I3(n558), .O(n12_adj_4786));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i12_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i37458_3_lut (.I0(n12_adj_4786), .I1(n87), .I2(n35_adj_4802), 
            .I3(GND_net), .O(n44583));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37458_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_add_1519_10_lut (.I0(GND_net), .I1(n2251), .I2(VCC_net), 
            .I3(n31281), .O(n2318)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_6_lut (.I0(GND_net), .I1(n2854), .I2(GND_net), 
            .I3(n31002), .O(n2921)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13992_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n14536), .I3(GND_net), .O(n19024));   // verilog/coms.v(126[12] 289[6])
    defparam i13992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13993_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n14536), .I3(GND_net), .O(n19025));   // verilog/coms.v(126[12] 289[6])
    defparam i13993_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_6 (.CI(n31002), .I0(n2854), .I1(GND_net), 
            .CO(n31003));
    SB_LUT4 rem_4_add_1921_5_lut (.I0(GND_net), .I1(n2855), .I2(GND_net), 
            .I3(n31001), .O(n2922)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_5 (.CI(n31001), .I0(n2855), .I1(GND_net), 
            .CO(n31002));
    SB_LUT4 i14095_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n14536), .I3(GND_net), .O(n19127));   // verilog/coms.v(126[12] 289[6])
    defparam i14095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1606_i38_3_lut (.I0(n20_adj_4793), .I1(n83), 
            .I2(n43_adj_4807), .I3(GND_net), .O(n38_adj_4804));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37459_3_lut (.I0(n44583), .I1(n86), .I2(n37_adj_4803), .I3(GND_net), 
            .O(n44584));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37459_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36153_4_lut (.I0(n41_adj_4806), .I1(n39_adj_4805), .I2(n37_adj_4803), 
            .I3(n43289), .O(n43277));
    defparam i36153_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 displacement_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4427));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_1921_4_lut (.I0(GND_net), .I1(n2856), .I2(VCC_net), 
            .I3(n31000), .O(n2923)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37703_4_lut (.I0(n38_adj_4804), .I1(n18_adj_4791), .I2(n43_adj_4807), 
            .I3(n43260), .O(n44828));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37703_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36861_3_lut (.I0(n44584), .I1(n85), .I2(n39_adj_4805), .I3(GND_net), 
            .O(n43986));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36861_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i14096_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n14536), .I3(GND_net), .O(n19128));   // verilog/coms.v(126[12] 289[6])
    defparam i14096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1606_i24_3_lut (.I0(n16_adj_4789), .I1(n91), 
            .I2(n27_adj_4798), .I3(GND_net), .O(n24_adj_4796));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37783_4_lut (.I0(n24_adj_4796), .I1(n14_adj_4787), .I2(n27_adj_4798), 
            .I3(n43307), .O(n44908));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37783_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY rem_4_add_1921_4 (.CI(n31000), .I0(n2856), .I1(VCC_net), 
            .CO(n31001));
    SB_LUT4 rem_4_add_1921_3_lut (.I0(GND_net), .I1(n2857_adj_4442), .I2(VCC_net), 
            .I3(n30999), .O(n2924)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14097_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n14536), .I3(GND_net), .O(n19129));   // verilog/coms.v(126[12] 289[6])
    defparam i14097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37784_3_lut (.I0(n44908), .I1(n90), .I2(n29_adj_4799), .I3(GND_net), 
            .O(n44909));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37784_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_1519_10 (.CI(n31281), .I0(n2251), .I1(VCC_net), 
            .CO(n31282));
    SB_CARRY rem_4_add_1921_3 (.CI(n30999), .I0(n2857_adj_4442), .I1(VCC_net), 
            .CO(n31000));
    SB_LUT4 i37678_3_lut (.I0(n44909), .I1(n89), .I2(n31_adj_4800), .I3(GND_net), 
            .O(n44803));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37678_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_add_1921_2_lut (.I0(GND_net), .I1(n2858), .I2(GND_net), 
            .I3(VCC_net), .O(n2925)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37581_4_lut (.I0(n41_adj_4806), .I1(n39_adj_4805), .I2(n37_adj_4803), 
            .I3(n43291), .O(n44706));
    defparam i37581_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1921_2 (.CI(VCC_net), .I0(n2858), .I1(GND_net), 
            .CO(n30999));
    SB_LUT4 rem_4_add_1988_27_lut (.I0(n2966), .I1(n2933), .I2(VCC_net), 
            .I3(n30998), .O(n3032)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1988_26_lut (.I0(GND_net), .I1(n2934), .I2(VCC_net), 
            .I3(n30997), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_9_lut (.I0(GND_net), .I1(n2252), .I2(VCC_net), 
            .I3(n31280), .O(n2319)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_26 (.CI(n30997), .I0(n2934), .I1(VCC_net), 
            .CO(n30998));
    SB_LUT4 i14098_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n14536), .I3(GND_net), .O(n19130));   // verilog/coms.v(126[12] 289[6])
    defparam i14098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14099_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n14536), .I3(GND_net), .O(n19131));   // verilog/coms.v(126[12] 289[6])
    defparam i14099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37901_4_lut (.I0(n43986), .I1(n44828), .I2(n43_adj_4807), 
            .I3(n43277), .O(n45026));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37901_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36859_3_lut (.I0(n44803), .I1(n88), .I2(n33_adj_4801), .I3(GND_net), 
            .O(n43984));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36859_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37993_4_lut (.I0(n43984), .I1(n45026), .I2(n43_adj_4807), 
            .I3(n44706), .O(n45118));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37993_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i37994_3_lut (.I0(n45118), .I1(n82), .I2(n2448), .I3(GND_net), 
            .O(n45119));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37994_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 rem_4_add_1988_25_lut (.I0(GND_net), .I1(n2935), .I2(VCC_net), 
            .I3(n30996), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14100_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n14536), .I3(GND_net), .O(n19132));   // verilog/coms.v(126[12] 289[6])
    defparam i14100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14101_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n14536), .I3(GND_net), .O(n19133));   // verilog/coms.v(126[12] 289[6])
    defparam i14101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14102_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n14536), .I3(GND_net), .O(n19134));   // verilog/coms.v(126[12] 289[6])
    defparam i14102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1676 (.I0(n45119), .I1(n17236), .I2(n81), .I3(n2447), 
            .O(n2471));
    defparam i1_4_lut_adj_1676.LUT_INIT = 16'hceef;
    SB_CARRY rem_4_add_1988_25 (.CI(n30996), .I0(n2935), .I1(VCC_net), 
            .CO(n30997));
    SB_LUT4 i14103_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n14536), .I3(GND_net), .O(n19135));   // verilog/coms.v(126[12] 289[6])
    defparam i14103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14104_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n14536), .I3(GND_net), .O(n19136));   // verilog/coms.v(126[12] 289[6])
    defparam i14104_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14105_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n14536), .I3(GND_net), .O(n19137));   // verilog/coms.v(126[12] 289[6])
    defparam i14105_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1988_24_lut (.I0(GND_net), .I1(n2936), .I2(VCC_net), 
            .I3(n30995), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14106_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n14536), .I3(GND_net), .O(n19138));   // verilog/coms.v(126[12] 289[6])
    defparam i14106_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14107_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n14536), .I3(GND_net), .O(n19139));   // verilog/coms.v(126[12] 289[6])
    defparam i14107_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14108_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n14536), .I3(GND_net), .O(n19140));   // verilog/coms.v(126[12] 289[6])
    defparam i14108_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14109_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n14536), .I3(GND_net), .O(n19141));   // verilog/coms.v(126[12] 289[6])
    defparam i14109_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14110_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n14536), .I3(GND_net), .O(n19142));   // verilog/coms.v(126[12] 289[6])
    defparam i14110_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1988_24 (.CI(n30995), .I0(n2936), .I1(VCC_net), 
            .CO(n30996));
    SB_LUT4 i14111_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n14536), .I3(GND_net), .O(n19143));   // verilog/coms.v(126[12] 289[6])
    defparam i14111_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14112_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n14536), .I3(GND_net), .O(n19144));   // verilog/coms.v(126[12] 289[6])
    defparam i14112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14113_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n14536), .I3(GND_net), .O(n19145));   // verilog/coms.v(126[12] 289[6])
    defparam i14113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1988_23_lut (.I0(GND_net), .I1(n2937), .I2(VCC_net), 
            .I3(n30994), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4950), .I3(n32321), .O(n14_adj_4398)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_9 (.CI(n31280), .I0(n2252), .I1(VCC_net), 
            .CO(n31281));
    SB_CARRY rem_4_add_1988_23 (.CI(n30994), .I0(n2937), .I1(VCC_net), 
            .CO(n30995));
    SB_LUT4 rem_4_add_1988_22_lut (.I0(GND_net), .I1(n2938), .I2(VCC_net), 
            .I3(n30993), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_22 (.CI(n30993), .I0(n2938), .I1(VCC_net), 
            .CO(n30994));
    SB_LUT4 div_36_LessThan_1545_i41_2_lut (.I0(n2360), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4778));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1545_i45_2_lut (.I0(n2358), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4780));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1545_i39_2_lut (.I0(n2361), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4776));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_mux_3_i6_3_lut (.I0(encoder0_position[5]), .I1(n20_adj_4342), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n386));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1545_i43_2_lut (.I0(n2359), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4779));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1988_21_lut (.I0(GND_net), .I1(n2939), .I2(VCC_net), 
            .I3(n30992), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_1545_i33_2_lut (.I0(n2364), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4773));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i33_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_unary_minus_2_add_3_21 (.CI(n32321), .I0(GND_net), .I1(n14_adj_4950), 
            .CO(n32322));
    SB_LUT4 rem_4_add_1519_8_lut (.I0(GND_net), .I1(n2253), .I2(VCC_net), 
            .I3(n31279), .O(n2320)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_21 (.CI(n30992), .I0(n2939), .I1(VCC_net), 
            .CO(n30993));
    SB_CARRY rem_4_add_1519_8 (.CI(n31279), .I0(n2253), .I1(VCC_net), 
            .CO(n31280));
    SB_LUT4 rem_4_unary_minus_2_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4951), .I3(n32320), .O(n15_adj_4397)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_20 (.CI(n32320), .I0(GND_net), .I1(n15_adj_4951), 
            .CO(n32321));
    SB_LUT4 rem_4_add_1988_20_lut (.I0(GND_net), .I1(n2940), .I2(VCC_net), 
            .I3(n30991), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_20 (.CI(n30991), .I0(n2940), .I1(VCC_net), 
            .CO(n30992));
    SB_LUT4 rem_4_unary_minus_2_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4952), .I3(n32319), .O(n16_adj_4396)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_1545_i35_2_lut (.I0(n2363), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4774));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1545_i17_2_lut (.I0(n2372), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4761));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1545_i19_2_lut (.I0(n2371), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4763));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1519_7_lut (.I0(GND_net), .I1(n2254), .I2(GND_net), 
            .I3(n31278), .O(n2321)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_19 (.CI(n32319), .I0(GND_net), .I1(n16_adj_4952), 
            .CO(n32320));
    SB_LUT4 rem_4_add_1988_19_lut (.I0(GND_net), .I1(n2941), .I2(VCC_net), 
            .I3(n30990), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_19 (.CI(n30990), .I0(n2941), .I1(VCC_net), 
            .CO(n30991));
    SB_CARRY rem_4_add_1519_7 (.CI(n31278), .I0(n2254), .I1(GND_net), 
            .CO(n31279));
    SB_LUT4 rem_4_add_1988_18_lut (.I0(GND_net), .I1(n2942), .I2(VCC_net), 
            .I3(n30989), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_6_lut (.I0(GND_net), .I1(n2255), .I2(GND_net), 
            .I3(n31277), .O(n2322)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_18 (.CI(n30989), .I0(n2942), .I1(VCC_net), 
            .CO(n30990));
    SB_CARRY rem_4_add_1519_6 (.CI(n31277), .I0(n2255), .I1(GND_net), 
            .CO(n31278));
    SB_LUT4 rem_4_add_1519_5_lut (.I0(GND_net), .I1(n2256), .I2(VCC_net), 
            .I3(n31276), .O(n2323)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_1545_i21_2_lut (.I0(n2370), .I1(n95_adj_4360), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4765));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_unary_minus_2_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4953), .I3(n32318), .O(n17_adj_4395)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_1545_i23_2_lut (.I0(n2369), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4767));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i23_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1519_5 (.CI(n31276), .I0(n2256), .I1(VCC_net), 
            .CO(n31277));
    SB_CARRY rem_4_unary_minus_2_add_3_18 (.CI(n32318), .I0(GND_net), .I1(n17_adj_4953), 
            .CO(n32319));
    SB_LUT4 div_36_LessThan_1545_i25_2_lut (.I0(n2368), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4768));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1519_4_lut (.I0(GND_net), .I1(n2257), .I2(VCC_net), 
            .I3(n31275), .O(n2324)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_17_lut (.I0(GND_net), .I1(n2943), .I2(VCC_net), 
            .I3(n30988), .O(n3010)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_4 (.CI(n31275), .I0(n2257), .I1(VCC_net), 
            .CO(n31276));
    SB_LUT4 div_36_LessThan_1545_i37_2_lut (.I0(n2362), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4775));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i37_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1988_17 (.CI(n30988), .I0(n2943), .I1(VCC_net), 
            .CO(n30989));
    SB_LUT4 rem_4_unary_minus_2_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4954), .I3(n32317), .O(n18_adj_4394)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_3_lut (.I0(GND_net), .I1(n2258), .I2(GND_net), 
            .I3(n31274), .O(n2325)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_17 (.CI(n32317), .I0(GND_net), .I1(n18_adj_4954), 
            .CO(n32318));
    SB_LUT4 div_36_LessThan_1545_i27_2_lut (.I0(n2367), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4770));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_unary_minus_2_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4955), .I3(n32316), .O(n19_adj_4393)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_3 (.CI(n31274), .I0(n2258), .I1(GND_net), 
            .CO(n31275));
    SB_CARRY rem_4_add_1519_2 (.CI(VCC_net), .I0(n2358_adj_4588), .I1(VCC_net), 
            .CO(n31274));
    SB_LUT4 rem_4_add_1988_16_lut (.I0(GND_net), .I1(n2944), .I2(VCC_net), 
            .I3(n30987), .O(n3011)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_16 (.CI(n32316), .I0(GND_net), .I1(n19_adj_4955), 
            .CO(n32317));
    SB_LUT4 div_36_unary_minus_2_add_3_25_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(n2_adj_4545), .I3(n31273), .O(n224)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_1988_16 (.CI(n30987), .I0(n2944), .I1(VCC_net), 
            .CO(n30988));
    SB_LUT4 rem_4_unary_minus_2_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4956), .I3(n32315), .O(n20_adj_4392)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_unary_minus_2_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4546), .I3(n31272), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_15 (.CI(n32315), .I0(GND_net), .I1(n20_adj_4956), 
            .CO(n32316));
    SB_LUT4 div_36_LessThan_1545_i29_2_lut (.I0(n2366), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4771));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1545_i31_2_lut (.I0(n2365), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4772));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_i1547_1_lut (.I0(n2381), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2382));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1547_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13994_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position[16]), 
            .I2(n14536), .I3(GND_net), .O(n19026));   // verilog/coms.v(126[12] 289[6])
    defparam i13994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36259_4_lut (.I0(n37_adj_4775), .I1(n25_adj_4768), .I2(n23_adj_4767), 
            .I3(n21_adj_4765), .O(n43384));
    defparam i36259_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36966_4_lut (.I0(n19_adj_4763), .I1(n17_adj_4761), .I2(n2373), 
            .I3(n98), .O(n44091));
    defparam i36966_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 rem_4_add_1988_15_lut (.I0(GND_net), .I1(n2945), .I2(VCC_net), 
            .I3(n30986), .O(n3012)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_2_add_3_24 (.CI(n31272), .I0(GND_net), .I1(n3_adj_4546), 
            .CO(n31273));
    SB_LUT4 i37322_4_lut (.I0(n25_adj_4768), .I1(n23_adj_4767), .I2(n21_adj_4765), 
            .I3(n44091), .O(n44447));
    defparam i37322_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i37320_4_lut (.I0(n31_adj_4772), .I1(n29_adj_4771), .I2(n27_adj_4770), 
            .I3(n44447), .O(n44445));
    defparam i37320_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 rem_4_unary_minus_2_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4957), .I3(n32314), .O(n21_adj_4391)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_15 (.CI(n30986), .I0(n2945), .I1(VCC_net), 
            .CO(n30987));
    SB_LUT4 i36265_4_lut (.I0(n37_adj_4775), .I1(n35_adj_4774), .I2(n33_adj_4773), 
            .I3(n44445), .O(n43390));
    defparam i36265_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY rem_4_unary_minus_2_add_3_14 (.CI(n32314), .I0(GND_net), .I1(n21_adj_4957), 
            .CO(n32315));
    SB_LUT4 rem_4_add_1988_14_lut (.I0(GND_net), .I1(n2946), .I2(VCC_net), 
            .I3(n30985), .O(n3013)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_unary_minus_2_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4547), .I3(n31271), .O(n4_adj_4326)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4958), .I3(n32313), .O(n22_adj_4390)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_2_add_3_23 (.CI(n31271), .I0(GND_net), .I1(n4_adj_4547), 
            .CO(n31272));
    SB_LUT4 div_36_LessThan_1545_i14_4_lut (.I0(n386), .I1(n99), .I2(n2374), 
            .I3(n558), .O(n14_adj_4759));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i14_4_lut.LUT_INIT = 16'h0317;
    SB_IO PIN_22_pad (.PACKAGE_PIN(PIN_22), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_22_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_22_pad.PIN_TYPE = 6'b011001;
    defparam PIN_22_pad.PULLUP = 1'b0;
    defparam PIN_22_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i37462_3_lut (.I0(n14_adj_4759), .I1(n87), .I2(n37_adj_4775), 
            .I3(GND_net), .O(n44587));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37462_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37463_3_lut (.I0(n44587), .I1(n86), .I2(n39_adj_4776), .I3(GND_net), 
            .O(n44588));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37463_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 displacement_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4426));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_unary_minus_2_add_3_13 (.CI(n32313), .I0(GND_net), .I1(n22_adj_4958), 
            .CO(n32314));
    SB_LUT4 div_36_unary_minus_2_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4548), .I3(n31270), .O(n5_adj_4358)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_14 (.CI(n30985), .I0(n2946), .I1(VCC_net), 
            .CO(n30986));
    SB_LUT4 rem_4_unary_minus_2_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4959), .I3(n32312), .O(n23_adj_4389)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_1545_i40_3_lut (.I0(n22_adj_4766), .I1(n83), 
            .I2(n45_adj_4780), .I3(GND_net), .O(n40_adj_4777));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY div_36_unary_minus_2_add_3_22 (.CI(n31270), .I0(GND_net), .I1(n5_adj_4548), 
            .CO(n31271));
    SB_LUT4 i14325_3_lut (.I0(encoder0_position[3]), .I1(n2886), .I2(count_enable), 
            .I3(GND_net), .O(n19357));   // quad.v(35[10] 41[6])
    defparam i14325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_unary_minus_2_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4549), .I3(n31269), .O(n6_adj_4431)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_12 (.CI(n32312), .I0(GND_net), .I1(n23_adj_4959), 
            .CO(n32313));
    SB_LUT4 i14324_3_lut (.I0(encoder0_position[2]), .I1(n2887), .I2(count_enable), 
            .I3(GND_net), .O(n19356));   // quad.v(35[10] 41[6])
    defparam i14324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36210_4_lut (.I0(n43_adj_4779), .I1(n41_adj_4778), .I2(n39_adj_4776), 
            .I3(n43384), .O(n43334));
    defparam i36210_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37553_4_lut (.I0(n40_adj_4777), .I1(n20_adj_4764), .I2(n45_adj_4780), 
            .I3(n43327), .O(n44678));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37553_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 rem_4_unary_minus_2_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4960), .I3(n32311), .O(n24_adj_4386)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36855_3_lut (.I0(n44588), .I1(n85), .I2(n41_adj_4778), .I3(GND_net), 
            .O(n43980));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36855_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_unary_minus_2_add_3_11 (.CI(n32311), .I0(GND_net), .I1(n24_adj_4960), 
            .CO(n32312));
    SB_LUT4 i14323_3_lut (.I0(encoder0_position[1]), .I1(n2888), .I2(count_enable), 
            .I3(GND_net), .O(n19355));   // quad.v(35[10] 41[6])
    defparam i14323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14327_3_lut (.I0(encoder0_position[5]), .I1(n2884), .I2(count_enable), 
            .I3(GND_net), .O(n19359));   // quad.v(35[10] 41[6])
    defparam i14327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14326_3_lut (.I0(encoder0_position[4]), .I1(n2885), .I2(count_enable), 
            .I3(GND_net), .O(n19358));   // quad.v(35[10] 41[6])
    defparam i14326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1545_i26_3_lut (.I0(n18_adj_4762), .I1(n91), 
            .I2(n29_adj_4771), .I3(GND_net), .O(n26_adj_4769));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37775_4_lut (.I0(n26_adj_4769), .I1(n16_adj_4760), .I2(n29_adj_4771), 
            .I3(n43406), .O(n44900));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37775_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i37776_3_lut (.I0(n44900), .I1(n90), .I2(n31_adj_4772), .I3(GND_net), 
            .O(n44901));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37776_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37680_3_lut (.I0(n44901), .I1(n89), .I2(n33_adj_4773), .I3(GND_net), 
            .O(n44805));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37680_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37613_4_lut (.I0(n43_adj_4779), .I1(n41_adj_4778), .I2(n39_adj_4776), 
            .I3(n43390), .O(n44738));
    defparam i37613_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i37877_4_lut (.I0(n43980), .I1(n44678), .I2(n45_adj_4780), 
            .I3(n43334), .O(n45002));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37877_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36853_3_lut (.I0(n44805), .I1(n88), .I2(n35_adj_4774), .I3(GND_net), 
            .O(n43978));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36853_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i14329_3_lut (.I0(encoder0_position[7]), .I1(n2882), .I2(count_enable), 
            .I3(GND_net), .O(n19361));   // quad.v(35[10] 41[6])
    defparam i14329_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37879_4_lut (.I0(n43978), .I1(n45002), .I2(n45_adj_4780), 
            .I3(n44738), .O(n45004));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37879_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14328_3_lut (.I0(encoder0_position[6]), .I1(n2883), .I2(count_enable), 
            .I3(GND_net), .O(n19360));   // quad.v(35[10] 41[6])
    defparam i14328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i991_rep_46_3_lut (.I0(n1454), .I1(n1521), .I2(n1481), 
            .I3(GND_net), .O(n1553_adj_4493));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i991_rep_46_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1677 (.I0(n45004), .I1(n17311), .I2(n82), .I3(n2357), 
            .O(n2381));
    defparam i1_4_lut_adj_1677.LUT_INIT = 16'hceef;
    SB_LUT4 i14331_3_lut (.I0(encoder0_position[9]), .I1(n2880), .I2(count_enable), 
            .I3(GND_net), .O(n19363));   // quad.v(35[10] 41[6])
    defparam i14331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14330_3_lut (.I0(encoder0_position[8]), .I1(n2881), .I2(count_enable), 
            .I3(GND_net), .O(n19362));   // quad.v(35[10] 41[6])
    defparam i14330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1482_i37_2_lut (.I0(n2269), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4755));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i990_3_lut (.I0(n1453), .I1(n1520), .I2(n1481), .I3(GND_net), 
            .O(n1552));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14333_3_lut (.I0(encoder0_position[11]), .I1(n2878), .I2(count_enable), 
            .I3(GND_net), .O(n19365));   // quad.v(35[10] 41[6])
    defparam i14333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1482_i43_2_lut (.I0(n2266), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4758));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i14332_3_lut (.I0(encoder0_position[10]), .I1(n2879), .I2(count_enable), 
            .I3(GND_net), .O(n19364));   // quad.v(35[10] 41[6])
    defparam i14332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1482_i41_2_lut (.I0(n2267), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4757));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1482_i39_2_lut (.I0(n2268), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4756));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_mux_3_i7_3_lut (.I0(encoder0_position[6]), .I1(n19_adj_4343), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n385));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4425));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_1482_i19_2_lut (.I0(n2278), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4743));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1482_i21_2_lut (.I0(n2277), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4745));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i14335_3_lut (.I0(encoder0_position[13]), .I1(n2876), .I2(count_enable), 
            .I3(GND_net), .O(n19367));   // quad.v(35[10] 41[6])
    defparam i14335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14334_3_lut (.I0(encoder0_position[12]), .I1(n2877), .I2(count_enable), 
            .I3(GND_net), .O(n19366));   // quad.v(35[10] 41[6])
    defparam i14334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1482_i31_2_lut (.I0(n2272), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4752));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1482_i33_2_lut (.I0(n2271), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4753));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1482_i35_2_lut (.I0(n2270), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4754));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1482_i23_2_lut (.I0(n2276), .I1(n95_adj_4360), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4747));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1482_i25_2_lut (.I0(n2275), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4748));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1482_i27_2_lut (.I0(n2274), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4749));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1482_i29_2_lut (.I0(n2273), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4751));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_i1484_1_lut (.I0(n2288), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2289));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1484_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_1482_i17_2_lut (.I0(n2279), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4741));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i36390_4_lut (.I0(n23_adj_4747), .I1(n21_adj_4745), .I2(n19_adj_4743), 
            .I3(n17_adj_4741), .O(n43515));
    defparam i36390_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36382_4_lut (.I0(n29_adj_4751), .I1(n27_adj_4749), .I2(n25_adj_4748), 
            .I3(n43515), .O(n43507));
    defparam i36382_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37623_4_lut (.I0(n35_adj_4754), .I1(n33_adj_4753), .I2(n31_adj_4752), 
            .I3(n43507), .O(n44748));
    defparam i37623_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(n10_adj_4350), .I1(one_wire_N_513[11]), .I2(one_wire_N_513[7]), 
            .I3(GND_net), .O(n12_adj_4435));
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_2_lut_adj_1678 (.I0(one_wire_N_513[5]), .I1(n8_adj_4437), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4436));
    defparam i4_2_lut_adj_1678.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1679 (.I0(state[1]), .I1(n11_adj_4436), .I2(start), 
            .I3(n12_adj_4435), .O(n38192));
    defparam i2_4_lut_adj_1679.LUT_INIT = 16'hfffe;
    SB_LUT4 div_36_LessThan_1482_i16_4_lut (.I0(n385), .I1(n99), .I2(n2280), 
            .I3(n558), .O(n16_adj_4740));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i16_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i37468_3_lut (.I0(n16_adj_4740), .I1(n87), .I2(n39_adj_4756), 
            .I3(GND_net), .O(n44593));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37468_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37469_3_lut (.I0(n44593), .I1(n86), .I2(n41_adj_4757), .I3(GND_net), 
            .O(n44594));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37469_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36982_4_lut (.I0(n41_adj_4757), .I1(n39_adj_4756), .I2(n27_adj_4749), 
            .I3(n43509), .O(n44107));
    defparam i36982_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i37551_3_lut (.I0(n22_adj_4746), .I1(n93), .I2(n27_adj_4749), 
            .I3(GND_net), .O(n44676));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37551_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36845_3_lut (.I0(n44594), .I1(n85), .I2(n43_adj_4758), .I3(GND_net), 
            .O(n43970));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36845_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_i855_3_lut (.I0(n1254), .I1(n1321), .I2(n1283), .I3(GND_net), 
            .O(n1353));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i919_3_lut (.I0(n1350), .I1(n1417_adj_4496), .I2(n1382), 
            .I3(GND_net), .O(n1449));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i923_3_lut (.I0(n1354), .I1(n1421), .I2(n1382), .I3(GND_net), 
            .O(n1453));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i854_3_lut (.I0(n1253), .I1(n1320), .I2(n1283), .I3(GND_net), 
            .O(n1352));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1482_i28_3_lut (.I0(n20_adj_4744), .I1(n91), 
            .I2(n31_adj_4752), .I3(GND_net), .O(n28_adj_4750));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37855_4_lut (.I0(n28_adj_4750), .I1(n18_adj_4742), .I2(n31_adj_4752), 
            .I3(n43505), .O(n44980));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37855_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 rem_4_i920_3_lut (.I0(n1351), .I1(n1418_adj_4497), .I2(n1382), 
            .I3(GND_net), .O(n1450));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i921_3_lut (.I0(n1352), .I1(n1419_adj_4498), .I2(n1382), 
            .I3(GND_net), .O(n1451));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i852_3_lut (.I0(n1251), .I1(n1318), .I2(n1283), .I3(GND_net), 
            .O(n1350));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i857_3_lut (.I0(n1256), .I1(n1323), .I2(n1283), .I3(GND_net), 
            .O(n1355));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i856_3_lut (.I0(n1255), .I1(n1322), .I2(n1283), .I3(GND_net), 
            .O(n1354));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i853_3_lut (.I0(n1252), .I1(n1319), .I2(n1283), .I3(GND_net), 
            .O(n1351));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i789_3_lut (.I0(n1156), .I1(n1223), .I2(n1184), .I3(GND_net), 
            .O(n1255));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i788_3_lut (.I0(n1155), .I1(n1222), .I2(n1184), .I3(GND_net), 
            .O(n1254));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i791_3_lut (.I0(n1158), .I1(n1225), .I2(n1184), .I3(GND_net), 
            .O(n1257));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i790_3_lut (.I0(n1157), .I1(n1224), .I2(n1184), .I3(GND_net), 
            .O(n1256));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i718_3_lut (.I0(n1053), .I1(n1120), .I2(n1085), .I3(GND_net), 
            .O(n1152));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i651_3_lut (.I0(n954), .I1(n1021), .I2(n986), .I3(GND_net), 
            .O(n1053));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i653_3_lut (.I0(n956), .I1(n1023), .I2(n986), .I3(GND_net), 
            .O(n1055));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i652_3_lut (.I0(n955), .I1(n1022), .I2(n986), .I3(GND_net), 
            .O(n1054));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37856_3_lut (.I0(n44980), .I1(n90), .I2(n33_adj_4753), .I3(GND_net), 
            .O(n44981));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37856_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37688_3_lut (.I0(n44981), .I1(n89), .I2(n35_adj_4754), .I3(GND_net), 
            .O(n44813));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37688_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36988_4_lut (.I0(n41_adj_4757), .I1(n39_adj_4756), .I2(n37_adj_4755), 
            .I3(n44748), .O(n44113));
    defparam i36988_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i14339_3_lut (.I0(encoder0_position[17]), .I1(n2872), .I2(count_enable), 
            .I3(GND_net), .O(n19371));   // quad.v(35[10] 41[6])
    defparam i14339_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37681_4_lut (.I0(n43970), .I1(n44676), .I2(n43_adj_4758), 
            .I3(n44107), .O(n44806));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37681_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 unary_minus_18_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36843_3_lut (.I0(n44813), .I1(n88), .I2(n37_adj_4755), .I3(GND_net), 
            .O(n43968));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36843_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i14338_3_lut (.I0(encoder0_position[16]), .I1(n2873), .I2(count_enable), 
            .I3(GND_net), .O(n19370));   // quad.v(35[10] 41[6])
    defparam i14338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i28_3_lut (.I0(communication_counter[27]), .I1(n6_adj_4406), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n855));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i29_3_lut (.I0(communication_counter[28]), .I1(n5_adj_4407), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n749));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i31_3_lut (.I0(communication_counter[30]), .I1(n3_adj_4409), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n852));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1680 (.I0(n852), .I1(n749), .I2(n748), .I3(n855), 
            .O(n40223));
    defparam i1_4_lut_adj_1680.LUT_INIT = 16'haaa8;
    SB_LUT4 rem_4_mux_3_i30_3_lut (.I0(communication_counter[29]), .I1(n4_adj_4408), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n748));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i30984_2_lut (.I0(n39906), .I1(n746), .I2(GND_net), .I3(GND_net), 
            .O(n953));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i30984_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_3_lut_adj_1681 (.I0(n956), .I1(n957), .I2(n958), .I3(GND_net), 
            .O(n38251));
    defparam i1_3_lut_adj_1681.LUT_INIT = 16'hfefe;
    SB_LUT4 i22453_4_lut (.I0(n954), .I1(n953), .I2(n38251), .I3(n955), 
            .O(n986));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i22453_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 rem_4_mux_3_i27_3_lut (.I0(communication_counter[26]), .I1(n7_adj_4405), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n958));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i655_3_lut (.I0(n958), .I1(n1025), .I2(n986), .I3(GND_net), 
            .O(n1057));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14337_3_lut (.I0(encoder0_position[15]), .I1(n2874), .I2(count_enable), 
            .I3(GND_net), .O(n19369));   // quad.v(35[10] 41[6])
    defparam i14337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37926_4_lut (.I0(n43968), .I1(n44806), .I2(n43_adj_4758), 
            .I3(n44113), .O(n45051));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37926_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 rem_4_add_1988_13_lut (.I0(GND_net), .I1(n2947), .I2(VCC_net), 
            .I3(n30984), .O(n3014)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37927_3_lut (.I0(n45051), .I1(n84), .I2(n2265), .I3(GND_net), 
            .O(n45052));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37927_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1682 (.I0(n45052), .I1(n17308), .I2(n83), .I3(n2264), 
            .O(n2288));
    defparam i1_4_lut_adj_1682.LUT_INIT = 16'hceef;
    SB_LUT4 i14336_3_lut (.I0(encoder0_position[14]), .I1(n2875), .I2(count_enable), 
            .I3(GND_net), .O(n19368));   // quad.v(35[10] 41[6])
    defparam i14336_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i654_3_lut (.I0(n957), .I1(n1024), .I2(n986), .I3(GND_net), 
            .O(n1056));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1683 (.I0(n1056), .I1(n1057), .I2(n1058), .I3(GND_net), 
            .O(n38249));
    defparam i1_3_lut_adj_1683.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1684 (.I0(n1054), .I1(n1055), .I2(GND_net), .I3(GND_net), 
            .O(n40249));
    defparam i1_2_lut_adj_1684.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1685 (.I0(n1052), .I1(n40249), .I2(n1053), .I3(n38249), 
            .O(n1085));
    defparam i1_4_lut_adj_1685.LUT_INIT = 16'hfefa;
    SB_LUT4 rem_4_mux_3_i26_3_lut (.I0(communication_counter[25]), .I1(n8_adj_4404), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1058));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i723_3_lut (.I0(n1058), .I1(n1125), .I2(n1085), .I3(GND_net), 
            .O(n1157));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i721_3_lut (.I0(n1056), .I1(n1123), .I2(n1085), .I3(GND_net), 
            .O(n1155));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i720_3_lut (.I0(n1055), .I1(n1122), .I2(n1085), .I3(GND_net), 
            .O(n1154));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i25_3_lut (.I0(communication_counter[24]), .I1(n9_adj_4403), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1158));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i722_3_lut (.I0(n1057), .I1(n1124), .I2(n1085), .I3(GND_net), 
            .O(n1156));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1686 (.I0(n1156), .I1(n1158), .I2(GND_net), .I3(GND_net), 
            .O(n40253));
    defparam i1_2_lut_adj_1686.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1687 (.I0(n1154), .I1(n40253), .I2(n1155), .I3(n1157), 
            .O(n38245));
    defparam i1_4_lut_adj_1687.LUT_INIT = 16'ha080;
    SB_LUT4 i3_4_lut_adj_1688 (.I0(n38245), .I1(n1152), .I2(n1151), .I3(n1153), 
            .O(n1184));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i3_4_lut_adj_1688.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i719_3_lut (.I0(n1054), .I1(n1121), .I2(n1085), .I3(GND_net), 
            .O(n1153));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i786_3_lut (.I0(n1153), .I1(n1220), .I2(n1184), .I3(GND_net), 
            .O(n1252));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i787_3_lut (.I0(n1154), .I1(n1221), .I2(n1184), .I3(GND_net), 
            .O(n1253));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1417_i39_2_lut (.I0(n2172), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4734));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1417_i45_2_lut (.I0(n2169), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4737));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i785_3_lut (.I0(n1152), .I1(n1219), .I2(n1184), .I3(GND_net), 
            .O(n1251));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1689 (.I0(n1256), .I1(n1257), .I2(n1258), .I3(GND_net), 
            .O(n38243));
    defparam i1_3_lut_adj_1689.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1690 (.I0(n1254), .I1(n1250), .I2(n38243), .I3(n1255), 
            .O(n6_adj_4922));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i1_4_lut_adj_1690.LUT_INIT = 16'heccc;
    SB_LUT4 i4_4_lut_adj_1691 (.I0(n1251), .I1(n1253), .I2(n1252), .I3(n6_adj_4922), 
            .O(n1283));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i4_4_lut_adj_1691.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i24_3_lut (.I0(communication_counter[23]), .I1(n10_adj_4402), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1258));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i859_3_lut (.I0(n1258), .I1(n1325), .I2(n1283), .I3(GND_net), 
            .O(n1357));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i858_3_lut (.I0(n1257), .I1(n1324), .I2(n1283), .I3(GND_net), 
            .O(n1356));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1692 (.I0(n1356), .I1(n1357), .I2(n1358), .I3(GND_net), 
            .O(n38239));
    defparam i1_3_lut_adj_1692.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut_adj_1693 (.I0(n1351), .I1(n1354), .I2(n38239), .I3(n1355), 
            .O(n8_adj_4917));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i2_4_lut_adj_1693.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_2_lut_adj_1694 (.I0(n1350), .I1(n1349), .I2(GND_net), .I3(GND_net), 
            .O(n7_adj_4918));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i1_2_lut_adj_1694.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut_adj_1695 (.I0(n1352), .I1(n7_adj_4918), .I2(n1353), 
            .I3(n8_adj_4917), .O(n1382));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i5_4_lut_adj_1695.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i23_3_lut (.I0(communication_counter[22]), .I1(n11_adj_4401), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1358));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i927_3_lut (.I0(n1358), .I1(n1425), .I2(n1382), .I3(GND_net), 
            .O(n1457));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i925_3_lut (.I0(n1356), .I1(n1423), .I2(n1382), .I3(GND_net), 
            .O(n1455));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i924_3_lut (.I0(n1355), .I1(n1422), .I2(n1382), .I3(GND_net), 
            .O(n1454));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i22_3_lut (.I0(communication_counter[21]), .I1(n12_adj_4400), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1458));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i926_3_lut (.I0(n1357), .I1(n1424), .I2(n1382), .I3(GND_net), 
            .O(n1456));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1417_i43_2_lut (.I0(n2170), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4736));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1417_i41_2_lut (.I0(n2171), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4735));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_mux_3_i8_3_lut (.I0(encoder0_position[7]), .I1(n18_adj_4344), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n384));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1696 (.I0(n1456), .I1(n1458), .I2(GND_net), .I3(GND_net), 
            .O(n40389));
    defparam i1_2_lut_adj_1696.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1697 (.I0(n1454), .I1(n40389), .I2(n1455), .I3(n1457), 
            .O(n38273));
    defparam i1_4_lut_adj_1697.LUT_INIT = 16'ha080;
    SB_LUT4 i5_4_lut_adj_1698 (.I0(n38273), .I1(n1451), .I2(n1450), .I3(n1452), 
            .O(n12_adj_4590));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i5_4_lut_adj_1698.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1699 (.I0(n1453), .I1(n12_adj_4590), .I2(n1449), 
            .I3(n1448), .O(n1481));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i6_4_lut_adj_1699.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i922_3_lut (.I0(n1353), .I1(n1420_adj_4499), .I2(n1382), 
            .I3(GND_net), .O(n1452));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i989_3_lut (.I0(n1452), .I1(n1519), .I2(n1481), .I3(GND_net), 
            .O(n1551));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1417_i33_2_lut (.I0(n2175), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4731));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1417_i35_2_lut (.I0(n2174), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4732));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 displacement_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4424));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_1417_i37_2_lut (.I0(n2173), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4733));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i1729_3_lut (.I0(n2544_adj_4518), .I1(n2611), .I2(n2570), 
            .I3(GND_net), .O(n2643_adj_4489));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1729_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1417_i29_2_lut (.I0(n2177), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4728));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1417_i31_2_lut (.I0(n2176), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4730));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i1730_3_lut (.I0(n2545_adj_4517), .I1(n2612), .I2(n2570), 
            .I3(GND_net), .O(n2644));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1730_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1417_i27_2_lut (.I0(n2178), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4727));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i1728_3_lut (.I0(n2543_adj_4519), .I1(n2610), .I2(n2570), 
            .I3(GND_net), .O(n2642_adj_4490));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1417_i21_2_lut (.I0(n2181), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4721));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1417_i23_2_lut (.I0(n2180), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4723));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1417_i25_2_lut (.I0(n2179), .I1(n95_adj_4360), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4725));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i1734_3_lut (.I0(n2549_adj_4513), .I1(n2616), .I2(n2570), 
            .I3(GND_net), .O(n2648));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1733_3_lut (.I0(n2548_adj_4514), .I1(n2615), .I2(n2570), 
            .I3(GND_net), .O(n2647));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1419_1_lut (.I0(n2192), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2193));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1419_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_1417_i19_2_lut (.I0(n2182), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4719));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i36454_4_lut (.I0(n25_adj_4725), .I1(n23_adj_4723), .I2(n21_adj_4721), 
            .I3(n19_adj_4719), .O(n43579));
    defparam i36454_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36439_4_lut (.I0(n31_adj_4730), .I1(n29_adj_4728), .I2(n27_adj_4727), 
            .I3(n43579), .O(n43564));
    defparam i36439_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37629_4_lut (.I0(n37_adj_4733), .I1(n35_adj_4732), .I2(n33_adj_4731), 
            .I3(n43564), .O(n44754));
    defparam i37629_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_36_LessThan_1417_i18_4_lut (.I0(n384), .I1(n99), .I2(n2183), 
            .I3(n558), .O(n18_adj_4718));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i18_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i37474_3_lut (.I0(n18_adj_4718), .I1(n87), .I2(n41_adj_4735), 
            .I3(GND_net), .O(n44599));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37474_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_1988_13 (.CI(n30984), .I0(n2947), .I1(VCC_net), 
            .CO(n30985));
    SB_LUT4 i37475_3_lut (.I0(n44599), .I1(n86), .I2(n43_adj_4736), .I3(GND_net), 
            .O(n44600));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37475_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37024_4_lut (.I0(n43_adj_4736), .I1(n41_adj_4735), .I2(n29_adj_4728), 
            .I3(n43577), .O(n44149));
    defparam i37024_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_36_LessThan_1417_i26_3_lut (.I0(n24_adj_4724), .I1(n93), 
            .I2(n29_adj_4728), .I3(GND_net), .O(n26_adj_4726));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i14350_3_lut (.I0(encoder1_position[4]), .I1(n2835), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19382));   // quad.v(35[10] 41[6])
    defparam i14350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36839_3_lut (.I0(n44600), .I1(n85), .I2(n45_adj_4737), .I3(GND_net), 
            .O(n43964));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36839_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i14349_3_lut (.I0(encoder1_position[3]), .I1(n2836), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19381));   // quad.v(35[10] 41[6])
    defparam i14349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14348_3_lut (.I0(encoder1_position[2]), .I1(n2837), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19380));   // quad.v(35[10] 41[6])
    defparam i14348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1736_3_lut (.I0(n2551_adj_4511), .I1(n2618_adj_4507), 
            .I2(n2570), .I3(GND_net), .O(n2650));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1736_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1417_i30_3_lut (.I0(n22_adj_4722), .I1(n91), 
            .I2(n33_adj_4731), .I3(GND_net), .O(n30_adj_4729));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37853_4_lut (.I0(n30_adj_4729), .I1(n20_adj_4720), .I2(n33_adj_4731), 
            .I3(n43562), .O(n44978));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37853_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i14347_3_lut (.I0(encoder1_position[1]), .I1(n2838), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19379));   // quad.v(35[10] 41[6])
    defparam i14347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37854_3_lut (.I0(n44978), .I1(n90), .I2(n35_adj_4732), .I3(GND_net), 
            .O(n44979));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37854_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37698_3_lut (.I0(n44979), .I1(n89), .I2(n37_adj_4733), .I3(GND_net), 
            .O(n44823));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37698_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37026_4_lut (.I0(n43_adj_4736), .I1(n41_adj_4735), .I2(n39_adj_4734), 
            .I3(n44754), .O(n44151));
    defparam i37026_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i37546_4_lut (.I0(n43964), .I1(n26_adj_4726), .I2(n45_adj_4737), 
            .I3(n44149), .O(n44671));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37546_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36837_3_lut (.I0(n44823), .I1(n88), .I2(n39_adj_4734), .I3(GND_net), 
            .O(n43962));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36837_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37548_4_lut (.I0(n43962), .I1(n44671), .I2(n45_adj_4737), 
            .I3(n44151), .O(n44673));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37548_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 rem_4_i1738_3_lut (.I0(n2553_adj_4509), .I1(n2620_adj_4502), 
            .I2(n2570), .I3(GND_net), .O(n2652));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1700 (.I0(n44673), .I1(n17231), .I2(n84), .I3(n2168), 
            .O(n2192));
    defparam i1_4_lut_adj_1700.LUT_INIT = 16'hceef;
    SB_LUT4 div_36_LessThan_1350_i41_2_lut (.I0(n2072), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4716));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1350_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1350_i39_2_lut (.I0(n2073), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4715));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1350_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1988_12_lut (.I0(GND_net), .I1(n2948), .I2(VCC_net), 
            .I3(n30983), .O(n3015)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_1350_i37_2_lut (.I0(n2074), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4714));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1350_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1350_i35_2_lut (.I0(n2075), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4713));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1350_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_mux_3_i9_3_lut (.I0(encoder0_position[8]), .I1(n17_adj_4410), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n383));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1350_i31_2_lut (.I0(n2077), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4710));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1350_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1350_i33_2_lut (.I0(n2076), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4712));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1350_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1350_i29_2_lut (.I0(n2078), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4709));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1350_i29_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY div_36_unary_minus_2_add_3_21 (.CI(n31269), .I0(GND_net), .I1(n6_adj_4549), 
            .CO(n31270));
    SB_LUT4 div_36_unary_minus_2_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4550), .I3(n31268), .O(n7_adj_4432)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4961), .I3(n32310), .O(n25_adj_4385)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_2_add_3_20 (.CI(n31268), .I0(GND_net), .I1(n7_adj_4550), 
            .CO(n31269));
    SB_CARRY rem_4_add_1988_12 (.CI(n30983), .I0(n2948), .I1(VCC_net), 
            .CO(n30984));
    SB_CARRY rem_4_unary_minus_2_add_3_10 (.CI(n32310), .I0(GND_net), .I1(n25_adj_4961), 
            .CO(n32311));
    SB_LUT4 rem_4_unary_minus_2_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n26_adj_4962), .I3(n32309), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_9 (.CI(n32309), .I0(GND_net), .I1(n26_adj_4962), 
            .CO(n32310));
    SB_LUT4 rem_4_add_1988_11_lut (.I0(GND_net), .I1(n2949), .I2(VCC_net), 
            .I3(n30982), .O(n3016)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_1350_i23_2_lut (.I0(n2081), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4703));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1350_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1350_i25_2_lut (.I0(n2080), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4705));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1350_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_unary_minus_2_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4551), .I3(n31267), .O(n8_adj_4369)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_11 (.CI(n30982), .I0(n2949), .I1(VCC_net), 
            .CO(n30983));
    SB_LUT4 div_36_LessThan_1350_i27_2_lut (.I0(n2079), .I1(n95_adj_4360), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4707));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1350_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_unary_minus_2_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n27_adj_4963), .I3(n32308), .O(n27_adj_4381)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_2_add_3_19 (.CI(n31267), .I0(GND_net), .I1(n8_adj_4551), 
            .CO(n31268));
    SB_LUT4 div_36_unary_minus_2_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4552), .I3(n31266), .O(n9_adj_4370)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_10_lut (.I0(GND_net), .I1(n2950), .I2(VCC_net), 
            .I3(n30981), .O(n3017)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_10 (.CI(n30981), .I0(n2950), .I1(VCC_net), 
            .CO(n30982));
    SB_CARRY rem_4_unary_minus_2_add_3_8 (.CI(n32308), .I0(GND_net), .I1(n27_adj_4963), 
            .CO(n32309));
    SB_LUT4 rem_4_unary_minus_2_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n28_adj_4964), .I3(n32307), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_2_add_3_18 (.CI(n31266), .I0(GND_net), .I1(n9_adj_4552), 
            .CO(n31267));
    SB_CARRY rem_4_unary_minus_2_add_3_7 (.CI(n32307), .I0(GND_net), .I1(n28_adj_4964), 
            .CO(n32308));
    SB_LUT4 div_36_i1352_1_lut (.I0(n2093), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2094));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1352_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_1350_i21_2_lut (.I0(n2082), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4701));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1350_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i36506_4_lut (.I0(n27_adj_4707), .I1(n25_adj_4705), .I2(n23_adj_4703), 
            .I3(n21_adj_4701), .O(n43631));
    defparam i36506_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36491_4_lut (.I0(n33_adj_4712), .I1(n31_adj_4710), .I2(n29_adj_4709), 
            .I3(n43631), .O(n43616));
    defparam i36491_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 rem_4_add_1988_9_lut (.I0(GND_net), .I1(n2951), .I2(VCC_net), 
            .I3(n30980), .O(n3018)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_9 (.CI(n30980), .I0(n2951), .I1(VCC_net), 
            .CO(n30981));
    SB_LUT4 div_36_unary_minus_2_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4553), .I3(n31265), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_8_lut (.I0(GND_net), .I1(n2952), .I2(VCC_net), 
            .I3(n30979), .O(n3019)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n29_adj_4965), .I3(n32306), .O(n29_adj_4380)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_2_add_3_17 (.CI(n31265), .I0(GND_net), .I1(n10_adj_4553), 
            .CO(n31266));
    SB_LUT4 div_36_unary_minus_2_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4554), .I3(n31264), .O(n11_adj_4382)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_8 (.CI(n30979), .I0(n2952), .I1(VCC_net), 
            .CO(n30980));
    SB_CARRY rem_4_unary_minus_2_add_3_6 (.CI(n32306), .I0(GND_net), .I1(n29_adj_4965), 
            .CO(n32307));
    SB_LUT4 rem_4_unary_minus_2_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n30_adj_4966), .I3(n32305), .O(n30_adj_4379)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_2_add_3_16 (.CI(n31264), .I0(GND_net), .I1(n11_adj_4554), 
            .CO(n31265));
    SB_CARRY rem_4_unary_minus_2_add_3_5 (.CI(n32305), .I0(GND_net), .I1(n30_adj_4966), 
            .CO(n32306));
    SB_LUT4 div_36_unary_minus_2_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4555), .I3(n31263), .O(n12_adj_4366)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n31_adj_4967), .I3(n32304), .O(n31_adj_4378)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_7_lut (.I0(GND_net), .I1(n2953), .I2(VCC_net), 
            .I3(n30978), .O(n3020)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_7 (.CI(n30978), .I0(n2953), .I1(VCC_net), 
            .CO(n30979));
    SB_LUT4 rem_4_add_1988_6_lut (.I0(GND_net), .I1(n2954), .I2(GND_net), 
            .I3(n30977), .O(n3021)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_2_add_3_15 (.CI(n31263), .I0(GND_net), .I1(n12_adj_4555), 
            .CO(n31264));
    SB_CARRY rem_4_add_1988_6 (.CI(n30977), .I0(n2954), .I1(GND_net), 
            .CO(n30978));
    SB_CARRY rem_4_unary_minus_2_add_3_4 (.CI(n32304), .I0(GND_net), .I1(n31_adj_4967), 
            .CO(n32305));
    SB_LUT4 rem_4_add_1988_5_lut (.I0(GND_net), .I1(n2955), .I2(GND_net), 
            .I3(n30976), .O(n3022)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_5 (.CI(n30976), .I0(n2955), .I1(GND_net), 
            .CO(n30977));
    SB_LUT4 rem_4_add_1988_4_lut (.I0(GND_net), .I1(n2956), .I2(VCC_net), 
            .I3(n30975), .O(n3023)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_4 (.CI(n30975), .I0(n2956), .I1(VCC_net), 
            .CO(n30976));
    SB_LUT4 div_36_unary_minus_2_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4556), .I3(n31262), .O(n13_adj_4375)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_3_lut (.I0(GND_net), .I1(n2957), .I2(VCC_net), 
            .I3(n30974), .O(n3024)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_3 (.CI(n30974), .I0(n2957), .I1(VCC_net), 
            .CO(n30975));
    SB_LUT4 rem_4_add_1988_2_lut (.I0(GND_net), .I1(n2958), .I2(GND_net), 
            .I3(VCC_net), .O(n3025)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_2 (.CI(VCC_net), .I0(n2958), .I1(GND_net), 
            .CO(n30974));
    SB_CARRY div_36_unary_minus_2_add_3_14 (.CI(n31262), .I0(GND_net), .I1(n13_adj_4556), 
            .CO(n31263));
    SB_LUT4 rem_4_unary_minus_2_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n32_adj_4968), .I3(n32303), .O(n32_adj_4377)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3167_25_lut (.I0(n249), .I1(n45862), .I2(n248), .I3(n30973), 
            .O(displacement_23__N_229[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3167_24_lut (.I0(n393), .I1(n45862), .I2(n392), .I3(n30972), 
            .O(displacement_23__N_229[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3167_24 (.CI(n30972), .I0(n45862), .I1(n392), .CO(n30973));
    SB_LUT4 add_3167_23_lut (.I0(n534), .I1(n45862), .I2(n533), .I3(n30971), 
            .O(displacement_23__N_229[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_36_unary_minus_2_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4557), .I3(n31261), .O(n14)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_3 (.CI(n32303), .I0(GND_net), .I1(n32_adj_4968), 
            .CO(n32304));
    SB_CARRY add_3167_23 (.CI(n30971), .I0(n45862), .I1(n533), .CO(n30972));
    SB_LUT4 add_3167_22_lut (.I0(n672), .I1(n45862), .I2(n671), .I3(n30970), 
            .O(displacement_23__N_229[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY div_36_unary_minus_2_add_3_13 (.CI(n31261), .I0(GND_net), .I1(n14_adj_4557), 
            .CO(n31262));
    SB_LUT4 div_36_LessThan_1350_i20_4_lut (.I0(n383), .I1(n99), .I2(n2083), 
            .I3(n558), .O(n20_adj_4700));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1350_i20_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_36_LessThan_1350_i28_3_lut (.I0(n26_adj_4706), .I1(n93), 
            .I2(n31_adj_4710), .I3(GND_net), .O(n28_adj_4708));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1350_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_unary_minus_2_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n33_adj_4969), .I3(VCC_net), .O(n33_adj_4376)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3167_22 (.CI(n30970), .I0(n45862), .I1(n671), .CO(n30971));
    SB_LUT4 add_3167_21_lut (.I0(n807), .I1(n45862), .I2(n806), .I3(n30969), 
            .O(displacement_23__N_229[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_unary_minus_2_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n33_adj_4969), 
            .CO(n32303));
    SB_LUT4 div_36_unary_minus_2_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4558), .I3(n31260), .O(n15_adj_4363)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3167_21 (.CI(n30969), .I0(n45862), .I1(n806), .CO(n30970));
    SB_LUT4 add_3167_20_lut (.I0(n939), .I1(n45862), .I2(n938), .I3(n30968), 
            .O(displacement_23__N_229[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY div_36_unary_minus_2_add_3_12 (.CI(n31260), .I0(GND_net), .I1(n15_adj_4558), 
            .CO(n31261));
    SB_CARRY add_3167_20 (.CI(n30968), .I0(n45862), .I1(n938), .CO(n30969));
    SB_LUT4 div_36_unary_minus_2_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4559), .I3(n31259), .O(n16_adj_4411)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_2_add_3_11 (.CI(n31259), .I0(GND_net), .I1(n16_adj_4559), 
            .CO(n31260));
    SB_LUT4 add_3167_19_lut (.I0(n1068), .I1(n45862), .I2(n1067), .I3(n30967), 
            .O(displacement_23__N_229[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3167_19 (.CI(n30967), .I0(n45862), .I1(n1067), .CO(n30968));
    SB_LUT4 div_36_unary_minus_2_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4560), .I3(n31258), .O(n17_adj_4410)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3167_18_lut (.I0(n1194), .I1(n45862), .I2(n1193), .I3(n30966), 
            .O(displacement_23__N_229[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3167_18 (.CI(n30966), .I0(n45862), .I1(n1193), .CO(n30967));
    SB_CARRY div_36_unary_minus_2_add_3_10 (.CI(n31258), .I0(GND_net), .I1(n17_adj_4560), 
            .CO(n31259));
    SB_LUT4 div_36_unary_minus_2_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4561), .I3(n31257), .O(n18_adj_4344)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3167_17_lut (.I0(n1317), .I1(n45862), .I2(n1316), .I3(n30965), 
            .O(displacement_23__N_229[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY div_36_unary_minus_2_add_3_9 (.CI(n31257), .I0(GND_net), .I1(n18_adj_4561), 
            .CO(n31258));
    SB_CARRY add_3167_17 (.CI(n30965), .I0(n45862), .I1(n1316), .CO(n30966));
    SB_LUT4 div_36_unary_minus_2_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4562), .I3(n31256), .O(n19_adj_4343)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3167_16_lut (.I0(n1437), .I1(n45862), .I2(n1436), .I3(n30964), 
            .O(displacement_23__N_229[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3167_16 (.CI(n30964), .I0(n45862), .I1(n1436), .CO(n30965));
    SB_LUT4 add_3167_15_lut (.I0(n1554), .I1(n45862), .I2(n1553), .I3(n30963), 
            .O(displacement_23__N_229[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3167_15 (.CI(n30963), .I0(n45862), .I1(n1553), .CO(n30964));
    SB_LUT4 add_3167_14_lut (.I0(n1668), .I1(n45862), .I2(n1667), .I3(n30962), 
            .O(displacement_23__N_229[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3167_14 (.CI(n30962), .I0(n45862), .I1(n1667), .CO(n30963));
    SB_LUT4 add_3167_13_lut (.I0(n1779), .I1(n45862), .I2(n1778), .I3(n30961), 
            .O(displacement_23__N_229[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY div_36_unary_minus_2_add_3_8 (.CI(n31256), .I0(GND_net), .I1(n19_adj_4562), 
            .CO(n31257));
    SB_LUT4 div_36_unary_minus_2_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4563), .I3(n31255), .O(n20_adj_4342)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_2_add_3_7 (.CI(n31255), .I0(GND_net), .I1(n20_adj_4563), 
            .CO(n31256));
    SB_CARRY add_3167_13 (.CI(n30961), .I0(n45862), .I1(n1778), .CO(n30962));
    SB_LUT4 add_3167_12_lut (.I0(n1887), .I1(n45862), .I2(n1886), .I3(n30960), 
            .O(displacement_23__N_229[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3167_12 (.CI(n30960), .I0(n45862), .I1(n1886), .CO(n30961));
    SB_LUT4 add_3167_11_lut (.I0(n1992), .I1(n45862), .I2(n1991), .I3(n30959), 
            .O(displacement_23__N_229[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3167_11 (.CI(n30959), .I0(n45862), .I1(n1991), .CO(n30960));
    SB_LUT4 add_3167_10_lut (.I0(n2094), .I1(n45862), .I2(n2093), .I3(n30958), 
            .O(displacement_23__N_229[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3167_10 (.CI(n30958), .I0(n45862), .I1(n2093), .CO(n30959));
    SB_LUT4 add_3167_9_lut (.I0(n2193), .I1(n45862), .I2(n2192), .I3(n30957), 
            .O(displacement_23__N_229[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3167_9 (.CI(n30957), .I0(n45862), .I1(n2192), .CO(n30958));
    SB_LUT4 add_3167_8_lut (.I0(n2289), .I1(n45862), .I2(n2288), .I3(n30956), 
            .O(displacement_23__N_229[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3167_8 (.CI(n30956), .I0(n45862), .I1(n2288), .CO(n30957));
    SB_LUT4 add_3167_7_lut (.I0(n2382), .I1(n45862), .I2(n2381), .I3(n30955), 
            .O(displacement_23__N_229[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3167_7 (.CI(n30955), .I0(n45862), .I1(n2381), .CO(n30956));
    SB_LUT4 add_3167_6_lut (.I0(n2472), .I1(n45862), .I2(n2471), .I3(n30954), 
            .O(displacement_23__N_229[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3167_6 (.CI(n30954), .I0(n45862), .I1(n2471), .CO(n30955));
    SB_LUT4 div_36_unary_minus_2_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4564), .I3(n31254), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_2_add_3_6 (.CI(n31254), .I0(GND_net), .I1(n21_adj_4564), 
            .CO(n31255));
    SB_LUT4 div_36_unary_minus_2_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4565), .I3(n31253), .O(n22)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_2_add_3_5 (.CI(n31253), .I0(GND_net), .I1(n22_adj_4565), 
            .CO(n31254));
    SB_LUT4 div_36_unary_minus_2_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4566), .I3(n31252), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_2_add_3_4 (.CI(n31252), .I0(GND_net), .I1(n23_adj_4566), 
            .CO(n31253));
    SB_LUT4 div_36_unary_minus_2_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4567), .I3(n31251), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_2_add_3_3 (.CI(n31251), .I0(GND_net), .I1(n24_adj_4567), 
            .CO(n31252));
    SB_LUT4 div_36_LessThan_1350_i32_3_lut (.I0(n24_adj_4704), .I1(n91), 
            .I2(n35_adj_4713), .I3(GND_net), .O(n32_adj_4711));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1350_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37845_4_lut (.I0(n32_adj_4711), .I1(n22_adj_4702), .I2(n35_adj_4713), 
            .I3(n43613), .O(n44970));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37845_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i37846_3_lut (.I0(n44970), .I1(n90), .I2(n37_adj_4714), .I3(GND_net), 
            .O(n44971));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37846_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3167_5_lut (.I0(n2559), .I1(n45862), .I2(n2558), .I3(n30953), 
            .O(displacement_23__N_229[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_5_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_36_unary_minus_2_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4568), .I3(VCC_net), .O(n25_adj_4364)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37718_3_lut (.I0(n44971), .I1(n89), .I2(n39_adj_4715), .I3(GND_net), 
            .O(n44843));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37718_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3167_5 (.CI(n30953), .I0(n45862), .I1(n2558), .CO(n30954));
    SB_CARRY div_36_unary_minus_2_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4568), 
            .CO(n31251));
    SB_LUT4 div_36_unary_minus_4_add_3_25_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(n2_adj_4521), .I3(n31250), .O(n77)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_553_24_lut (.I0(duty[22]), .I1(n45865), .I2(n3_adj_4327), 
            .I3(n30454), .O(pwm_setpoint_22__N_57[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_36_unary_minus_4_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4522), .I3(n31249), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37639_4_lut (.I0(n39_adj_4715), .I1(n37_adj_4714), .I2(n35_adj_4713), 
            .I3(n43616), .O(n44764));
    defparam i37639_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i37847_4_lut (.I0(n28_adj_4708), .I1(n20_adj_4700), .I2(n31_adj_4710), 
            .I3(n43625), .O(n44972));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37847_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36823_3_lut (.I0(n44843), .I1(n88), .I2(n41_adj_4716), .I3(GND_net), 
            .O(n43948));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36823_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37928_4_lut (.I0(n43948), .I1(n44972), .I2(n41_adj_4716), 
            .I3(n44764), .O(n45053));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37928_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i37929_3_lut (.I0(n45053), .I1(n87), .I2(n2071), .I3(GND_net), 
            .O(n45054));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37929_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i37872_3_lut (.I0(n45054), .I1(n86), .I2(n2070), .I3(GND_net), 
            .O(n44997));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37872_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1701 (.I0(n44997), .I1(n17305), .I2(n85), .I3(n2069), 
            .O(n2093));
    defparam i1_4_lut_adj_1701.LUT_INIT = 16'hceef;
    SB_LUT4 div_36_LessThan_1281_i43_2_lut (.I0(n1969), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4698));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1281_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1281_i41_2_lut (.I0(n1970), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4697));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1281_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1281_i39_2_lut (.I0(n1971), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4696));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1281_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1281_i37_2_lut (.I0(n1972), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4695));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1281_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_mux_3_i10_3_lut (.I0(encoder0_position[9]), .I1(n16_adj_4411), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n382));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1281_i31_2_lut (.I0(n1975), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4691));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1281_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1281_i33_2_lut (.I0(n1974), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4692));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1281_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1281_i35_2_lut (.I0(n1973), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4694));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1281_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1281_i25_2_lut (.I0(n1978), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4685));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1281_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1281_i27_2_lut (.I0(n1977), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4687));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1281_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1281_i29_2_lut (.I0(n1976), .I1(n95_adj_4360), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4689));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1281_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_i1283_1_lut (.I0(n1991), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1992));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1283_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_1281_i23_2_lut (.I0(n1979), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4683));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1281_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i36559_4_lut (.I0(n29_adj_4689), .I1(n27_adj_4687), .I2(n25_adj_4685), 
            .I3(n23_adj_4683), .O(n43684));
    defparam i36559_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36553_4_lut (.I0(n35_adj_4694), .I1(n33_adj_4692), .I2(n31_adj_4691), 
            .I3(n43684), .O(n43678));
    defparam i36553_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_36_LessThan_1281_i22_4_lut (.I0(n382), .I1(n99), .I2(n1980), 
            .I3(n558), .O(n22_adj_4682));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1281_i22_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_36_LessThan_1281_i30_3_lut (.I0(n28_adj_4688), .I1(n93), 
            .I2(n33_adj_4692), .I3(GND_net), .O(n30_adj_4690));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1281_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_36_LessThan_1281_i34_3_lut (.I0(n26_adj_4686), .I1(n91), 
            .I2(n37_adj_4695), .I3(GND_net), .O(n34_adj_4693));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1281_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37843_4_lut (.I0(n34_adj_4693), .I1(n24_adj_4684), .I2(n37_adj_4695), 
            .I3(n43676), .O(n44968));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37843_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i37844_3_lut (.I0(n44968), .I1(n90), .I2(n39_adj_4696), .I3(GND_net), 
            .O(n44969));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37844_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37724_3_lut (.I0(n44969), .I1(n89), .I2(n41_adj_4697), .I3(GND_net), 
            .O(n44849));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37724_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37645_4_lut (.I0(n41_adj_4697), .I1(n39_adj_4696), .I2(n37_adj_4695), 
            .I3(n43678), .O(n44770));
    defparam i37645_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i37831_4_lut (.I0(n30_adj_4690), .I1(n22_adj_4682), .I2(n33_adj_4692), 
            .I3(n43680), .O(n44956));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37831_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY div_36_unary_minus_4_add_3_24 (.CI(n31249), .I0(GND_net), .I1(n3_adj_4522), 
            .CO(n31250));
    SB_LUT4 add_553_23_lut (.I0(duty[21]), .I1(n45865), .I2(n4_adj_4328), 
            .I3(n30453), .O(pwm_setpoint_22__N_57[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3167_4_lut (.I0(n2643), .I1(n45862), .I2(n2642), .I3(n30952), 
            .O(displacement_23__N_229[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i36819_3_lut (.I0(n44849), .I1(n88), .I2(n43_adj_4698), .I3(GND_net), 
            .O(n43944));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36819_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_36_unary_minus_4_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4523), .I3(n31248), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37920_4_lut (.I0(n43944), .I1(n44956), .I2(n43_adj_4698), 
            .I3(n44770), .O(n45045));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37920_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i37921_3_lut (.I0(n45045), .I1(n87), .I2(n1968), .I3(GND_net), 
            .O(n45046));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37921_3_lut.LUT_INIT = 16'h2b2b;
    SB_CARRY div_36_unary_minus_4_add_3_23 (.CI(n31248), .I0(GND_net), .I1(n4_adj_4523), 
            .CO(n31249));
    SB_LUT4 div_36_unary_minus_4_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4524), .I3(n31247), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3167_4 (.CI(n30952), .I0(n45862), .I1(n2642), .CO(n30953));
    SB_LUT4 add_3167_3_lut (.I0(n2724), .I1(n45862), .I2(n2723), .I3(n30951), 
            .O(displacement_23__N_229[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_3_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_4_lut_adj_1702 (.I0(n45046), .I1(n17302), .I2(n86), .I3(n1967), 
            .O(n1991));
    defparam i1_4_lut_adj_1702.LUT_INIT = 16'hceef;
    SB_CARRY add_553_23 (.CI(n30453), .I0(n45865), .I1(n4_adj_4328), .CO(n30454));
    SB_CARRY div_36_unary_minus_4_add_3_22 (.CI(n31247), .I0(GND_net), .I1(n5_adj_4524), 
            .CO(n31248));
    SB_LUT4 rem_4_i1732_3_lut (.I0(n2547_adj_4515), .I1(n2614), .I2(n2570), 
            .I3(GND_net), .O(n2646));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1210_i45_2_lut (.I0(n1863), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4680));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1210_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1210_i43_2_lut (.I0(n1864), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4679));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1210_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i1735_3_lut (.I0(n2550_adj_4512), .I1(n2617), .I2(n2570), 
            .I3(GND_net), .O(n2649));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1210_i41_2_lut (.I0(n1865), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4678));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1210_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i1737_3_lut (.I0(n2552_adj_4510), .I1(n2619_adj_4506), 
            .I2(n2570), .I3(GND_net), .O(n2651));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1210_i39_2_lut (.I0(n1866), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4677));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1210_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_mux_3_i11_3_lut (.I0(encoder0_position[10]), .I1(n15_adj_4363), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n381));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1210_i33_2_lut (.I0(n1869), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4673));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1210_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1210_i35_2_lut (.I0(n1868), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4674));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1210_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1210_i37_2_lut (.I0(n1867), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4676));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1210_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1210_i27_2_lut (.I0(n1872), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4667));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1210_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1210_i29_2_lut (.I0(n1871), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4669));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1210_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1210_i31_2_lut (.I0(n1870), .I1(n95_adj_4360), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4671));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1210_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_i1212_1_lut (.I0(n1886), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1887));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1212_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_1210_i25_2_lut (.I0(n1873), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4665));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1210_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i35880_4_lut (.I0(n31_adj_4671), .I1(n29_adj_4669), .I2(n27_adj_4667), 
            .I3(n25_adj_4665), .O(n43004));
    defparam i35880_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35869_4_lut (.I0(n37_adj_4676), .I1(n35_adj_4674), .I2(n33_adj_4673), 
            .I3(n43004), .O(n42993));
    defparam i35869_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_36_LessThan_1210_i24_4_lut (.I0(n381), .I1(n99), .I2(n1874), 
            .I3(n558), .O(n24_adj_4664));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1210_i24_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_36_LessThan_1210_i32_3_lut (.I0(n30_adj_4670), .I1(n93), 
            .I2(n35_adj_4674), .I3(GND_net), .O(n32_adj_4672));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1210_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_36_LessThan_1210_i36_3_lut (.I0(n28_adj_4668), .I1(n91), 
            .I2(n39_adj_4677), .I3(GND_net), .O(n36_adj_4675));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1210_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37841_4_lut (.I0(n36_adj_4675), .I1(n26_adj_4666), .I2(n39_adj_4677), 
            .I3(n43727), .O(n44966));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37841_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i37842_3_lut (.I0(n44966), .I1(n90), .I2(n41_adj_4678), .I3(GND_net), 
            .O(n44967));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37842_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37728_3_lut (.I0(n44967), .I1(n89), .I2(n43_adj_4679), .I3(GND_net), 
            .O(n44853));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37728_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37428_4_lut (.I0(n43_adj_4679), .I1(n41_adj_4678), .I2(n39_adj_4677), 
            .I3(n42993), .O(n44553));
    defparam i37428_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i37536_4_lut (.I0(n32_adj_4672), .I1(n24_adj_4664), .I2(n35_adj_4674), 
            .I3(n43002), .O(n44661));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37536_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36815_3_lut (.I0(n44853), .I1(n88), .I2(n45_adj_4680), .I3(GND_net), 
            .O(n43940));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36815_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37538_4_lut (.I0(n43940), .I1(n44661), .I2(n45_adj_4680), 
            .I3(n44553), .O(n44663));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37538_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1703 (.I0(n44663), .I1(n17225), .I2(n87), .I3(n1862), 
            .O(n1886));
    defparam i1_4_lut_adj_1703.LUT_INIT = 16'hceef;
    SB_CARRY add_3167_3 (.CI(n30951), .I0(n45862), .I1(n2723), .CO(n30952));
    SB_LUT4 add_3167_2_lut (.I0(n2802), .I1(n45862), .I2(n2801), .I3(VCC_net), 
            .O(displacement_23__N_229[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3167_2_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_36_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4563));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3167_2 (.CI(VCC_net), .I0(n45862), .I1(n2801), .CO(n30951));
    SB_LUT4 div_36_unary_minus_4_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4525), .I3(n31246), .O(n56)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3166_25_lut (.I0(GND_net), .I1(n2699), .I2(n78), .I3(n30950), 
            .O(n7160)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3166_24_lut (.I0(GND_net), .I1(n2700), .I2(n79), .I3(n30949), 
            .O(n7161)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13726_2_lut (.I0(n18897), .I1(n18756), .I2(GND_net), .I3(GND_net), 
            .O(n18758));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13726_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3166_24 (.CI(n30949), .I0(n2700), .I1(n79), .CO(n30950));
    SB_CARRY div_36_unary_minus_4_add_3_21 (.CI(n31246), .I0(GND_net), .I1(n6_adj_4525), 
            .CO(n31247));
    SB_LUT4 div_36_unary_minus_4_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4526), .I3(n31245), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_4_add_3_20 (.CI(n31245), .I0(GND_net), .I1(n7_adj_4526), 
            .CO(n31246));
    SB_LUT4 add_3166_23_lut (.I0(GND_net), .I1(n2701), .I2(n80), .I3(n30948), 
            .O(n7162)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_23 (.CI(n30948), .I0(n2701), .I1(n80), .CO(n30949));
    SB_LUT4 add_3166_22_lut (.I0(GND_net), .I1(n2702), .I2(n81), .I3(n30947), 
            .O(n7163)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_1137_i37_2_lut (.I0(n1759), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4660));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1137_i37_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3166_22 (.CI(n30947), .I0(n2702), .I1(n81), .CO(n30948));
    SB_LUT4 add_3166_21_lut (.I0(GND_net), .I1(n2703), .I2(n82), .I3(n30946), 
            .O(n7164)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_21 (.CI(n30946), .I0(n2703), .I1(n82), .CO(n30947));
    SB_LUT4 add_3166_20_lut (.I0(GND_net), .I1(n2704), .I2(n83), .I3(n30945), 
            .O(n7165)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_20 (.CI(n30945), .I0(n2704), .I1(n83), .CO(n30946));
    SB_LUT4 add_3166_19_lut (.I0(GND_net), .I1(n2705), .I2(n84), .I3(n30944), 
            .O(n7166)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_19 (.CI(n30944), .I0(n2705), .I1(n84), .CO(n30945));
    SB_LUT4 add_553_22_lut (.I0(duty[20]), .I1(n45865), .I2(n5), .I3(n30452), 
            .O(pwm_setpoint_22__N_57[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_36_unary_minus_4_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4527), .I3(n31244), .O(n58)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_553_22 (.CI(n30452), .I0(n45865), .I1(n5), .CO(n30453));
    SB_LUT4 add_3166_18_lut (.I0(GND_net), .I1(n2706), .I2(n85), .I3(n30943), 
            .O(n7167)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_18 (.CI(n30943), .I0(n2706), .I1(n85), .CO(n30944));
    SB_LUT4 add_3166_17_lut (.I0(GND_net), .I1(n2707), .I2(n86), .I3(n30942), 
            .O(n7168)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_17 (.CI(n30942), .I0(n2707), .I1(n86), .CO(n30943));
    SB_LUT4 add_3166_16_lut (.I0(GND_net), .I1(n2708), .I2(n87), .I3(n30941), 
            .O(n7169)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_16 (.CI(n30941), .I0(n2708), .I1(n87), .CO(n30942));
    SB_LUT4 add_3166_15_lut (.I0(GND_net), .I1(n2709), .I2(n88), .I3(n30940), 
            .O(n7170)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_15 (.CI(n30940), .I0(n2709), .I1(n88), .CO(n30941));
    SB_LUT4 div_36_LessThan_1137_i35_2_lut (.I0(n1760), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4659));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1137_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_553_21_lut (.I0(duty[19]), .I1(n45865), .I2(n6), .I3(n30451), 
            .O(pwm_setpoint_22__N_57[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_553_21 (.CI(n30451), .I0(n45865), .I1(n6), .CO(n30452));
    SB_CARRY div_36_unary_minus_4_add_3_19 (.CI(n31244), .I0(GND_net), .I1(n8_adj_4527), 
            .CO(n31245));
    SB_LUT4 div_36_unary_minus_4_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4528), .I3(n31243), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_4_add_3_18 (.CI(n31243), .I0(GND_net), .I1(n9_adj_4528), 
            .CO(n31244));
    SB_LUT4 add_553_20_lut (.I0(duty[18]), .I1(n45865), .I2(n7_adj_4329), 
            .I3(n30450), .O(pwm_setpoint_22__N_57[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3166_14_lut (.I0(GND_net), .I1(n2710), .I2(n89), .I3(n30939), 
            .O(n7171)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_unary_minus_4_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4529), .I3(n31242), .O(n60)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_14 (.CI(n30939), .I0(n2710), .I1(n89), .CO(n30940));
    SB_CARRY div_36_unary_minus_4_add_3_17 (.CI(n31242), .I0(GND_net), .I1(n10_adj_4529), 
            .CO(n31243));
    SB_LUT4 add_3166_13_lut (.I0(GND_net), .I1(n2711), .I2(n90), .I3(n30938), 
            .O(n7172)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_13 (.CI(n30938), .I0(n2711), .I1(n90), .CO(n30939));
    SB_LUT4 add_3166_12_lut (.I0(GND_net), .I1(n2712), .I2(n91), .I3(n30937), 
            .O(n7173)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_12 (.CI(n30937), .I0(n2712), .I1(n91), .CO(n30938));
    SB_LUT4 add_3166_11_lut (.I0(GND_net), .I1(n2713), .I2(n92), .I3(n30936), 
            .O(n7174)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_11 (.CI(n30936), .I0(n2713), .I1(n92), .CO(n30937));
    SB_LUT4 add_3166_10_lut (.I0(GND_net), .I1(n2714), .I2(n93), .I3(n30935), 
            .O(n7175)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_10 (.CI(n30935), .I0(n2714), .I1(n93), .CO(n30936));
    SB_LUT4 add_3166_9_lut (.I0(GND_net), .I1(n2715), .I2(n94), .I3(n30934), 
            .O(n7176)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_9 (.CI(n30934), .I0(n2715), .I1(n94), .CO(n30935));
    SB_LUT4 add_3166_8_lut (.I0(GND_net), .I1(n2716), .I2(n95_adj_4360), 
            .I3(n30933), .O(n7177)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_8 (.CI(n30933), .I0(n2716), .I1(n95_adj_4360), .CO(n30934));
    SB_LUT4 add_3166_7_lut (.I0(GND_net), .I1(n2717), .I2(n96), .I3(n30932), 
            .O(n7178)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_7 (.CI(n30932), .I0(n2717), .I1(n96), .CO(n30933));
    SB_LUT4 add_3166_6_lut (.I0(GND_net), .I1(n2718), .I2(n97), .I3(n30931), 
            .O(n7179)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_6 (.CI(n30931), .I0(n2718), .I1(n97), .CO(n30932));
    SB_LUT4 add_3166_5_lut (.I0(GND_net), .I1(n2719), .I2(n98), .I3(n30930), 
            .O(n7180)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_5 (.CI(n30930), .I0(n2719), .I1(n98), .CO(n30931));
    SB_LUT4 add_3166_4_lut (.I0(GND_net), .I1(n2720), .I2(n99), .I3(n30929), 
            .O(n7181)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_4 (.CI(n30929), .I0(n2720), .I1(n99), .CO(n30930));
    SB_LUT4 add_3166_3_lut (.I0(GND_net), .I1(n390), .I2(n558), .I3(n30928), 
            .O(n7182)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3166_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3166_3 (.CI(n30928), .I0(n390), .I1(n558), .CO(n30929));
    SB_CARRY add_3166_2 (.CI(VCC_net), .I0(n391), .I1(VCC_net), .CO(n30928));
    SB_LUT4 add_3165_23_lut (.I0(GND_net), .I1(n2618), .I2(n79), .I3(n30927), 
            .O(n7136)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3165_22_lut (.I0(GND_net), .I1(n2619), .I2(n80), .I3(n30926), 
            .O(n7137)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_22 (.CI(n30926), .I0(n2619), .I1(n80), .CO(n30927));
    SB_LUT4 add_3165_21_lut (.I0(GND_net), .I1(n2620), .I2(n81), .I3(n30925), 
            .O(n7138)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_21 (.CI(n30925), .I0(n2620), .I1(n81), .CO(n30926));
    SB_LUT4 add_3165_20_lut (.I0(GND_net), .I1(n2621), .I2(n82), .I3(n30924), 
            .O(n7139)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_20 (.CI(n30924), .I0(n2621), .I1(n82), .CO(n30925));
    SB_LUT4 add_3165_19_lut (.I0(GND_net), .I1(n2622), .I2(n83), .I3(n30923), 
            .O(n7140)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_unary_minus_4_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4530), .I3(n31241), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_4_add_3_16 (.CI(n31241), .I0(GND_net), .I1(n11_adj_4530), 
            .CO(n31242));
    SB_LUT4 div_36_unary_minus_4_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4531), .I3(n31240), .O(n62)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_4_add_3_15 (.CI(n31240), .I0(GND_net), .I1(n12_adj_4531), 
            .CO(n31241));
    SB_LUT4 div_36_unary_minus_4_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4532), .I3(n31239), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_mux_3_i12_3_lut (.I0(encoder0_position[11]), .I1(n14), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n380));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_36_unary_minus_4_add_3_14 (.CI(n31239), .I0(GND_net), .I1(n13_adj_4532), 
            .CO(n31240));
    SB_LUT4 div_36_LessThan_1137_i41_2_lut (.I0(n1757), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4663));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1137_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1137_i39_2_lut (.I0(n1758), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4662));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1137_i39_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3165_19 (.CI(n30923), .I0(n2622), .I1(n83), .CO(n30924));
    SB_LUT4 add_3165_18_lut (.I0(GND_net), .I1(n2623), .I2(n84), .I3(n30922), 
            .O(n7141)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_18 (.CI(n30922), .I0(n2623), .I1(n84), .CO(n30923));
    SB_LUT4 add_3165_17_lut (.I0(GND_net), .I1(n2624), .I2(n85), .I3(n30921), 
            .O(n7142)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_17 (.CI(n30921), .I0(n2624), .I1(n85), .CO(n30922));
    SB_LUT4 add_3165_16_lut (.I0(GND_net), .I1(n2625), .I2(n86), .I3(n30920), 
            .O(n7143)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_16 (.CI(n30920), .I0(n2625), .I1(n86), .CO(n30921));
    SB_LUT4 add_3165_15_lut (.I0(GND_net), .I1(n2626), .I2(n87), .I3(n30919), 
            .O(n7144)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_15 (.CI(n30919), .I0(n2626), .I1(n87), .CO(n30920));
    SB_LUT4 add_3165_14_lut (.I0(GND_net), .I1(n2627), .I2(n88), .I3(n30918), 
            .O(n7145)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_14 (.CI(n30918), .I0(n2627), .I1(n88), .CO(n30919));
    SB_LUT4 add_3165_13_lut (.I0(GND_net), .I1(n2628), .I2(n89), .I3(n30917), 
            .O(n7146)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_13 (.CI(n30917), .I0(n2628), .I1(n89), .CO(n30918));
    SB_LUT4 add_3165_12_lut (.I0(GND_net), .I1(n2629), .I2(n90), .I3(n30916), 
            .O(n7147)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_12 (.CI(n30916), .I0(n2629), .I1(n90), .CO(n30917));
    SB_LUT4 add_3165_11_lut (.I0(GND_net), .I1(n2630), .I2(n91), .I3(n30915), 
            .O(n7148)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_11 (.CI(n30915), .I0(n2630), .I1(n91), .CO(n30916));
    SB_LUT4 add_3165_10_lut (.I0(GND_net), .I1(n2631), .I2(n92), .I3(n30914), 
            .O(n7149)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_10 (.CI(n30914), .I0(n2631), .I1(n92), .CO(n30915));
    SB_LUT4 add_3165_9_lut (.I0(GND_net), .I1(n2632), .I2(n93), .I3(n30913), 
            .O(n7150)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_9 (.CI(n30913), .I0(n2632), .I1(n93), .CO(n30914));
    SB_LUT4 add_3165_8_lut (.I0(GND_net), .I1(n2633), .I2(n94), .I3(n30912), 
            .O(n7151)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_8 (.CI(n30912), .I0(n2633), .I1(n94), .CO(n30913));
    SB_LUT4 add_3165_7_lut (.I0(GND_net), .I1(n2634), .I2(n95_adj_4360), 
            .I3(n30911), .O(n7152)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_7 (.CI(n30911), .I0(n2634), .I1(n95_adj_4360), .CO(n30912));
    SB_LUT4 add_3165_6_lut (.I0(GND_net), .I1(n2635), .I2(n96), .I3(n30910), 
            .O(n7153)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_1137_i29_2_lut (.I0(n1763), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4655));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1137_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1137_i31_2_lut (.I0(n1762), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4657));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1137_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1137_i33_2_lut (.I0(n1761), .I1(n95_adj_4360), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4658));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1137_i33_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3165_6 (.CI(n30910), .I0(n2635), .I1(n96), .CO(n30911));
    SB_LUT4 add_3165_5_lut (.I0(GND_net), .I1(n2636), .I2(n97), .I3(n30909), 
            .O(n7154)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i1139_1_lut (.I0(n1778), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1779));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1139_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_4_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4533), .I3(n31238), .O(n64)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_553_20 (.CI(n30450), .I0(n45865), .I1(n7_adj_4329), .CO(n30451));
    SB_CARRY div_36_unary_minus_4_add_3_13 (.CI(n31238), .I0(GND_net), .I1(n14_adj_4533), 
            .CO(n31239));
    SB_CARRY add_3165_5 (.CI(n30909), .I0(n2636), .I1(n97), .CO(n30910));
    SB_LUT4 add_3165_4_lut (.I0(GND_net), .I1(n2637), .I2(n98), .I3(n30908), 
            .O(n7155)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_4 (.CI(n30908), .I0(n2637), .I1(n98), .CO(n30909));
    SB_LUT4 add_3165_3_lut (.I0(GND_net), .I1(n2638), .I2(n99), .I3(n30907), 
            .O(n7156)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_3 (.CI(n30907), .I0(n2638), .I1(n99), .CO(n30908));
    SB_LUT4 add_3165_2_lut (.I0(GND_net), .I1(n389), .I2(n558), .I3(VCC_net), 
            .O(n7157)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3165_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3165_2 (.CI(VCC_net), .I0(n389), .I1(n558), .CO(n30907));
    SB_LUT4 add_3164_22_lut (.I0(GND_net), .I1(n2534), .I2(n80), .I3(n30906), 
            .O(n7113)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3164_21_lut (.I0(GND_net), .I1(n2535), .I2(n81), .I3(n30905), 
            .O(n7114)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_21 (.CI(n30905), .I0(n2535), .I1(n81), .CO(n30906));
    SB_LUT4 add_3164_20_lut (.I0(GND_net), .I1(n2536), .I2(n82), .I3(n30904), 
            .O(n7115)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_20 (.CI(n30904), .I0(n2536), .I1(n82), .CO(n30905));
    SB_LUT4 add_3164_19_lut (.I0(GND_net), .I1(n2537), .I2(n83), .I3(n30903), 
            .O(n7116)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_19 (.CI(n30903), .I0(n2537), .I1(n83), .CO(n30904));
    SB_LUT4 add_3164_18_lut (.I0(GND_net), .I1(n2538), .I2(n84), .I3(n30902), 
            .O(n7117)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_18 (.CI(n30902), .I0(n2538), .I1(n84), .CO(n30903));
    SB_LUT4 div_36_LessThan_1137_i27_2_lut (.I0(n1764), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4653));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1137_i27_2_lut.LUT_INIT = 16'h9999;
    SB_DFF communication_counter_1146__i1 (.Q(communication_counter[1]), .C(LED_c), 
           .D(n164));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_LUT4 i35910_4_lut (.I0(n33_adj_4658), .I1(n31_adj_4657), .I2(n29_adj_4655), 
            .I3(n27_adj_4653), .O(n43034));
    defparam i35910_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_36_LessThan_1137_i38_3_lut (.I0(n30_adj_4656), .I1(n91), 
            .I2(n41_adj_4663), .I3(GND_net), .O(n38_adj_4661));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1137_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_36_LessThan_1137_i26_4_lut (.I0(n380), .I1(n99), .I2(n1765), 
            .I3(n558), .O(n26_adj_4652));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1137_i26_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 add_3164_17_lut (.I0(GND_net), .I1(n2539), .I2(n85), .I3(n30901), 
            .O(n7118)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_17 (.CI(n30901), .I0(n2539), .I1(n85), .CO(n30902));
    SB_LUT4 add_3164_16_lut (.I0(GND_net), .I1(n2540), .I2(n86), .I3(n30900), 
            .O(n7119)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_16 (.CI(n30900), .I0(n2540), .I1(n86), .CO(n30901));
    SB_LUT4 add_3164_15_lut (.I0(GND_net), .I1(n2541), .I2(n87), .I3(n30899), 
            .O(n7120)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_15 (.CI(n30899), .I0(n2541), .I1(n87), .CO(n30900));
    SB_LUT4 add_3164_14_lut (.I0(GND_net), .I1(n2542), .I2(n88), .I3(n30898), 
            .O(n7121)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_14 (.CI(n30898), .I0(n2542), .I1(n88), .CO(n30899));
    SB_LUT4 add_3164_13_lut (.I0(GND_net), .I1(n2543), .I2(n89), .I3(n30897), 
            .O(n7122)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_13 (.CI(n30897), .I0(n2543), .I1(n89), .CO(n30898));
    SB_LUT4 add_3164_12_lut (.I0(GND_net), .I1(n2544), .I2(n90), .I3(n30896), 
            .O(n7123)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_12 (.CI(n30896), .I0(n2544), .I1(n90), .CO(n30897));
    SB_LUT4 add_3164_11_lut (.I0(GND_net), .I1(n2545), .I2(n91), .I3(n30895), 
            .O(n7124)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_11 (.CI(n30895), .I0(n2545), .I1(n91), .CO(n30896));
    SB_LUT4 add_3164_10_lut (.I0(GND_net), .I1(n2546), .I2(n92), .I3(n30894), 
            .O(n7125)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_10 (.CI(n30894), .I0(n2546), .I1(n92), .CO(n30895));
    SB_LUT4 add_3164_9_lut (.I0(GND_net), .I1(n2547), .I2(n93), .I3(n30893), 
            .O(n7126)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_9 (.CI(n30893), .I0(n2547), .I1(n93), .CO(n30894));
    SB_LUT4 add_3164_8_lut (.I0(GND_net), .I1(n2548), .I2(n94), .I3(n30892), 
            .O(n7127)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_8 (.CI(n30892), .I0(n2548), .I1(n94), .CO(n30893));
    SB_LUT4 add_3164_7_lut (.I0(GND_net), .I1(n2549), .I2(n95_adj_4360), 
            .I3(n30891), .O(n7128)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_7 (.CI(n30891), .I0(n2549), .I1(n95_adj_4360), .CO(n30892));
    SB_LUT4 add_3164_6_lut (.I0(GND_net), .I1(n2550), .I2(n96), .I3(n30890), 
            .O(n7129)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_6 (.CI(n30890), .I0(n2550), .I1(n96), .CO(n30891));
    SB_LUT4 add_3164_5_lut (.I0(GND_net), .I1(n2551), .I2(n97), .I3(n30889), 
            .O(n7130)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_5 (.CI(n30889), .I0(n2551), .I1(n97), .CO(n30890));
    SB_LUT4 add_3164_4_lut (.I0(GND_net), .I1(n2552), .I2(n98), .I3(n30888), 
            .O(n7131)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_4 (.CI(n30888), .I0(n2552), .I1(n98), .CO(n30889));
    SB_LUT4 add_3164_3_lut (.I0(GND_net), .I1(n2553), .I2(n99), .I3(n30887), 
            .O(n7132)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_3 (.CI(n30887), .I0(n2553), .I1(n99), .CO(n30888));
    SB_LUT4 add_3164_2_lut (.I0(GND_net), .I1(n388), .I2(n558), .I3(VCC_net), 
            .O(n7133)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3164_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3164_2 (.CI(VCC_net), .I0(n388), .I1(n558), .CO(n30887));
    SB_LUT4 add_3163_21_lut (.I0(GND_net), .I1(n2447), .I2(n81), .I3(n30886), 
            .O(n7091)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3163_20_lut (.I0(GND_net), .I1(n2448), .I2(n82), .I3(n30885), 
            .O(n7092)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_20 (.CI(n30885), .I0(n2448), .I1(n82), .CO(n30886));
    SB_LUT4 add_3163_19_lut (.I0(GND_net), .I1(n2449), .I2(n83), .I3(n30884), 
            .O(n7093)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_19 (.CI(n30884), .I0(n2449), .I1(n83), .CO(n30885));
    SB_LUT4 add_3163_18_lut (.I0(GND_net), .I1(n2450), .I2(n84), .I3(n30883), 
            .O(n7094)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_18 (.CI(n30883), .I0(n2450), .I1(n84), .CO(n30884));
    SB_LUT4 add_3163_17_lut (.I0(GND_net), .I1(n2451), .I2(n85), .I3(n30882), 
            .O(n7095)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_17 (.CI(n30882), .I0(n2451), .I1(n85), .CO(n30883));
    SB_LUT4 add_3163_16_lut (.I0(GND_net), .I1(n2452), .I2(n86), .I3(n30881), 
            .O(n7096)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_16 (.CI(n30881), .I0(n2452), .I1(n86), .CO(n30882));
    SB_LUT4 add_3163_15_lut (.I0(GND_net), .I1(n2453), .I2(n87), .I3(n30880), 
            .O(n7097)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_15 (.CI(n30880), .I0(n2453), .I1(n87), .CO(n30881));
    SB_LUT4 add_3163_14_lut (.I0(GND_net), .I1(n2454), .I2(n88), .I3(n30879), 
            .O(n7098)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_14 (.CI(n30879), .I0(n2454), .I1(n88), .CO(n30880));
    SB_LUT4 add_3163_13_lut (.I0(GND_net), .I1(n2455), .I2(n89), .I3(n30878), 
            .O(n7099)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_13 (.CI(n30878), .I0(n2455), .I1(n89), .CO(n30879));
    SB_LUT4 add_3163_12_lut (.I0(GND_net), .I1(n2456), .I2(n90), .I3(n30877), 
            .O(n7100)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_12 (.CI(n30877), .I0(n2456), .I1(n90), .CO(n30878));
    SB_LUT4 add_3163_11_lut (.I0(GND_net), .I1(n2457), .I2(n91), .I3(n30876), 
            .O(n7101)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_11 (.CI(n30876), .I0(n2457), .I1(n91), .CO(n30877));
    SB_LUT4 add_3163_10_lut (.I0(GND_net), .I1(n2458), .I2(n92), .I3(n30875), 
            .O(n7102)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_10 (.CI(n30875), .I0(n2458), .I1(n92), .CO(n30876));
    SB_LUT4 add_3163_9_lut (.I0(GND_net), .I1(n2459), .I2(n93), .I3(n30874), 
            .O(n7103)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_9 (.CI(n30874), .I0(n2459), .I1(n93), .CO(n30875));
    SB_LUT4 add_3163_8_lut (.I0(GND_net), .I1(n2460), .I2(n94), .I3(n30873), 
            .O(n7104)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_8 (.CI(n30873), .I0(n2460), .I1(n94), .CO(n30874));
    SB_LUT4 add_3163_7_lut (.I0(GND_net), .I1(n2461), .I2(n95_adj_4360), 
            .I3(n30872), .O(n7105)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_7 (.CI(n30872), .I0(n2461), .I1(n95_adj_4360), .CO(n30873));
    SB_LUT4 add_3163_6_lut (.I0(GND_net), .I1(n2462), .I2(n96), .I3(n30871), 
            .O(n7106)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_6 (.CI(n30871), .I0(n2462), .I1(n96), .CO(n30872));
    SB_LUT4 add_3163_5_lut (.I0(GND_net), .I1(n2463), .I2(n97), .I3(n30870), 
            .O(n7107)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_5 (.CI(n30870), .I0(n2463), .I1(n97), .CO(n30871));
    SB_LUT4 add_3163_4_lut (.I0(GND_net), .I1(n2464), .I2(n98), .I3(n30869), 
            .O(n7108)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_4 (.CI(n30869), .I0(n2464), .I1(n98), .CO(n30870));
    SB_LUT4 add_3163_3_lut (.I0(GND_net), .I1(n2465), .I2(n99), .I3(n30868), 
            .O(n7109)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_3 (.CI(n30868), .I0(n2465), .I1(n99), .CO(n30869));
    SB_LUT4 add_3163_2_lut (.I0(GND_net), .I1(n387), .I2(n558), .I3(VCC_net), 
            .O(n7110)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3163_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3163_2 (.CI(VCC_net), .I0(n387), .I1(n558), .CO(n30868));
    SB_LUT4 rem_4_add_2055_28_lut (.I0(n3065), .I1(n3032), .I2(VCC_net), 
            .I3(n30867), .O(n3131)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_2055_27_lut (.I0(GND_net), .I1(n3033), .I2(VCC_net), 
            .I3(n30866), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_27 (.CI(n30866), .I0(n3033), .I1(VCC_net), 
            .CO(n30867));
    SB_LUT4 rem_4_add_2055_26_lut (.I0(GND_net), .I1(n3034), .I2(VCC_net), 
            .I3(n30865), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_26 (.CI(n30865), .I0(n3034), .I1(VCC_net), 
            .CO(n30866));
    SB_LUT4 rem_4_add_2055_25_lut (.I0(GND_net), .I1(n3035), .I2(VCC_net), 
            .I3(n30864), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_25 (.CI(n30864), .I0(n3035), .I1(VCC_net), 
            .CO(n30865));
    SB_LUT4 i37715_3_lut (.I0(n26_adj_4652), .I1(n95_adj_4360), .I2(n33_adj_4658), 
            .I3(GND_net), .O(n44840));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37715_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37716_3_lut (.I0(n44840), .I1(n94), .I2(n35_adj_4659), .I3(GND_net), 
            .O(n44841));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37716_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35900_4_lut (.I0(n39_adj_4662), .I1(n37_adj_4660), .I2(n35_adj_4659), 
            .I3(n43034), .O(n43024));
    defparam i35900_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37910_4_lut (.I0(n38_adj_4661), .I1(n28_adj_4654), .I2(n41_adj_4663), 
            .I3(n43022), .O(n45035));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37910_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i37533_3_lut (.I0(n44841), .I1(n93), .I2(n37_adj_4660), .I3(GND_net), 
            .O(n44658));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37533_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37983_4_lut (.I0(n44658), .I1(n45035), .I2(n41_adj_4663), 
            .I3(n43024), .O(n45108));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37983_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 rem_4_add_2055_24_lut (.I0(GND_net), .I1(n3036), .I2(VCC_net), 
            .I3(n30863), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_24 (.CI(n30863), .I0(n3036), .I1(VCC_net), 
            .CO(n30864));
    SB_LUT4 rem_4_add_2055_23_lut (.I0(GND_net), .I1(n3037), .I2(VCC_net), 
            .I3(n30862), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_23 (.CI(n30862), .I0(n3037), .I1(VCC_net), 
            .CO(n30863));
    SB_LUT4 rem_4_add_2055_22_lut (.I0(GND_net), .I1(n3038), .I2(VCC_net), 
            .I3(n30861), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_22 (.CI(n30861), .I0(n3038), .I1(VCC_net), 
            .CO(n30862));
    SB_LUT4 rem_4_add_2055_21_lut (.I0(GND_net), .I1(n3039), .I2(VCC_net), 
            .I3(n30860), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_21 (.CI(n30860), .I0(n3039), .I1(VCC_net), 
            .CO(n30861));
    SB_LUT4 rem_4_add_2055_20_lut (.I0(GND_net), .I1(n3040), .I2(VCC_net), 
            .I3(n30859), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_20 (.CI(n30859), .I0(n3040), .I1(VCC_net), 
            .CO(n30860));
    SB_LUT4 rem_4_add_2055_19_lut (.I0(GND_net), .I1(n3041), .I2(VCC_net), 
            .I3(n30858), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_19 (.CI(n30858), .I0(n3041), .I1(VCC_net), 
            .CO(n30859));
    SB_LUT4 rem_4_add_2055_18_lut (.I0(GND_net), .I1(n3042), .I2(VCC_net), 
            .I3(n30857), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_18 (.CI(n30857), .I0(n3042), .I1(VCC_net), 
            .CO(n30858));
    SB_LUT4 rem_4_add_2055_17_lut (.I0(GND_net), .I1(n3043), .I2(VCC_net), 
            .I3(n30856), .O(n3110)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_17 (.CI(n30856), .I0(n3043), .I1(VCC_net), 
            .CO(n30857));
    SB_LUT4 rem_4_add_2055_16_lut (.I0(GND_net), .I1(n3044), .I2(VCC_net), 
            .I3(n30855), .O(n3111)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_16 (.CI(n30855), .I0(n3044), .I1(VCC_net), 
            .CO(n30856));
    SB_LUT4 rem_4_add_2055_15_lut (.I0(GND_net), .I1(n3045), .I2(VCC_net), 
            .I3(n30854), .O(n3112)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_15 (.CI(n30854), .I0(n3045), .I1(VCC_net), 
            .CO(n30855));
    SB_LUT4 rem_4_add_2055_14_lut (.I0(GND_net), .I1(n3046), .I2(VCC_net), 
            .I3(n30853), .O(n3113)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_14 (.CI(n30853), .I0(n3046), .I1(VCC_net), 
            .CO(n30854));
    SB_LUT4 rem_4_add_2055_13_lut (.I0(GND_net), .I1(n3047), .I2(VCC_net), 
            .I3(n30852), .O(n3114)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_13 (.CI(n30852), .I0(n3047), .I1(VCC_net), 
            .CO(n30853));
    SB_LUT4 rem_4_add_2055_12_lut (.I0(GND_net), .I1(n3048), .I2(VCC_net), 
            .I3(n30851), .O(n3115)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_12 (.CI(n30851), .I0(n3048), .I1(VCC_net), 
            .CO(n30852));
    SB_LUT4 rem_4_add_2055_11_lut (.I0(GND_net), .I1(n3049), .I2(VCC_net), 
            .I3(n30850), .O(n3116)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_11 (.CI(n30850), .I0(n3049), .I1(VCC_net), 
            .CO(n30851));
    SB_LUT4 rem_4_add_2055_10_lut (.I0(GND_net), .I1(n3050), .I2(VCC_net), 
            .I3(n30849), .O(n3117)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_10 (.CI(n30849), .I0(n3050), .I1(VCC_net), 
            .CO(n30850));
    SB_LUT4 rem_4_add_2055_9_lut (.I0(GND_net), .I1(n3051), .I2(VCC_net), 
            .I3(n30848), .O(n3118)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_9 (.CI(n30848), .I0(n3051), .I1(VCC_net), 
            .CO(n30849));
    SB_LUT4 rem_4_add_2055_8_lut (.I0(GND_net), .I1(n3052), .I2(VCC_net), 
            .I3(n30847), .O(n3119)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_8 (.CI(n30847), .I0(n3052), .I1(VCC_net), 
            .CO(n30848));
    SB_LUT4 rem_4_add_2055_7_lut (.I0(GND_net), .I1(n3053), .I2(VCC_net), 
            .I3(n30846), .O(n3120)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_7 (.CI(n30846), .I0(n3053), .I1(VCC_net), 
            .CO(n30847));
    SB_LUT4 rem_4_add_2055_6_lut (.I0(GND_net), .I1(n3054), .I2(GND_net), 
            .I3(n30845), .O(n3121)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_6 (.CI(n30845), .I0(n3054), .I1(GND_net), 
            .CO(n30846));
    SB_LUT4 rem_4_add_2055_5_lut (.I0(GND_net), .I1(n3055), .I2(GND_net), 
            .I3(n30844), .O(n3122)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_5 (.CI(n30844), .I0(n3055), .I1(GND_net), 
            .CO(n30845));
    SB_LUT4 rem_4_add_2055_4_lut (.I0(GND_net), .I1(n3056), .I2(VCC_net), 
            .I3(n30843), .O(n3123)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_4 (.CI(n30843), .I0(n3056), .I1(VCC_net), 
            .CO(n30844));
    SB_LUT4 rem_4_add_2055_3_lut (.I0(GND_net), .I1(n3057), .I2(VCC_net), 
            .I3(n30842), .O(n3124)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_3 (.CI(n30842), .I0(n3057), .I1(VCC_net), 
            .CO(n30843));
    SB_LUT4 rem_4_add_2055_2_lut (.I0(GND_net), .I1(n3058), .I2(GND_net), 
            .I3(VCC_net), .O(n3125)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_2 (.CI(VCC_net), .I0(n3058), .I1(GND_net), 
            .CO(n30842));
    SB_LUT4 add_3162_20_lut (.I0(GND_net), .I1(n2357), .I2(n82), .I3(n30841), 
            .O(n7070)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3162_19_lut (.I0(GND_net), .I1(n2358), .I2(n83), .I3(n30840), 
            .O(n7071)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_19 (.CI(n30840), .I0(n2358), .I1(n83), .CO(n30841));
    SB_LUT4 add_3162_18_lut (.I0(GND_net), .I1(n2359), .I2(n84), .I3(n30839), 
            .O(n7072)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_18 (.CI(n30839), .I0(n2359), .I1(n84), .CO(n30840));
    SB_LUT4 add_3162_17_lut (.I0(GND_net), .I1(n2360), .I2(n85), .I3(n30838), 
            .O(n7073)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_17 (.CI(n30838), .I0(n2360), .I1(n85), .CO(n30839));
    SB_LUT4 add_3162_16_lut (.I0(GND_net), .I1(n2361), .I2(n86), .I3(n30837), 
            .O(n7074)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_16 (.CI(n30837), .I0(n2361), .I1(n86), .CO(n30838));
    SB_LUT4 add_3162_15_lut (.I0(GND_net), .I1(n2362), .I2(n87), .I3(n30836), 
            .O(n7075)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_15 (.CI(n30836), .I0(n2362), .I1(n87), .CO(n30837));
    SB_LUT4 add_3162_14_lut (.I0(GND_net), .I1(n2363), .I2(n88), .I3(n30835), 
            .O(n7076)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_14 (.CI(n30835), .I0(n2363), .I1(n88), .CO(n30836));
    SB_LUT4 add_3162_13_lut (.I0(GND_net), .I1(n2364), .I2(n89), .I3(n30834), 
            .O(n7077)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_13 (.CI(n30834), .I0(n2364), .I1(n89), .CO(n30835));
    SB_LUT4 add_3162_12_lut (.I0(GND_net), .I1(n2365), .I2(n90), .I3(n30833), 
            .O(n7078)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_12 (.CI(n30833), .I0(n2365), .I1(n90), .CO(n30834));
    SB_LUT4 add_3162_11_lut (.I0(GND_net), .I1(n2366), .I2(n91), .I3(n30832), 
            .O(n7079)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_11 (.CI(n30832), .I0(n2366), .I1(n91), .CO(n30833));
    SB_LUT4 add_3162_10_lut (.I0(GND_net), .I1(n2367), .I2(n92), .I3(n30831), 
            .O(n7080)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_10 (.CI(n30831), .I0(n2367), .I1(n92), .CO(n30832));
    SB_LUT4 add_3162_9_lut (.I0(GND_net), .I1(n2368), .I2(n93), .I3(n30830), 
            .O(n7081)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_9 (.CI(n30830), .I0(n2368), .I1(n93), .CO(n30831));
    SB_LUT4 add_3162_8_lut (.I0(GND_net), .I1(n2369), .I2(n94), .I3(n30829), 
            .O(n7082)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_8 (.CI(n30829), .I0(n2369), .I1(n94), .CO(n30830));
    SB_LUT4 add_3162_7_lut (.I0(GND_net), .I1(n2370), .I2(n95_adj_4360), 
            .I3(n30828), .O(n7083)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_7 (.CI(n30828), .I0(n2370), .I1(n95_adj_4360), .CO(n30829));
    SB_LUT4 add_3162_6_lut (.I0(GND_net), .I1(n2371), .I2(n96), .I3(n30827), 
            .O(n7084)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_6 (.CI(n30827), .I0(n2371), .I1(n96), .CO(n30828));
    SB_LUT4 add_3162_5_lut (.I0(GND_net), .I1(n2372), .I2(n97), .I3(n30826), 
            .O(n7085)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_5 (.CI(n30826), .I0(n2372), .I1(n97), .CO(n30827));
    SB_LUT4 add_3162_4_lut (.I0(GND_net), .I1(n2373), .I2(n98), .I3(n30825), 
            .O(n7086)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_4 (.CI(n30825), .I0(n2373), .I1(n98), .CO(n30826));
    SB_LUT4 add_3162_3_lut (.I0(GND_net), .I1(n2374), .I2(n99), .I3(n30824), 
            .O(n7087)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_3 (.CI(n30824), .I0(n2374), .I1(n99), .CO(n30825));
    SB_LUT4 add_3162_2_lut (.I0(GND_net), .I1(n386), .I2(n558), .I3(VCC_net), 
            .O(n7088)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3162_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3162_2 (.CI(VCC_net), .I0(n386), .I1(n558), .CO(n30824));
    SB_LUT4 add_3161_19_lut (.I0(GND_net), .I1(n2264), .I2(n83), .I3(n30823), 
            .O(n7050)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3161_18_lut (.I0(GND_net), .I1(n2265), .I2(n84), .I3(n30822), 
            .O(n7051)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_18 (.CI(n30822), .I0(n2265), .I1(n84), .CO(n30823));
    SB_LUT4 add_3161_17_lut (.I0(GND_net), .I1(n2266), .I2(n85), .I3(n30821), 
            .O(n7052)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_17 (.CI(n30821), .I0(n2266), .I1(n85), .CO(n30822));
    SB_LUT4 add_3161_16_lut (.I0(GND_net), .I1(n2267), .I2(n86), .I3(n30820), 
            .O(n7053)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_16 (.CI(n30820), .I0(n2267), .I1(n86), .CO(n30821));
    SB_LUT4 add_3161_15_lut (.I0(GND_net), .I1(n2268), .I2(n87), .I3(n30819), 
            .O(n7054)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_15 (.CI(n30819), .I0(n2268), .I1(n87), .CO(n30820));
    SB_LUT4 add_3161_14_lut (.I0(GND_net), .I1(n2269), .I2(n88), .I3(n30818), 
            .O(n7055)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_14 (.CI(n30818), .I0(n2269), .I1(n88), .CO(n30819));
    SB_LUT4 add_3161_13_lut (.I0(GND_net), .I1(n2270), .I2(n89), .I3(n30817), 
            .O(n7056)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_13 (.CI(n30817), .I0(n2270), .I1(n89), .CO(n30818));
    SB_LUT4 add_3161_12_lut (.I0(GND_net), .I1(n2271), .I2(n90), .I3(n30816), 
            .O(n7057)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_12 (.CI(n30816), .I0(n2271), .I1(n90), .CO(n30817));
    SB_LUT4 add_3161_11_lut (.I0(GND_net), .I1(n2272), .I2(n91), .I3(n30815), 
            .O(n7058)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_11 (.CI(n30815), .I0(n2272), .I1(n91), .CO(n30816));
    SB_LUT4 add_3161_10_lut (.I0(GND_net), .I1(n2273), .I2(n92), .I3(n30814), 
            .O(n7059)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_10 (.CI(n30814), .I0(n2273), .I1(n92), .CO(n30815));
    SB_LUT4 add_3161_9_lut (.I0(GND_net), .I1(n2274), .I2(n93), .I3(n30813), 
            .O(n7060)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_9 (.CI(n30813), .I0(n2274), .I1(n93), .CO(n30814));
    SB_LUT4 add_3161_8_lut (.I0(GND_net), .I1(n2275), .I2(n94), .I3(n30812), 
            .O(n7061)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_8 (.CI(n30812), .I0(n2275), .I1(n94), .CO(n30813));
    SB_LUT4 add_3161_7_lut (.I0(GND_net), .I1(n2276), .I2(n95_adj_4360), 
            .I3(n30811), .O(n7062)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_7 (.CI(n30811), .I0(n2276), .I1(n95_adj_4360), .CO(n30812));
    SB_LUT4 add_3161_6_lut (.I0(GND_net), .I1(n2277), .I2(n96), .I3(n30810), 
            .O(n7063)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_6 (.CI(n30810), .I0(n2277), .I1(n96), .CO(n30811));
    SB_LUT4 add_3161_5_lut (.I0(GND_net), .I1(n2278), .I2(n97), .I3(n30809), 
            .O(n7064)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_5 (.CI(n30809), .I0(n2278), .I1(n97), .CO(n30810));
    SB_LUT4 add_3161_4_lut (.I0(GND_net), .I1(n2279), .I2(n98), .I3(n30808), 
            .O(n7065)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_4 (.CI(n30808), .I0(n2279), .I1(n98), .CO(n30809));
    SB_LUT4 add_3161_3_lut (.I0(GND_net), .I1(n2280), .I2(n99), .I3(n30807), 
            .O(n7066)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_3 (.CI(n30807), .I0(n2280), .I1(n99), .CO(n30808));
    SB_LUT4 add_3161_2_lut (.I0(GND_net), .I1(n385), .I2(n558), .I3(VCC_net), 
            .O(n7067)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3161_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3161_2 (.CI(VCC_net), .I0(n385), .I1(n558), .CO(n30807));
    SB_LUT4 add_3160_18_lut (.I0(GND_net), .I1(n2168), .I2(n84), .I3(n30806), 
            .O(n7031)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3160_17_lut (.I0(GND_net), .I1(n2169), .I2(n85), .I3(n30805), 
            .O(n7032)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3160_17 (.CI(n30805), .I0(n2169), .I1(n85), .CO(n30806));
    SB_LUT4 add_3160_16_lut (.I0(GND_net), .I1(n2170), .I2(n86), .I3(n30804), 
            .O(n7033)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3160_16 (.CI(n30804), .I0(n2170), .I1(n86), .CO(n30805));
    SB_LUT4 add_3160_15_lut (.I0(GND_net), .I1(n2171), .I2(n87), .I3(n30803), 
            .O(n7034)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3160_15 (.CI(n30803), .I0(n2171), .I1(n87), .CO(n30804));
    SB_LUT4 add_3160_14_lut (.I0(GND_net), .I1(n2172), .I2(n88), .I3(n30802), 
            .O(n7035)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3160_14 (.CI(n30802), .I0(n2172), .I1(n88), .CO(n30803));
    SB_LUT4 add_3160_13_lut (.I0(GND_net), .I1(n2173), .I2(n89), .I3(n30801), 
            .O(n7036)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3160_13 (.CI(n30801), .I0(n2173), .I1(n89), .CO(n30802));
    SB_LUT4 add_3160_12_lut (.I0(GND_net), .I1(n2174), .I2(n90), .I3(n30800), 
            .O(n7037)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3160_12 (.CI(n30800), .I0(n2174), .I1(n90), .CO(n30801));
    SB_LUT4 add_3160_11_lut (.I0(GND_net), .I1(n2175), .I2(n91), .I3(n30799), 
            .O(n7038)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3160_11 (.CI(n30799), .I0(n2175), .I1(n91), .CO(n30800));
    SB_LUT4 add_3160_10_lut (.I0(GND_net), .I1(n2176), .I2(n92), .I3(n30798), 
            .O(n7039)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3160_10 (.CI(n30798), .I0(n2176), .I1(n92), .CO(n30799));
    SB_LUT4 add_3160_9_lut (.I0(GND_net), .I1(n2177), .I2(n93), .I3(n30797), 
            .O(n7040)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3160_9 (.CI(n30797), .I0(n2177), .I1(n93), .CO(n30798));
    SB_LUT4 add_3160_8_lut (.I0(GND_net), .I1(n2178), .I2(n94), .I3(n30796), 
            .O(n7041)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3160_8 (.CI(n30796), .I0(n2178), .I1(n94), .CO(n30797));
    SB_LUT4 i37984_3_lut (.I0(n45108), .I1(n90), .I2(n1756), .I3(GND_net), 
            .O(n45109));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37984_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i37964_3_lut (.I0(n45109), .I1(n89), .I2(n1755), .I3(GND_net), 
            .O(n45089));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37964_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 rem_4_i1731_3_lut (.I0(n2546_adj_4516), .I1(n2613), .I2(n2570), 
            .I3(GND_net), .O(n2645));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1704 (.I0(n45089), .I1(n17299), .I2(n88), .I3(n1754), 
            .O(n1778));
    defparam i1_4_lut_adj_1704.LUT_INIT = 16'hceef;
    SB_LUT4 div_36_LessThan_1062_i39_2_lut (.I0(n1647), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4648));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1062_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1062_i37_2_lut (.I0(n1648), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4647));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1062_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_mux_3_i13_3_lut (.I0(encoder0_position[12]), .I1(n13_adj_4375), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n379));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1062_i43_2_lut (.I0(n1645), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4651));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1062_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1062_i41_2_lut (.I0(n1646), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4650));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1062_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1062_i31_2_lut (.I0(n1651), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4643));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1062_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1062_i33_2_lut (.I0(n1650), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4645));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1062_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1062_i35_2_lut (.I0(n1649), .I1(n95_adj_4360), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4646));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1062_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_i1064_1_lut (.I0(n1667), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1668));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1064_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_1062_i29_2_lut (.I0(n1652), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4641));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1062_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i35932_4_lut (.I0(n35_adj_4646), .I1(n33_adj_4645), .I2(n31_adj_4643), 
            .I3(n29_adj_4641), .O(n43056));
    defparam i35932_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_36_LessThan_1062_i40_3_lut (.I0(n32_adj_4644), .I1(n91), 
            .I2(n43_adj_4651), .I3(GND_net), .O(n40_adj_4649));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1062_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_36_LessThan_1062_i28_4_lut (.I0(n379), .I1(n99), .I2(n1653), 
            .I3(n558), .O(n28_adj_4640));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1062_i28_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i37721_3_lut (.I0(n28_adj_4640), .I1(n95_adj_4360), .I2(n35_adj_4646), 
            .I3(GND_net), .O(n44846));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37721_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3160_7_lut (.I0(GND_net), .I1(n2179), .I2(n95_adj_4360), 
            .I3(n30795), .O(n7042)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_unary_minus_4_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4534), .I3(n31237), .O(n65)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_4_add_3_12 (.CI(n31237), .I0(GND_net), .I1(n15_adj_4534), 
            .CO(n31238));
    SB_LUT4 i37722_3_lut (.I0(n44846), .I1(n94), .I2(n37_adj_4647), .I3(GND_net), 
            .O(n44847));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37722_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_36_unary_minus_4_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4535), .I3(n31236), .O(n66)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35924_4_lut (.I0(n41_adj_4650), .I1(n39_adj_4648), .I2(n37_adj_4647), 
            .I3(n43056), .O(n43048));
    defparam i35924_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_3160_7 (.CI(n30795), .I0(n2179), .I1(n95_adj_4360), .CO(n30796));
    SB_LUT4 add_3160_6_lut (.I0(GND_net), .I1(n2180), .I2(n96), .I3(n30794), 
            .O(n7043)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37719_4_lut (.I0(n40_adj_4649), .I1(n30_adj_4642), .I2(n43_adj_4651), 
            .I3(n43044), .O(n44844));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37719_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY div_36_unary_minus_4_add_3_11 (.CI(n31236), .I0(GND_net), .I1(n16_adj_4535), 
            .CO(n31237));
    SB_CARRY add_3160_6 (.CI(n30794), .I0(n2180), .I1(n96), .CO(n30795));
    SB_LUT4 i37529_3_lut (.I0(n44847), .I1(n93), .I2(n39_adj_4648), .I3(GND_net), 
            .O(n44654));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37529_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3160_5_lut (.I0(GND_net), .I1(n2181), .I2(n97), .I3(n30793), 
            .O(n7044)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_unary_minus_4_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4536), .I3(n31235), .O(n67)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_4_add_3_10 (.CI(n31235), .I0(GND_net), .I1(n17_adj_4536), 
            .CO(n31236));
    SB_LUT4 add_553_19_lut (.I0(duty[17]), .I1(n45865), .I2(n8), .I3(n30449), 
            .O(pwm_setpoint_22__N_57[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i37903_4_lut (.I0(n44654), .I1(n44844), .I2(n43_adj_4651), 
            .I3(n43048), .O(n45028));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37903_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_3160_5 (.CI(n30793), .I0(n2181), .I1(n97), .CO(n30794));
    SB_LUT4 add_3160_4_lut (.I0(GND_net), .I1(n2182), .I2(n98), .I3(n30792), 
            .O(n7045)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_unary_minus_4_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4537), .I3(n31234), .O(n68)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3160_4 (.CI(n30792), .I0(n2182), .I1(n98), .CO(n30793));
    SB_CARRY div_36_unary_minus_4_add_3_9 (.CI(n31234), .I0(GND_net), .I1(n18_adj_4537), 
            .CO(n31235));
    SB_LUT4 i37904_3_lut (.I0(n45028), .I1(n90), .I2(n1644), .I3(GND_net), 
            .O(n45029));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37904_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 add_3160_3_lut (.I0(GND_net), .I1(n2183), .I2(n99), .I3(n30791), 
            .O(n7046)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1705 (.I0(n45029), .I1(n17296), .I2(n89), .I3(n1643), 
            .O(n1667));
    defparam i1_4_lut_adj_1705.LUT_INIT = 16'hceef;
    SB_CARRY add_3160_3 (.CI(n30791), .I0(n2183), .I1(n99), .CO(n30792));
    SB_CARRY add_553_19 (.CI(n30449), .I0(n45865), .I1(n8), .CO(n30450));
    SB_LUT4 div_36_unary_minus_4_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4538), .I3(n31233), .O(n69)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_4_add_3_8 (.CI(n31233), .I0(GND_net), .I1(n19_adj_4538), 
            .CO(n31234));
    SB_LUT4 div_36_LessThan_985_i41_2_lut (.I0(n1532), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4636));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_985_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_985_i39_2_lut (.I0(n1533), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4635));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_985_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_mux_3_i14_3_lut (.I0(encoder0_position[13]), .I1(n12_adj_4366), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n378));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_985_i45_2_lut (.I0(n1530), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4639));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_985_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3160_2_lut (.I0(GND_net), .I1(n384), .I2(n558), .I3(VCC_net), 
            .O(n7047)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3160_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_985_i35_2_lut (.I0(n1535), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4633));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_985_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_unary_minus_4_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4539), .I3(n31232), .O(n70)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_985_i37_2_lut (.I0(n1534), .I1(n95_adj_4360), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4634));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_985_i37_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3160_2 (.CI(VCC_net), .I0(n384), .I1(n558), .CO(n30791));
    SB_LUT4 add_3159_17_lut (.I0(GND_net), .I1(n2069), .I2(n85), .I3(n30790), 
            .O(n7013)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3159_16_lut (.I0(GND_net), .I1(n2070), .I2(n86), .I3(n30789), 
            .O(n7014)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3159_16 (.CI(n30789), .I0(n2070), .I1(n86), .CO(n30790));
    SB_LUT4 add_3159_15_lut (.I0(GND_net), .I1(n2071), .I2(n87), .I3(n30788), 
            .O(n7015)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_985_i33_2_lut (.I0(n1536), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4631));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_985_i33_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_3159_15 (.CI(n30788), .I0(n2071), .I1(n87), .CO(n30789));
    SB_LUT4 add_3159_14_lut (.I0(GND_net), .I1(n2072), .I2(n88), .I3(n30787), 
            .O(n7016)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3159_14 (.CI(n30787), .I0(n2072), .I1(n88), .CO(n30788));
    SB_LUT4 add_3159_13_lut (.I0(GND_net), .I1(n2073), .I2(n89), .I3(n30786), 
            .O(n7017)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3159_13 (.CI(n30786), .I0(n2073), .I1(n89), .CO(n30787));
    SB_LUT4 div_36_LessThan_985_i43_2_lut (.I0(n1531), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4638));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_985_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3159_12_lut (.I0(GND_net), .I1(n2074), .I2(n90), .I3(n30785), 
            .O(n7018)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_4_add_3_7 (.CI(n31232), .I0(GND_net), .I1(n20_adj_4539), 
            .CO(n31233));
    SB_LUT4 add_553_18_lut (.I0(duty[16]), .I1(n45865), .I2(n9), .I3(n30448), 
            .O(pwm_setpoint_22__N_57[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3159_12 (.CI(n30785), .I0(n2074), .I1(n90), .CO(n30786));
    SB_LUT4 div_36_unary_minus_4_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4540), .I3(n31231), .O(n71)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i987_1_lut (.I0(n1553), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1554));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i987_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_985_i31_2_lut (.I0(n1537), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4629));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_985_i31_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY div_36_unary_minus_4_add_3_6 (.CI(n31231), .I0(GND_net), .I1(n21_adj_4540), 
            .CO(n31232));
    SB_LUT4 i35968_4_lut (.I0(n37_adj_4634), .I1(n35_adj_4633), .I2(n33_adj_4631), 
            .I3(n31_adj_4629), .O(n43092));
    defparam i35968_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3159_11_lut (.I0(GND_net), .I1(n2075), .I2(n91), .I3(n30784), 
            .O(n7019)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_unary_minus_4_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4541), .I3(n31230), .O(n72)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_36_unary_minus_4_add_3_5 (.CI(n31230), .I0(GND_net), .I1(n22_adj_4541), 
            .CO(n31231));
    SB_LUT4 div_36_LessThan_985_i42_3_lut (.I0(n34_adj_4632), .I1(n91), 
            .I2(n45_adj_4639), .I3(GND_net), .O(n42_adj_4637));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_985_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_36_LessThan_985_i30_4_lut (.I0(n378), .I1(n99), .I2(n1538), 
            .I3(n558), .O(n30_adj_4628));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_985_i30_4_lut.LUT_INIT = 16'h0317;
    SB_CARRY add_3159_11 (.CI(n30784), .I0(n2075), .I1(n91), .CO(n30785));
    SB_LUT4 div_36_unary_minus_4_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4542), .I3(n31229), .O(n73)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_553_18 (.CI(n30448), .I0(n45865), .I1(n9), .CO(n30449));
    SB_LUT4 i37725_3_lut (.I0(n30_adj_4628), .I1(n95_adj_4360), .I2(n37_adj_4634), 
            .I3(GND_net), .O(n44850));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37725_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3159_10_lut (.I0(GND_net), .I1(n2076), .I2(n92), .I3(n30783), 
            .O(n7020)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3159_10 (.CI(n30783), .I0(n2076), .I1(n92), .CO(n30784));
    SB_LUT4 add_3159_9_lut (.I0(GND_net), .I1(n2077), .I2(n93), .I3(n30782), 
            .O(n7021)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3159_9 (.CI(n30782), .I0(n2077), .I1(n93), .CO(n30783));
    SB_LUT4 add_3159_8_lut (.I0(GND_net), .I1(n2078), .I2(n94), .I3(n30781), 
            .O(n7022)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37726_3_lut (.I0(n44850), .I1(n94), .I2(n39_adj_4635), .I3(GND_net), 
            .O(n44851));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37726_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35960_4_lut (.I0(n43_adj_4638), .I1(n41_adj_4636), .I2(n39_adj_4635), 
            .I3(n43092), .O(n43084));
    defparam i35960_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37272_4_lut (.I0(n42_adj_4637), .I1(n32_adj_4630), .I2(n45_adj_4639), 
            .I3(n43070), .O(n44397));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37272_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i37523_3_lut (.I0(n44851), .I1(n93), .I2(n41_adj_4636), .I3(GND_net), 
            .O(n44648));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37523_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_3159_8 (.CI(n30781), .I0(n2078), .I1(n94), .CO(n30782));
    SB_CARRY div_36_unary_minus_4_add_3_4 (.CI(n31229), .I0(GND_net), .I1(n23_adj_4542), 
            .CO(n31230));
    SB_LUT4 div_36_unary_minus_4_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4543), .I3(n31228), .O(n74)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37741_4_lut (.I0(n44648), .I1(n44397), .I2(n45_adj_4639), 
            .I3(n43084), .O(n44866));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37741_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1706 (.I0(n44866), .I1(n17293), .I2(n90), .I3(n1529), 
            .O(n1553));
    defparam i1_4_lut_adj_1706.LUT_INIT = 16'hceef;
    SB_LUT4 rem_4_i1743_3_lut (.I0(n2558_adj_4508), .I1(n2625_adj_4500), 
            .I2(n2570), .I3(GND_net), .O(n2657));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_906_i43_2_lut (.I0(n1414), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4625));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_906_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_3159_7_lut (.I0(GND_net), .I1(n2079), .I2(n95_adj_4360), 
            .I3(n30780), .O(n7023)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3159_7 (.CI(n30780), .I0(n2079), .I1(n95_adj_4360), .CO(n30781));
    SB_LUT4 rem_4_i1741_3_lut (.I0(n2556), .I1(n2623_adj_4503), .I2(n2570), 
            .I3(GND_net), .O(n2655));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1741_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_906_i37_2_lut (.I0(n1417), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4622));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_906_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_906_i41_2_lut (.I0(n1415), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4624));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_906_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_906_i39_2_lut (.I0(n1416), .I1(n95_adj_4360), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4623));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_906_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_mux_3_i15_3_lut (.I0(encoder0_position[14]), .I1(n11_adj_4382), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n377));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_36_unary_minus_4_add_3_3 (.CI(n31228), .I0(GND_net), .I1(n24_adj_4543), 
            .CO(n31229));
    SB_LUT4 add_3159_6_lut (.I0(GND_net), .I1(n2080), .I2(n96), .I3(n30779), 
            .O(n7024)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3159_6 (.CI(n30779), .I0(n2080), .I1(n96), .CO(n30780));
    SB_LUT4 div_36_i908_1_lut (.I0(n1436), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1437));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i908_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3159_5_lut (.I0(GND_net), .I1(n2081), .I2(n97), .I3(n30778), 
            .O(n7025)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3159_5 (.CI(n30778), .I0(n2081), .I1(n97), .CO(n30779));
    SB_LUT4 div_36_LessThan_906_i32_4_lut (.I0(n377), .I1(n99), .I2(n1420), 
            .I3(n558), .O(n32_adj_4620));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_906_i32_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 add_3159_4_lut (.I0(GND_net), .I1(n2082), .I2(n98), .I3(n30777), 
            .O(n7026)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_unary_minus_4_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4544), .I3(VCC_net), .O(n75)) /* synthesis syn_instantiated=1 */ ;
    defparam div_36_unary_minus_4_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3159_4 (.CI(n30777), .I0(n2082), .I1(n98), .CO(n30778));
    SB_LUT4 add_553_17_lut (.I0(duty[15]), .I1(n45865), .I2(n10_adj_4330), 
            .I3(n30447), .O(pwm_setpoint_22__N_57[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i37731_3_lut (.I0(n32_adj_4620), .I1(n95_adj_4360), .I2(n39_adj_4623), 
            .I3(GND_net), .O(n44856));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37731_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_3159_3_lut (.I0(GND_net), .I1(n2083), .I2(n99), .I3(n30776), 
            .O(n7027)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37732_3_lut (.I0(n44856), .I1(n94), .I2(n41_adj_4624), .I3(GND_net), 
            .O(n44857));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37732_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36710_4_lut (.I0(n41_adj_4624), .I1(n39_adj_4623), .I2(n37_adj_4622), 
            .I3(n43128), .O(n43835));
    defparam i36710_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i37270_3_lut (.I0(n34_adj_4621), .I1(n96), .I2(n37_adj_4622), 
            .I3(GND_net), .O(n44395));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37270_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37519_3_lut (.I0(n44857), .I1(n93), .I2(n43_adj_4625), .I3(GND_net), 
            .O(n44644));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37519_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37729_4_lut (.I0(n44644), .I1(n44395), .I2(n43_adj_4625), 
            .I3(n43835), .O(n44854));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37729_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i37730_3_lut (.I0(n44854), .I1(n92), .I2(n1413), .I3(GND_net), 
            .O(n44855));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37730_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1707 (.I0(n44855), .I1(n17211), .I2(n91), .I3(n1412), 
            .O(n1436));
    defparam i1_4_lut_adj_1707.LUT_INIT = 16'hceef;
    SB_LUT4 div_36_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4562));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_825_i45_2_lut (.I0(n1293), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4617));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_825_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i1740_3_lut (.I0(n2555), .I1(n2622_adj_4505), .I2(n2570), 
            .I3(GND_net), .O(n2654));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_825_i39_2_lut (.I0(n1296), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4613));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_825_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_825_i43_2_lut (.I0(n1294), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4615));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_825_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_825_i41_2_lut (.I0(n1295), .I1(n95_adj_4360), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4614));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_825_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_mux_3_i16_3_lut (.I0(encoder0_position[15]), .I1(n10), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n376));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_36_unary_minus_4_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4544), 
            .CO(n31228));
    SB_CARRY add_553_17 (.CI(n30447), .I0(n45865), .I1(n10_adj_4330), 
            .CO(n30448));
    SB_LUT4 add_553_16_lut (.I0(duty[14]), .I1(n45865), .I2(n11), .I3(n30446), 
            .O(pwm_setpoint_22__N_57[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1586_22_lut (.I0(n2372_adj_4587), .I1(n2339), .I2(VCC_net), 
            .I3(n31227), .O(n2438)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1586_21_lut (.I0(GND_net), .I1(n2340), .I2(VCC_net), 
            .I3(n31226), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3159_3 (.CI(n30776), .I0(n2083), .I1(n99), .CO(n30777));
    SB_CARRY rem_4_add_1586_21 (.CI(n31226), .I0(n2340), .I1(VCC_net), 
            .CO(n31227));
    SB_LUT4 div_36_i827_1_lut (.I0(n1316), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1317));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i827_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_1586_20_lut (.I0(GND_net), .I1(n2341), .I2(VCC_net), 
            .I3(n31225), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_20 (.CI(n31225), .I0(n2341), .I1(VCC_net), 
            .CO(n31226));
    SB_LUT4 rem_4_add_1586_19_lut (.I0(GND_net), .I1(n2342), .I2(VCC_net), 
            .I3(n31224), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3159_2_lut (.I0(GND_net), .I1(n383), .I2(n558), .I3(VCC_net), 
            .O(n7028)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3159_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3159_2 (.CI(VCC_net), .I0(n383), .I1(n558), .CO(n30776));
    SB_CARRY rem_4_add_1586_19 (.CI(n31224), .I0(n2342), .I1(VCC_net), 
            .CO(n31225));
    SB_LUT4 div_36_i723_3_lut_3_lut (.I0(n1067), .I1(n6899), .I2(n1047), 
            .I3(GND_net), .O(n1173));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i723_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_2122_29_lut (.I0(n3164), .I1(n3131), .I2(VCC_net), 
            .I3(n30775), .O(n3230)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_36_i722_3_lut_3_lut (.I0(n1067), .I1(n6898), .I2(n1046), 
            .I3(GND_net), .O(n1172));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i722_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1742_3_lut (.I0(n2557), .I1(n2624_adj_4501), .I2(n2570), 
            .I3(GND_net), .O(n2656));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1742_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1723_3_lut (.I0(n2538_adj_4572), .I1(n2605), .I2(n2570), 
            .I3(GND_net), .O(n2637_adj_4492));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_825_i34_4_lut (.I0(n376), .I1(n99), .I2(n1299), 
            .I3(n558), .O(n34_adj_4610));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_825_i34_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 rem_4_add_2122_28_lut (.I0(GND_net), .I1(n3132), .I2(VCC_net), 
            .I3(n30774), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_553_16 (.CI(n30446), .I0(n45865), .I1(n11), .CO(n30447));
    SB_CARRY rem_4_add_2122_28 (.CI(n30774), .I0(n3132), .I1(VCC_net), 
            .CO(n30775));
    SB_LUT4 rem_4_add_2122_27_lut (.I0(GND_net), .I1(n3133), .I2(VCC_net), 
            .I3(n30773), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_18_lut (.I0(GND_net), .I1(n2343), .I2(VCC_net), 
            .I3(n31223), .O(n2410)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_27 (.CI(n30773), .I0(n3133), .I1(VCC_net), 
            .CO(n30774));
    SB_LUT4 rem_4_add_2122_26_lut (.I0(GND_net), .I1(n3134), .I2(VCC_net), 
            .I3(n30772), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i724_3_lut_3_lut (.I0(n1067), .I1(n6900), .I2(n1048), 
            .I3(GND_net), .O(n1174));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i724_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_DFF communication_counter_1146__i2 (.Q(communication_counter[2]), .C(LED_c), 
           .D(n163));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_LUT4 i37733_3_lut (.I0(n34_adj_4610), .I1(n95_adj_4360), .I2(n41_adj_4614), 
            .I3(GND_net), .O(n44858));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37733_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_1586_18 (.CI(n31223), .I0(n2343), .I1(VCC_net), 
            .CO(n31224));
    SB_LUT4 rem_4_add_1586_17_lut (.I0(GND_net), .I1(n2344), .I2(VCC_net), 
            .I3(n31222), .O(n2411)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_26 (.CI(n30772), .I0(n3134), .I1(VCC_net), 
            .CO(n30773));
    SB_LUT4 add_553_15_lut (.I0(duty[13]), .I1(n45865), .I2(n12), .I3(n30445), 
            .O(pwm_setpoint_22__N_57[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i37734_3_lut (.I0(n44858), .I1(n94), .I2(n43_adj_4615), .I3(GND_net), 
            .O(n44859));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37734_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_add_2122_25_lut (.I0(GND_net), .I1(n3135), .I2(VCC_net), 
            .I3(n30771), .O(n3202)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_25 (.CI(n30771), .I0(n3135), .I1(VCC_net), 
            .CO(n30772));
    SB_CARRY rem_4_add_1586_17 (.CI(n31222), .I0(n2344), .I1(VCC_net), 
            .CO(n31223));
    SB_LUT4 rem_4_add_1586_16_lut (.I0(GND_net), .I1(n2345), .I2(VCC_net), 
            .I3(n31221), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_24_lut (.I0(GND_net), .I1(n3136), .I2(VCC_net), 
            .I3(n30770), .O(n3203)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_16 (.CI(n31221), .I0(n2345), .I1(VCC_net), 
            .CO(n31222));
    SB_LUT4 rem_4_add_1586_15_lut (.I0(GND_net), .I1(n2346), .I2(VCC_net), 
            .I3(n31220), .O(n2413)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_15 (.CI(n31220), .I0(n2346), .I1(VCC_net), 
            .CO(n31221));
    SB_CARRY rem_4_add_2122_24 (.CI(n30770), .I0(n3136), .I1(VCC_net), 
            .CO(n30771));
    SB_LUT4 rem_4_i1739_3_lut (.I0(n2554), .I1(n2621_adj_4504), .I2(n2570), 
            .I3(GND_net), .O(n2653));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1739_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2122_23_lut (.I0(GND_net), .I1(n3137), .I2(VCC_net), 
            .I3(n30769), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_14_lut (.I0(GND_net), .I1(n2347), .I2(VCC_net), 
            .I3(n31219), .O(n2414)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_23 (.CI(n30769), .I0(n3137), .I1(VCC_net), 
            .CO(n30770));
    SB_LUT4 rem_4_add_2122_22_lut (.I0(GND_net), .I1(n3138), .I2(VCC_net), 
            .I3(n30768), .O(n3205)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36722_4_lut (.I0(n43_adj_4615), .I1(n41_adj_4614), .I2(n39_adj_4613), 
            .I3(n43164), .O(n43847));
    defparam i36722_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_36_LessThan_825_i38_3_lut (.I0(n36_adj_4611), .I1(n96), 
            .I2(n39_adj_4613), .I3(GND_net), .O(n38_adj_4612));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_825_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37513_3_lut (.I0(n44859), .I1(n93), .I2(n45_adj_4617), .I3(GND_net), 
            .O(n44_adj_4616));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37513_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFF communication_counter_1146__i3 (.Q(communication_counter[3]), .C(LED_c), 
           .D(n162));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i4 (.Q(communication_counter[4]), .C(LED_c), 
           .D(n161));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i5 (.Q(communication_counter[5]), .C(LED_c), 
           .D(n160));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i6 (.Q(communication_counter[6]), .C(LED_c), 
           .D(n159));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i7 (.Q(communication_counter[7]), .C(LED_c), 
           .D(n158));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i8 (.Q(communication_counter[8]), .C(LED_c), 
           .D(n157));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i9 (.Q(communication_counter[9]), .C(LED_c), 
           .D(n156));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i10 (.Q(communication_counter[10]), 
           .C(LED_c), .D(n155));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i11 (.Q(communication_counter[11]), 
           .C(LED_c), .D(n154));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i12 (.Q(communication_counter[12]), 
           .C(LED_c), .D(n153));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i13 (.Q(communication_counter[13]), 
           .C(LED_c), .D(n152));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i14 (.Q(communication_counter[14]), 
           .C(LED_c), .D(n151));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i15 (.Q(communication_counter[15]), 
           .C(LED_c), .D(n150));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i16 (.Q(communication_counter[16]), 
           .C(LED_c), .D(n149));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i17 (.Q(communication_counter[17]), 
           .C(LED_c), .D(n148));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i18 (.Q(communication_counter[18]), 
           .C(LED_c), .D(n147));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i19 (.Q(communication_counter[19]), 
           .C(LED_c), .D(n146));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i20 (.Q(communication_counter[20]), 
           .C(LED_c), .D(n145));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i21 (.Q(communication_counter[21]), 
           .C(LED_c), .D(n144));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i22 (.Q(communication_counter[22]), 
           .C(LED_c), .D(n143));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i23 (.Q(communication_counter[23]), 
           .C(LED_c), .D(n142));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i24 (.Q(communication_counter[24]), 
           .C(LED_c), .D(n141));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i25 (.Q(communication_counter[25]), 
           .C(LED_c), .D(n140));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i26 (.Q(communication_counter[26]), 
           .C(LED_c), .D(n139));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i27 (.Q(communication_counter[27]), 
           .C(LED_c), .D(n138));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i28 (.Q(communication_counter[28]), 
           .C(LED_c), .D(n137));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i29 (.Q(communication_counter[29]), 
           .C(LED_c), .D(n136));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i30 (.Q(communication_counter[30]), 
           .C(LED_c), .D(n135));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_DFF communication_counter_1146__i31 (.Q(communication_counter[31]), 
           .C(LED_c), .D(n134));   // verilog/TinyFPGA_B.v(49[28:51])
    SB_CARRY add_553_15 (.CI(n30445), .I0(n45865), .I1(n12), .CO(n30446));
    SB_CARRY rem_4_add_2122_22 (.CI(n30768), .I0(n3138), .I1(VCC_net), 
            .CO(n30769));
    SB_LUT4 rem_4_add_2122_21_lut (.I0(GND_net), .I1(n3139), .I2(VCC_net), 
            .I3(n30767), .O(n3206)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_14 (.CI(n31219), .I0(n2347), .I1(VCC_net), 
            .CO(n31220));
    SB_LUT4 rem_4_add_1586_13_lut (.I0(GND_net), .I1(n2348), .I2(VCC_net), 
            .I3(n31218), .O(n2415)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_21 (.CI(n30767), .I0(n3139), .I1(VCC_net), 
            .CO(n30768));
    SB_CARRY rem_4_add_1586_13 (.CI(n31218), .I0(n2348), .I1(VCC_net), 
            .CO(n31219));
    SB_LUT4 rem_4_add_2122_20_lut (.I0(GND_net), .I1(n3140), .I2(VCC_net), 
            .I3(n30766), .O(n3207)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_20 (.CI(n30766), .I0(n3140), .I1(VCC_net), 
            .CO(n30767));
    SB_LUT4 rem_4_add_2122_19_lut (.I0(GND_net), .I1(n3141), .I2(VCC_net), 
            .I3(n30765), .O(n3208)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_19 (.CI(n30765), .I0(n3141), .I1(VCC_net), 
            .CO(n30766));
    SB_LUT4 rem_4_add_2122_18_lut (.I0(GND_net), .I1(n3142), .I2(VCC_net), 
            .I3(n30764), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_553_14_lut (.I0(duty[12]), .I1(n45865), .I2(n13_adj_4331), 
            .I3(n30444), .O(pwm_setpoint_22__N_57[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2122_18 (.CI(n30764), .I0(n3142), .I1(VCC_net), 
            .CO(n30765));
    SB_LUT4 rem_4_add_2122_17_lut (.I0(GND_net), .I1(n3143), .I2(VCC_net), 
            .I3(n30763), .O(n3210)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_17 (.CI(n30763), .I0(n3143), .I1(VCC_net), 
            .CO(n30764));
    SB_LUT4 div_36_i725_3_lut_3_lut (.I0(n1067), .I1(n6901), .I2(n374), 
            .I3(GND_net), .O(n1175));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i725_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i721_3_lut_3_lut (.I0(n1067), .I1(n6897), .I2(n1045), 
            .I3(GND_net), .O(n1171));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i721_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i719_3_lut_3_lut (.I0(n1067), .I1(n6895), .I2(n1043), 
            .I3(GND_net), .O(n1169));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_2122_16_lut (.I0(GND_net), .I1(n3144), .I2(VCC_net), 
            .I3(n30762), .O(n3211)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_16 (.CI(n30762), .I0(n3144), .I1(VCC_net), 
            .CO(n30763));
    SB_LUT4 rem_4_add_2122_15_lut (.I0(GND_net), .I1(n3145), .I2(VCC_net), 
            .I3(n30761), .O(n3212)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_15 (.CI(n30761), .I0(n3145), .I1(VCC_net), 
            .CO(n30762));
    SB_LUT4 rem_4_add_2122_14_lut (.I0(GND_net), .I1(n3146), .I2(VCC_net), 
            .I3(n30760), .O(n3213)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37268_4_lut (.I0(n44_adj_4616), .I1(n38_adj_4612), .I2(n45_adj_4617), 
            .I3(n43847), .O(n44393));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37268_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_553_14 (.CI(n30444), .I0(n45865), .I1(n13_adj_4331), 
            .CO(n30445));
    SB_CARRY rem_4_add_2122_14 (.CI(n30760), .I0(n3146), .I1(VCC_net), 
            .CO(n30761));
    SB_LUT4 rem_4_add_1586_12_lut (.I0(GND_net), .I1(n2349), .I2(VCC_net), 
            .I3(n31217), .O(n2416)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_13_lut (.I0(GND_net), .I1(n3147), .I2(VCC_net), 
            .I3(n30759), .O(n3214)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_13 (.CI(n30759), .I0(n3147), .I1(VCC_net), 
            .CO(n30760));
    SB_CARRY rem_4_add_1586_12 (.CI(n31217), .I0(n2349), .I1(VCC_net), 
            .CO(n31218));
    SB_LUT4 i1_4_lut_adj_1708 (.I0(n44393), .I1(n17290), .I2(n92), .I3(n1292), 
            .O(n1316));
    defparam i1_4_lut_adj_1708.LUT_INIT = 16'hceef;
    SB_LUT4 rem_4_add_1586_11_lut (.I0(GND_net), .I1(n2350), .I2(VCC_net), 
            .I3(n31216), .O(n2417)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_12_lut (.I0(GND_net), .I1(n3148), .I2(VCC_net), 
            .I3(n30758), .O(n3215)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i720_3_lut_3_lut (.I0(n1067), .I1(n6896), .I2(n1044), 
            .I3(GND_net), .O(n1170));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i720_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_2122_12 (.CI(n30758), .I0(n3148), .I1(VCC_net), 
            .CO(n30759));
    SB_LUT4 add_553_13_lut (.I0(duty[11]), .I1(n45865), .I2(n14_adj_4332), 
            .I3(n30443), .O(pwm_setpoint_22__N_57[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_13_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_36_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4561));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1586_11 (.CI(n31216), .I0(n2350), .I1(VCC_net), 
            .CO(n31217));
    SB_LUT4 rem_4_add_1586_10_lut (.I0(GND_net), .I1(n2351), .I2(VCC_net), 
            .I3(n31215), .O(n2418)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_11_lut (.I0(GND_net), .I1(n3149), .I2(VCC_net), 
            .I3(n30757), .O(n3216)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_11 (.CI(n30757), .I0(n3149), .I1(VCC_net), 
            .CO(n30758));
    SB_LUT4 rem_4_add_2122_10_lut (.I0(GND_net), .I1(n3150), .I2(VCC_net), 
            .I3(n30756), .O(n3217)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_10 (.CI(n31215), .I0(n2351), .I1(VCC_net), 
            .CO(n31216));
    SB_CARRY rem_4_add_2122_10 (.CI(n30756), .I0(n3150), .I1(VCC_net), 
            .CO(n30757));
    SB_LUT4 rem_4_add_2122_9_lut (.I0(GND_net), .I1(n3151), .I2(VCC_net), 
            .I3(n30755), .O(n3218)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_553_13 (.CI(n30443), .I0(n45865), .I1(n14_adj_4332), 
            .CO(n30444));
    SB_LUT4 rem_4_add_1586_9_lut (.I0(GND_net), .I1(n2352), .I2(VCC_net), 
            .I3(n31214), .O(n2419)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_9 (.CI(n31214), .I0(n2352), .I1(VCC_net), 
            .CO(n31215));
    SB_CARRY rem_4_add_2122_9 (.CI(n30755), .I0(n3151), .I1(VCC_net), 
            .CO(n30756));
    SB_LUT4 rem_4_add_1586_8_lut (.I0(GND_net), .I1(n2353), .I2(VCC_net), 
            .I3(n31213), .O(n2420)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_8 (.CI(n31213), .I0(n2353), .I1(VCC_net), 
            .CO(n31214));
    SB_LUT4 rem_4_add_2122_8_lut (.I0(GND_net), .I1(n3152), .I2(VCC_net), 
            .I3(n30754), .O(n3219)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_8 (.CI(n30754), .I0(n3152), .I1(VCC_net), 
            .CO(n30755));
    SB_LUT4 rem_4_add_1586_7_lut (.I0(GND_net), .I1(n2354), .I2(GND_net), 
            .I3(n31212), .O(n2421)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_7_lut (.I0(GND_net), .I1(n3153), .I2(VCC_net), 
            .I3(n30753), .O(n3220)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_7 (.CI(n30753), .I0(n3153), .I1(VCC_net), 
            .CO(n30754));
    SB_LUT4 rem_4_add_2122_6_lut (.I0(GND_net), .I1(n3154), .I2(GND_net), 
            .I3(n30752), .O(n3221)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_6 (.CI(n30752), .I0(n3154), .I1(GND_net), 
            .CO(n30753));
    SB_LUT4 rem_4_add_2122_5_lut (.I0(GND_net), .I1(n3155), .I2(GND_net), 
            .I3(n30751), .O(n3222)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_mux_3_i17_3_lut (.I0(encoder0_position[16]), .I1(n9_adj_4370), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n375));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1586_7 (.CI(n31212), .I0(n2354), .I1(GND_net), 
            .CO(n31213));
    SB_LUT4 rem_4_add_1586_6_lut (.I0(GND_net), .I1(n2355), .I2(GND_net), 
            .I3(n31211), .O(n2422)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_742_i41_2_lut (.I0(n1172), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4607));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_742_i41_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_2122_5 (.CI(n30751), .I0(n3155), .I1(GND_net), 
            .CO(n30752));
    SB_LUT4 add_553_12_lut (.I0(duty[10]), .I1(n45865), .I2(n15), .I3(n30442), 
            .O(pwm_setpoint_22__N_57[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_2122_4_lut (.I0(GND_net), .I1(n3156), .I2(VCC_net), 
            .I3(n30750), .O(n3223)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_6 (.CI(n31211), .I0(n2355), .I1(GND_net), 
            .CO(n31212));
    SB_CARRY rem_4_add_2122_4 (.CI(n30750), .I0(n3156), .I1(VCC_net), 
            .CO(n30751));
    SB_LUT4 rem_4_i1727_3_lut (.I0(n2542_adj_4520), .I1(n2609), .I2(n2570), 
            .I3(GND_net), .O(n2641));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2122_3_lut (.I0(GND_net), .I1(n3157), .I2(VCC_net), 
            .I3(n30749), .O(n3224)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i744_1_lut (.I0(n1193), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1194));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i744_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_1586_5_lut (.I0(GND_net), .I1(n2356), .I2(VCC_net), 
            .I3(n31210), .O(n2423)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_657_i40_3_lut_3_lut (.I0(n1046), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n40_adj_4599));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_657_i40_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_36_LessThan_742_i36_4_lut (.I0(n375), .I1(n99), .I2(n1175), 
            .I3(n558), .O(n36_adj_4604));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_742_i36_4_lut.LUT_INIT = 16'h0317;
    SB_CARRY rem_4_add_1586_5 (.CI(n31210), .I0(n2356), .I1(VCC_net), 
            .CO(n31211));
    SB_CARRY rem_4_add_2122_3 (.CI(n30749), .I0(n3157), .I1(VCC_net), 
            .CO(n30750));
    SB_LUT4 rem_4_add_1586_4_lut (.I0(GND_net), .I1(n2357_adj_4589), .I2(VCC_net), 
            .I3(n31209), .O(n2424)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_2_lut (.I0(GND_net), .I1(n3158), .I2(GND_net), 
            .I3(VCC_net), .O(n3225)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_2 (.CI(VCC_net), .I0(n3158), .I1(GND_net), 
            .CO(n30749));
    SB_LUT4 rem_4_add_2189_30_lut (.I0(n3263), .I1(n3230), .I2(VCC_net), 
            .I3(n30748), .O(n40712)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_1586_4 (.CI(n31209), .I0(n2357_adj_4589), .I1(VCC_net), 
            .CO(n31210));
    SB_LUT4 i36079_3_lut_4_lut (.I0(n1046), .I1(n97), .I2(n98), .I3(n1047), 
            .O(n43203));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36079_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 rem_4_add_1586_3_lut (.I0(GND_net), .I1(n2358_adj_4588), .I2(GND_net), 
            .I3(n31208), .O(n2425)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_3 (.CI(n31208), .I0(n2358_adj_4588), .I1(GND_net), 
            .CO(n31209));
    SB_LUT4 rem_4_add_2189_29_lut (.I0(GND_net), .I1(n3231), .I2(VCC_net), 
            .I3(n30747), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_29 (.CI(n30747), .I0(n3231), .I1(VCC_net), 
            .CO(n30748));
    SB_CARRY rem_4_add_1586_2 (.CI(VCC_net), .I0(n2458_adj_4575), .I1(VCC_net), 
            .CO(n31208));
    SB_LUT4 div_36_LessThan_742_i40_3_lut (.I0(n38_adj_4605), .I1(n96), 
            .I2(n41_adj_4607), .I3(GND_net), .O(n40_adj_4606));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_742_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_add_2189_28_lut (.I0(GND_net), .I1(n3232), .I2(VCC_net), 
            .I3(n30746), .O(n3299)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_28 (.CI(n30746), .I0(n3232), .I1(VCC_net), 
            .CO(n30747));
    SB_LUT4 i37908_4_lut (.I0(n40_adj_4606), .I1(n36_adj_4604), .I2(n41_adj_4607), 
            .I3(n43178), .O(n45033));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37908_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i37909_3_lut (.I0(n45033), .I1(n95_adj_4360), .I2(n1171), 
            .I3(GND_net), .O(n45034));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37909_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_36_i808_3_lut_3_lut (.I0(n1193), .I1(n6910), .I2(n1175), 
            .I3(GND_net), .O(n1298));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i808_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_2189_27_lut (.I0(GND_net), .I1(n3233), .I2(VCC_net), 
            .I3(n30745), .O(n3300)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_27 (.CI(n30745), .I0(n3233), .I1(VCC_net), 
            .CO(n30746));
    SB_CARRY add_553_12 (.CI(n30442), .I0(n45865), .I1(n15), .CO(n30443));
    SB_LUT4 rem_4_add_2189_26_lut (.I0(GND_net), .I1(n3234), .I2(VCC_net), 
            .I3(n30744), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37840_3_lut (.I0(n45034), .I1(n94), .I2(n1170), .I3(GND_net), 
            .O(n44965));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37840_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1709 (.I0(n44965), .I1(n17287), .I2(n93), .I3(n1169), 
            .O(n1193));
    defparam i1_4_lut_adj_1709.LUT_INIT = 16'hceef;
    SB_LUT4 div_36_i807_3_lut_3_lut (.I0(n1193), .I1(n6909), .I2(n1174), 
            .I3(GND_net), .O(n1297));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i807_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_553_11_lut (.I0(duty[9]), .I1(n45865), .I2(n16_adj_4333), 
            .I3(n30441), .O(pwm_setpoint_22__N_57[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_11_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_36_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4560));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_2189_26 (.CI(n30744), .I0(n3234), .I1(VCC_net), 
            .CO(n30745));
    SB_LUT4 rem_4_add_2189_25_lut (.I0(GND_net), .I1(n3235), .I2(VCC_net), 
            .I3(n30743), .O(n3302)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_25 (.CI(n30743), .I0(n3235), .I1(VCC_net), 
            .CO(n30744));
    SB_LUT4 rem_4_add_2189_24_lut (.I0(GND_net), .I1(n3236), .I2(VCC_net), 
            .I3(n30742), .O(n3303)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_657_i43_2_lut (.I0(n1045), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_657_i43_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_2189_24 (.CI(n30742), .I0(n3236), .I1(VCC_net), 
            .CO(n30743));
    SB_LUT4 rem_4_i1725_3_lut (.I0(n2540_adj_4570), .I1(n2607), .I2(n2570), 
            .I3(GND_net), .O(n2639));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2189_23_lut (.I0(GND_net), .I1(n3237), .I2(VCC_net), 
            .I3(n30741), .O(n3304)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_23 (.CI(n30741), .I0(n3237), .I1(VCC_net), 
            .CO(n30742));
    SB_LUT4 div_36_mux_3_i18_3_lut (.I0(encoder0_position[17]), .I1(n8_adj_4369), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n374));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2189_22_lut (.I0(GND_net), .I1(n3238), .I2(VCC_net), 
            .I3(n30740), .O(n3305)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_553_11 (.CI(n30441), .I0(n45865), .I1(n16_adj_4333), 
            .CO(n30442));
    SB_CARRY rem_4_add_2189_22 (.CI(n30740), .I0(n3238), .I1(VCC_net), 
            .CO(n30741));
    SB_LUT4 rem_4_add_2189_21_lut (.I0(GND_net), .I1(n3239), .I2(VCC_net), 
            .I3(n30739), .O(n3306)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_553_10_lut (.I0(duty[8]), .I1(n45865), .I2(n17), .I3(n30440), 
            .O(pwm_setpoint_22__N_57[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_36_i809_3_lut_3_lut (.I0(n1193), .I1(n6911), .I2(n375), 
            .I3(GND_net), .O(n1299));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i809_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_2189_21 (.CI(n30739), .I0(n3239), .I1(VCC_net), 
            .CO(n30740));
    SB_LUT4 div_36_i659_1_lut (.I0(n1067), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1068));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i659_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_2189_20_lut (.I0(GND_net), .I1(n3240), .I2(VCC_net), 
            .I3(n30738), .O(n3307)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_20 (.CI(n30738), .I0(n3240), .I1(VCC_net), 
            .CO(n30739));
    SB_LUT4 rem_4_add_2189_19_lut (.I0(GND_net), .I1(n3241), .I2(VCC_net), 
            .I3(n30737), .O(n3308)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_553_10 (.CI(n30440), .I0(n45865), .I1(n17), .CO(n30441));
    SB_CARRY rem_4_add_2189_19 (.CI(n30737), .I0(n3241), .I1(VCC_net), 
            .CO(n30738));
    SB_LUT4 add_553_9_lut (.I0(duty[7]), .I1(n45865), .I2(n18_adj_4334), 
            .I3(n30439), .O(pwm_setpoint_22__N_57[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_2189_18_lut (.I0(GND_net), .I1(n3242), .I2(VCC_net), 
            .I3(n30736), .O(n3309)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_553_9 (.CI(n30439), .I0(n45865), .I1(n18_adj_4334), .CO(n30440));
    SB_CARRY rem_4_add_2189_18 (.CI(n30736), .I0(n3242), .I1(VCC_net), 
            .CO(n30737));
    SB_LUT4 rem_4_add_2189_17_lut (.I0(GND_net), .I1(n3243), .I2(VCC_net), 
            .I3(n30735), .O(n3310)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_17 (.CI(n30735), .I0(n3243), .I1(VCC_net), 
            .CO(n30736));
    SB_LUT4 add_553_8_lut (.I0(duty[6]), .I1(n45865), .I2(n19), .I3(n30438), 
            .O(pwm_setpoint_22__N_57[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_2189_16_lut (.I0(GND_net), .I1(n3244), .I2(VCC_net), 
            .I3(n30734), .O(n3311)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_16 (.CI(n30734), .I0(n3244), .I1(VCC_net), 
            .CO(n30735));
    SB_LUT4 div_36_LessThan_657_i38_4_lut (.I0(n374), .I1(n99), .I2(n1048), 
            .I3(n558), .O(n38_adj_4598));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_657_i38_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 rem_4_add_2189_15_lut (.I0(GND_net), .I1(n3245), .I2(VCC_net), 
            .I3(n30733), .O(n3312)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_LessThan_657_i42_3_lut (.I0(n40_adj_4599), .I1(n96), 
            .I2(n43), .I3(GND_net), .O(n42_adj_4600));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_657_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_2189_15 (.CI(n30733), .I0(n3245), .I1(VCC_net), 
            .CO(n30734));
    SB_LUT4 rem_4_add_2189_14_lut (.I0(GND_net), .I1(n3246), .I2(VCC_net), 
            .I3(n30732), .O(n3313)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_14 (.CI(n30732), .I0(n3246), .I1(VCC_net), 
            .CO(n30733));
    SB_LUT4 rem_4_add_2189_13_lut (.I0(GND_net), .I1(n3247), .I2(VCC_net), 
            .I3(n30731), .O(n3314)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_13 (.CI(n30731), .I0(n3247), .I1(VCC_net), 
            .CO(n30732));
    SB_LUT4 rem_4_add_2189_12_lut (.I0(GND_net), .I1(n3248), .I2(VCC_net), 
            .I3(n30730), .O(n3315)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37508_4_lut (.I0(n42_adj_4600), .I1(n38_adj_4598), .I2(n43), 
            .I3(n43203), .O(n44633));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37508_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY rem_4_add_2189_12 (.CI(n30730), .I0(n3248), .I1(VCC_net), 
            .CO(n30731));
    SB_LUT4 rem_4_add_2189_11_lut (.I0(GND_net), .I1(n3249), .I2(VCC_net), 
            .I3(n30729), .O(n3316)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37509_3_lut (.I0(n44633), .I1(n95_adj_4360), .I2(n1044), 
            .I3(GND_net), .O(n44634));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37509_3_lut.LUT_INIT = 16'h2b2b;
    SB_CARRY rem_4_add_2189_11 (.CI(n30729), .I0(n3249), .I1(VCC_net), 
            .CO(n30730));
    SB_LUT4 i1_4_lut_adj_1710 (.I0(n44634), .I1(n17284), .I2(n94), .I3(n1043), 
            .O(n1067));
    defparam i1_4_lut_adj_1710.LUT_INIT = 16'hceef;
    SB_LUT4 rem_4_add_2189_10_lut (.I0(GND_net), .I1(n3250), .I2(VCC_net), 
            .I3(n30728), .O(n3317)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_10 (.CI(n30728), .I0(n3250), .I1(VCC_net), 
            .CO(n30729));
    SB_CARRY add_553_8 (.CI(n30438), .I0(n45865), .I1(n19), .CO(n30439));
    SB_LUT4 rem_4_add_2189_9_lut (.I0(GND_net), .I1(n3251), .I2(VCC_net), 
            .I3(n30727), .O(n3318)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_9 (.CI(n30727), .I0(n3251), .I1(VCC_net), 
            .CO(n30728));
    SB_LUT4 rem_4_add_2189_8_lut (.I0(GND_net), .I1(n3252), .I2(VCC_net), 
            .I3(n30726), .O(n3319)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_8 (.CI(n30726), .I0(n3252), .I1(VCC_net), 
            .CO(n30727));
    SB_LUT4 rem_4_add_2189_7_lut (.I0(GND_net), .I1(n3253), .I2(VCC_net), 
            .I3(n30725), .O(n3320)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_7 (.CI(n30725), .I0(n3253), .I1(VCC_net), 
            .CO(n30726));
    SB_LUT4 rem_4_add_2189_6_lut (.I0(GND_net), .I1(n3254), .I2(GND_net), 
            .I3(n30724), .O(n3321)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_6 (.CI(n30724), .I0(n3254), .I1(GND_net), 
            .CO(n30725));
    SB_LUT4 rem_4_add_2189_5_lut (.I0(GND_net), .I1(n3255), .I2(GND_net), 
            .I3(n30723), .O(n3322)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_5 (.CI(n30723), .I0(n3255), .I1(GND_net), 
            .CO(n30724));
    SB_LUT4 rem_4_add_2189_4_lut (.I0(GND_net), .I1(n3256), .I2(VCC_net), 
            .I3(n30722), .O(n3323)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i805_3_lut_3_lut (.I0(n1193), .I1(n6907), .I2(n1172), 
            .I3(GND_net), .O(n1295));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i805_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_2189_4 (.CI(n30722), .I0(n3256), .I1(VCC_net), 
            .CO(n30723));
    SB_LUT4 rem_4_add_2189_3_lut (.I0(GND_net), .I1(n3257), .I2(VCC_net), 
            .I3(n30721), .O(n3324)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_3 (.CI(n30721), .I0(n3257), .I1(VCC_net), 
            .CO(n30722));
    SB_LUT4 rem_4_add_2189_2_lut (.I0(GND_net), .I1(n3258), .I2(GND_net), 
            .I3(VCC_net), .O(n3325)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_2 (.CI(VCC_net), .I0(n3258), .I1(GND_net), 
            .CO(n30721));
    SB_LUT4 add_3158_16_lut (.I0(GND_net), .I1(n1967), .I2(n86), .I3(n30720), 
            .O(n6996)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3158_15_lut (.I0(GND_net), .I1(n1968), .I2(n87), .I3(n30719), 
            .O(n6997)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3158_15 (.CI(n30719), .I0(n1968), .I1(n87), .CO(n30720));
    SB_LUT4 add_3158_14_lut (.I0(GND_net), .I1(n1969), .I2(n88), .I3(n30718), 
            .O(n6998)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_553_7_lut (.I0(duty[5]), .I1(n45865), .I2(n20), .I3(n30437), 
            .O(pwm_setpoint_22__N_57[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3158_14 (.CI(n30718), .I0(n1969), .I1(n88), .CO(n30719));
    SB_LUT4 add_3158_13_lut (.I0(GND_net), .I1(n1970), .I2(n89), .I3(n30717), 
            .O(n6999)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3158_13 (.CI(n30717), .I0(n1970), .I1(n89), .CO(n30718));
    SB_LUT4 add_3158_12_lut (.I0(GND_net), .I1(n1971), .I2(n90), .I3(n30716), 
            .O(n7000)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3158_12 (.CI(n30716), .I0(n1971), .I1(n90), .CO(n30717));
    SB_LUT4 add_3158_11_lut (.I0(GND_net), .I1(n1972), .I2(n91), .I3(n30715), 
            .O(n7001)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3158_11 (.CI(n30715), .I0(n1972), .I1(n91), .CO(n30716));
    SB_LUT4 add_3158_10_lut (.I0(GND_net), .I1(n1973), .I2(n92), .I3(n30714), 
            .O(n7002)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3158_10 (.CI(n30714), .I0(n1973), .I1(n92), .CO(n30715));
    SB_LUT4 add_3158_9_lut (.I0(GND_net), .I1(n1974), .I2(n93), .I3(n30713), 
            .O(n7003)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3158_9 (.CI(n30713), .I0(n1974), .I1(n93), .CO(n30714));
    SB_LUT4 add_3158_8_lut (.I0(GND_net), .I1(n1975), .I2(n94), .I3(n30712), 
            .O(n7004)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3158_8 (.CI(n30712), .I0(n1975), .I1(n94), .CO(n30713));
    SB_LUT4 add_3158_7_lut (.I0(GND_net), .I1(n1976), .I2(n95_adj_4360), 
            .I3(n30711), .O(n7005)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_553_7 (.CI(n30437), .I0(n45865), .I1(n20), .CO(n30438));
    SB_CARRY add_3158_7 (.CI(n30711), .I0(n1976), .I1(n95_adj_4360), .CO(n30712));
    SB_LUT4 add_553_6_lut (.I0(duty[4]), .I1(n45865), .I2(n21_adj_4335), 
            .I3(n30436), .O(pwm_setpoint_22__N_57[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_3158_6_lut (.I0(GND_net), .I1(n1977), .I2(n96), .I3(n30710), 
            .O(n7006)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3158_6 (.CI(n30710), .I0(n1977), .I1(n96), .CO(n30711));
    SB_LUT4 add_3158_5_lut (.I0(GND_net), .I1(n1978), .I2(n97), .I3(n30709), 
            .O(n7007)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i804_3_lut_3_lut (.I0(n1193), .I1(n6906), .I2(n1171), 
            .I3(GND_net), .O(n1294));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i804_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_553_6 (.CI(n30436), .I0(n45865), .I1(n21_adj_4335), .CO(n30437));
    SB_LUT4 div_36_i806_3_lut_3_lut (.I0(n1193), .I1(n6908), .I2(n1173), 
            .I3(GND_net), .O(n1296));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i806_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i802_3_lut_3_lut (.I0(n1193), .I1(n6904), .I2(n1169), 
            .I3(GND_net), .O(n1292));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i802_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3158_5 (.CI(n30709), .I0(n1978), .I1(n97), .CO(n30710));
    SB_LUT4 add_3158_4_lut (.I0(GND_net), .I1(n1979), .I2(n98), .I3(n30708), 
            .O(n7008)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3158_4 (.CI(n30708), .I0(n1979), .I1(n98), .CO(n30709));
    SB_LUT4 add_3158_3_lut (.I0(GND_net), .I1(n1980), .I2(n99), .I3(n30707), 
            .O(n7009)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3158_3 (.CI(n30707), .I0(n1980), .I1(n99), .CO(n30708));
    SB_LUT4 add_3158_2_lut (.I0(GND_net), .I1(n382), .I2(n558), .I3(VCC_net), 
            .O(n7010)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3158_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_553_5_lut (.I0(duty[3]), .I1(n45865), .I2(n22_adj_4336), 
            .I3(n30435), .O(pwm_setpoint_22__N_57[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3158_2 (.CI(VCC_net), .I0(n382), .I1(n558), .CO(n30707));
    SB_LUT4 div_36_i803_3_lut_3_lut (.I0(n1193), .I1(n6905), .I2(n1170), 
            .I3(GND_net), .O(n1293));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i803_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_LessThan_742_i38_3_lut_3_lut (.I0(n1173), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n38_adj_4605));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_742_i38_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 add_3157_15_lut (.I0(GND_net), .I1(n1862), .I2(n87), .I3(n30706), 
            .O(n6980)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3157_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3157_14_lut (.I0(GND_net), .I1(n1863), .I2(n88), .I3(n30705), 
            .O(n6981)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3157_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3157_14 (.CI(n30705), .I0(n1863), .I1(n88), .CO(n30706));
    SB_LUT4 add_3157_13_lut (.I0(GND_net), .I1(n1864), .I2(n89), .I3(n30704), 
            .O(n6982)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3157_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3157_13 (.CI(n30704), .I0(n1864), .I1(n89), .CO(n30705));
    SB_LUT4 add_3157_12_lut (.I0(GND_net), .I1(n1865), .I2(n90), .I3(n30703), 
            .O(n6983)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3157_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36054_3_lut_4_lut (.I0(n1173), .I1(n97), .I2(n98), .I3(n1174), 
            .O(n43178));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36054_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_CARRY add_553_5 (.CI(n30435), .I0(n45865), .I1(n22_adj_4336), .CO(n30436));
    SB_LUT4 div_36_i890_3_lut_3_lut (.I0(n1316), .I1(n6921), .I2(n1299), 
            .I3(GND_net), .O(n1419));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i890_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i891_3_lut_3_lut (.I0(n1316), .I1(n6922), .I2(n376), 
            .I3(GND_net), .O(n1420));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i891_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3157_12 (.CI(n30703), .I0(n1865), .I1(n90), .CO(n30704));
    SB_LUT4 add_3157_11_lut (.I0(GND_net), .I1(n1866), .I2(n91), .I3(n30702), 
            .O(n6984)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3157_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3157_11 (.CI(n30702), .I0(n1866), .I1(n91), .CO(n30703));
    SB_LUT4 rem_4_i1726_3_lut (.I0(n2541_adj_4569), .I1(n2608), .I2(n2570), 
            .I3(GND_net), .O(n2640));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3157_10_lut (.I0(GND_net), .I1(n1867), .I2(n92), .I3(n30701), 
            .O(n6985)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3157_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3157_10 (.CI(n30701), .I0(n1867), .I1(n92), .CO(n30702));
    SB_LUT4 add_3157_9_lut (.I0(GND_net), .I1(n1868), .I2(n93), .I3(n30700), 
            .O(n6986)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3157_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3157_9 (.CI(n30700), .I0(n1868), .I1(n93), .CO(n30701));
    SB_LUT4 div_36_i887_3_lut_3_lut (.I0(n1316), .I1(n6918), .I2(n1296), 
            .I3(GND_net), .O(n1416));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i887_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3157_8_lut (.I0(GND_net), .I1(n1869), .I2(n94), .I3(n30699), 
            .O(n6987)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3157_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3157_8 (.CI(n30699), .I0(n1869), .I1(n94), .CO(n30700));
    SB_LUT4 add_3157_7_lut (.I0(GND_net), .I1(n1870), .I2(n95_adj_4360), 
            .I3(n30698), .O(n6988)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3157_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3157_7 (.CI(n30698), .I0(n1870), .I1(n95_adj_4360), .CO(n30699));
    SB_LUT4 add_3157_6_lut (.I0(GND_net), .I1(n1871), .I2(n96), .I3(n30697), 
            .O(n6989)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3157_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_553_4_lut (.I0(duty[2]), .I1(n45865), .I2(n23_adj_4337), 
            .I3(n30434), .O(pwm_setpoint_22__N_57[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_3157_6 (.CI(n30697), .I0(n1871), .I1(n96), .CO(n30698));
    SB_LUT4 add_3157_5_lut (.I0(GND_net), .I1(n1872), .I2(n97), .I3(n30696), 
            .O(n6990)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3157_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3157_5 (.CI(n30696), .I0(n1872), .I1(n97), .CO(n30697));
    SB_LUT4 add_3157_4_lut (.I0(GND_net), .I1(n1873), .I2(n98), .I3(n30695), 
            .O(n6991)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3157_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1724_3_lut (.I0(n2539_adj_4571), .I1(n2606), .I2(n2570), 
            .I3(GND_net), .O(n2638_adj_4491));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i888_3_lut_3_lut (.I0(n1316), .I1(n6919), .I2(n1297), 
            .I3(GND_net), .O(n1417));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i888_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3157_4 (.CI(n30695), .I0(n1873), .I1(n98), .CO(n30696));
    SB_LUT4 add_3157_3_lut (.I0(GND_net), .I1(n1874), .I2(n99), .I3(n30694), 
            .O(n6992)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3157_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i886_3_lut_3_lut (.I0(n1316), .I1(n6917), .I2(n1295), 
            .I3(GND_net), .O(n1415));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i886_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_648_8_lut (.I0(n986), .I1(n953), .I2(VCC_net), .I3(n31448), 
            .O(n1052)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3157_3 (.CI(n30694), .I0(n1874), .I1(n99), .CO(n30695));
    SB_LUT4 rem_4_add_648_7_lut (.I0(GND_net), .I1(n954), .I2(GND_net), 
            .I3(n31447), .O(n1021)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_7 (.CI(n31447), .I0(n954), .I1(GND_net), .CO(n31448));
    SB_LUT4 add_3157_2_lut (.I0(GND_net), .I1(n381), .I2(n558), .I3(VCC_net), 
            .O(n6993)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3157_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3157_2 (.CI(VCC_net), .I0(n381), .I1(n558), .CO(n30694));
    SB_LUT4 add_3156_14_lut (.I0(GND_net), .I1(n1754), .I2(n88), .I3(n30693), 
            .O(n6965)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3156_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_648_6_lut (.I0(GND_net), .I1(n955), .I2(GND_net), 
            .I3(n31446), .O(n1022)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3156_13_lut (.I0(GND_net), .I1(n1755), .I2(n89), .I3(n30692), 
            .O(n6966)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3156_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3156_13 (.CI(n30692), .I0(n1755), .I1(n89), .CO(n30693));
    SB_LUT4 add_3156_12_lut (.I0(GND_net), .I1(n1756), .I2(n90), .I3(n30691), 
            .O(n6967)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3156_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_6 (.CI(n31446), .I0(n955), .I1(GND_net), .CO(n31447));
    SB_LUT4 div_36_i885_3_lut_3_lut (.I0(n1316), .I1(n6916), .I2(n1294), 
            .I3(GND_net), .O(n1414));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i885_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_648_5_lut (.I0(GND_net), .I1(n956), .I2(VCC_net), 
            .I3(n31445), .O(n1023)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1711 (.I0(n5_adj_4440), .I1(n63_adj_4439), .I2(n2664), 
            .I3(n20639), .O(n6_adj_4626));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1711.LUT_INIT = 16'heaaa;
    SB_CARRY rem_4_add_648_5 (.CI(n31445), .I0(n956), .I1(VCC_net), .CO(n31446));
    SB_CARRY add_3156_12 (.CI(n30691), .I0(n1756), .I1(n90), .CO(n30692));
    SB_LUT4 add_3156_11_lut (.I0(GND_net), .I1(n1757), .I2(n91), .I3(n30690), 
            .O(n6968)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3156_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3156_11 (.CI(n30690), .I0(n1757), .I1(n91), .CO(n30691));
    SB_LUT4 add_3156_10_lut (.I0(GND_net), .I1(n1758), .I2(n92), .I3(n30689), 
            .O(n6969)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3156_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3156_10 (.CI(n30689), .I0(n1758), .I1(n92), .CO(n30690));
    SB_LUT4 div_36_i883_3_lut_3_lut (.I0(n1316), .I1(n6914), .I2(n1292), 
            .I3(GND_net), .O(n1412));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i883_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_648_4_lut (.I0(GND_net), .I1(n957), .I2(VCC_net), 
            .I3(n31444), .O(n1024)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3156_9_lut (.I0(GND_net), .I1(n1759), .I2(n93), .I3(n30688), 
            .O(n6970)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3156_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_4 (.CI(n31444), .I0(n957), .I1(VCC_net), .CO(n31445));
    SB_LUT4 rem_4_add_648_3_lut (.I0(GND_net), .I1(n958), .I2(GND_net), 
            .I3(n31443), .O(n1025)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_3 (.CI(n31443), .I0(n958), .I1(GND_net), .CO(n31444));
    SB_CARRY add_3156_9 (.CI(n30688), .I0(n1759), .I1(n93), .CO(n30689));
    SB_CARRY rem_4_add_648_2 (.CI(VCC_net), .I0(n1058), .I1(VCC_net), 
            .CO(n31443));
    SB_LUT4 add_3156_8_lut (.I0(GND_net), .I1(n1760), .I2(n94), .I3(n30687), 
            .O(n6971)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3156_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3156_8 (.CI(n30687), .I0(n1760), .I1(n94), .CO(n30688));
    SB_LUT4 add_3156_7_lut (.I0(GND_net), .I1(n1761), .I2(n95_adj_4360), 
            .I3(n30686), .O(n6972)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3156_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3156_7 (.CI(n30686), .I0(n1761), .I1(n95_adj_4360), .CO(n30687));
    SB_LUT4 add_3156_6_lut (.I0(GND_net), .I1(n1762), .I2(n96), .I3(n30685), 
            .O(n6973)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3156_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11_4_lut_adj_1712 (.I0(n2638_adj_4491), .I1(n2640), .I2(n2639), 
            .I3(n2641), .O(n30));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i11_4_lut_adj_1712.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_715_9_lut (.I0(n1085), .I1(n1052), .I2(VCC_net), 
            .I3(n31442), .O(n1151)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3156_6 (.CI(n30685), .I0(n1762), .I1(n96), .CO(n30686));
    SB_LUT4 rem_4_add_715_8_lut (.I0(GND_net), .I1(n1053), .I2(VCC_net), 
            .I3(n31441), .O(n1120)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3156_5_lut (.I0(GND_net), .I1(n1763), .I2(n97), .I3(n30684), 
            .O(n6974)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3156_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_553_4 (.CI(n30434), .I0(n45865), .I1(n23_adj_4337), .CO(n30435));
    SB_CARRY add_3156_5 (.CI(n30684), .I0(n1763), .I1(n97), .CO(n30685));
    SB_LUT4 add_553_3_lut (.I0(duty[1]), .I1(n45865), .I2(n24_adj_4338), 
            .I3(n30433), .O(pwm_setpoint_22__N_57[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_715_8 (.CI(n31441), .I0(n1053), .I1(VCC_net), .CO(n31442));
    SB_LUT4 div_36_i884_3_lut_3_lut (.I0(n1316), .I1(n6915), .I2(n1293), 
            .I3(GND_net), .O(n1413));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i884_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i889_3_lut_3_lut (.I0(n1316), .I1(n6920), .I2(n1298), 
            .I3(GND_net), .O(n1418));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i889_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3156_4_lut (.I0(GND_net), .I1(n1764), .I2(n98), .I3(n30683), 
            .O(n6975)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3156_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_715_7_lut (.I0(GND_net), .I1(n1054), .I2(GND_net), 
            .I3(n31440), .O(n1121)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3156_4 (.CI(n30683), .I0(n1764), .I1(n98), .CO(n30684));
    SB_CARRY rem_4_add_715_7 (.CI(n31440), .I0(n1054), .I1(GND_net), .CO(n31441));
    SB_LUT4 i36040_3_lut_4_lut (.I0(n1297), .I1(n97), .I2(n98), .I3(n1298), 
            .O(n43164));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36040_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_36_LessThan_825_i36_3_lut_3_lut (.I0(n1297), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n36_adj_4611));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_825_i36_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 add_3156_3_lut (.I0(GND_net), .I1(n1765), .I2(n99), .I3(n30682), 
            .O(n6976)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3156_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i970_3_lut_3_lut (.I0(n1436), .I1(n6933), .I2(n1420), 
            .I3(GND_net), .O(n1537));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i970_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3156_3 (.CI(n30682), .I0(n1765), .I1(n99), .CO(n30683));
    SB_LUT4 add_3156_2_lut (.I0(GND_net), .I1(n380), .I2(n558), .I3(VCC_net), 
            .O(n6977)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3156_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3156_2 (.CI(VCC_net), .I0(n380), .I1(n558), .CO(n30682));
    SB_LUT4 rem_4_add_715_6_lut (.I0(GND_net), .I1(n1055), .I2(GND_net), 
            .I3(n31439), .O(n1122)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_6 (.CI(n31439), .I0(n1055), .I1(GND_net), .CO(n31440));
    SB_LUT4 add_3155_13_lut (.I0(GND_net), .I1(n1643), .I2(n89), .I3(n30681), 
            .O(n6951)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3155_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i964_3_lut_3_lut (.I0(n1436), .I1(n6927), .I2(n1414), 
            .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i964_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3155_12_lut (.I0(GND_net), .I1(n1644), .I2(n90), .I3(n30680), 
            .O(n6952)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3155_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3155_12 (.CI(n30680), .I0(n1644), .I1(n90), .CO(n30681));
    SB_LUT4 add_3155_11_lut (.I0(GND_net), .I1(n1645), .I2(n91), .I3(n30679), 
            .O(n6953)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3155_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_715_5_lut (.I0(GND_net), .I1(n1056), .I2(VCC_net), 
            .I3(n31438), .O(n1123)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3155_11 (.CI(n30679), .I0(n1645), .I1(n91), .CO(n30680));
    SB_LUT4 div_36_i969_3_lut_3_lut (.I0(n1436), .I1(n6932), .I2(n1419), 
            .I3(GND_net), .O(n1536));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i969_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3155_10_lut (.I0(GND_net), .I1(n1646), .I2(n92), .I3(n30678), 
            .O(n6954)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3155_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3155_10 (.CI(n30678), .I0(n1646), .I1(n92), .CO(n30679));
    SB_LUT4 div_36_i968_3_lut_3_lut (.I0(n1436), .I1(n6931), .I2(n1418), 
            .I3(GND_net), .O(n1535));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i968_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3155_9_lut (.I0(GND_net), .I1(n1647), .I2(n93), .I3(n30677), 
            .O(n6955)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3155_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3155_9 (.CI(n30677), .I0(n1647), .I1(n93), .CO(n30678));
    SB_CARRY rem_4_add_715_5 (.CI(n31438), .I0(n1056), .I1(VCC_net), .CO(n31439));
    SB_LUT4 add_3155_8_lut (.I0(GND_net), .I1(n1648), .I2(n94), .I3(n30676), 
            .O(n6956)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3155_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i967_3_lut_3_lut (.I0(n1436), .I1(n6930), .I2(n1417), 
            .I3(GND_net), .O(n1534));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i967_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3155_8 (.CI(n30676), .I0(n1648), .I1(n94), .CO(n30677));
    SB_CARRY add_553_3 (.CI(n30433), .I0(n45865), .I1(n24_adj_4338), .CO(n30434));
    SB_LUT4 add_3155_7_lut (.I0(GND_net), .I1(n1649), .I2(n95_adj_4360), 
            .I3(n30675), .O(n6957)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3155_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3155_7 (.CI(n30675), .I0(n1649), .I1(n95_adj_4360), .CO(n30676));
    SB_LUT4 rem_4_add_715_4_lut (.I0(GND_net), .I1(n1057), .I2(VCC_net), 
            .I3(n31437), .O(n1124)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_4 (.CI(n31437), .I0(n1057), .I1(VCC_net), .CO(n31438));
    SB_LUT4 rem_4_add_715_3_lut (.I0(GND_net), .I1(n1058), .I2(GND_net), 
            .I3(n31436), .O(n1125)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3155_6_lut (.I0(GND_net), .I1(n1650), .I2(n96), .I3(n30674), 
            .O(n6958)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3155_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_3 (.CI(n31436), .I0(n1058), .I1(GND_net), .CO(n31437));
    SB_CARRY add_3155_6 (.CI(n30674), .I0(n1650), .I1(n96), .CO(n30675));
    SB_LUT4 add_3155_5_lut (.I0(GND_net), .I1(n1651), .I2(n97), .I3(n30673), 
            .O(n6959)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3155_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3155_5 (.CI(n30673), .I0(n1651), .I1(n97), .CO(n30674));
    SB_LUT4 add_3155_4_lut (.I0(GND_net), .I1(n1652), .I2(n98), .I3(n30672), 
            .O(n6960)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3155_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3155_4 (.CI(n30672), .I0(n1652), .I1(n98), .CO(n30673));
    SB_CARRY rem_4_add_715_2 (.CI(VCC_net), .I0(n1158), .I1(VCC_net), 
            .CO(n31436));
    SB_LUT4 rem_4_add_782_10_lut (.I0(n1184), .I1(n1151), .I2(VCC_net), 
            .I3(n31435), .O(n1250)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_782_9_lut (.I0(GND_net), .I1(n1152), .I2(VCC_net), 
            .I3(n31434), .O(n1219)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3155_3_lut (.I0(GND_net), .I1(n1653), .I2(n99), .I3(n30671), 
            .O(n6961)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3155_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_9 (.CI(n31434), .I0(n1152), .I1(VCC_net), .CO(n31435));
    SB_LUT4 rem_4_add_782_8_lut (.I0(GND_net), .I1(n1153), .I2(VCC_net), 
            .I3(n31433), .O(n1220)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i963_3_lut_3_lut (.I0(n1436), .I1(n6926), .I2(n1413), 
            .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i963_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3155_3 (.CI(n30671), .I0(n1653), .I1(n99), .CO(n30672));
    SB_LUT4 add_3155_2_lut (.I0(GND_net), .I1(n379), .I2(n558), .I3(VCC_net), 
            .O(n6962)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3155_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3155_2 (.CI(VCC_net), .I0(n379), .I1(n558), .CO(n30671));
    SB_LUT4 rem_4_add_2298_9_lut (.I0(n45142), .I1(n2_adj_4938), .I2(n3452), 
            .I3(n30670), .O(color_23__N_164[7])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_2298_8_lut (.I0(n45146), .I1(n2_adj_4938), .I2(n3453), 
            .I3(n30669), .O(color_23__N_164[6])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_8 (.CI(n30669), .I0(n2_adj_4938), .I1(n3453), 
            .CO(n30670));
    SB_CARRY rem_4_add_782_8 (.CI(n31433), .I0(n1153), .I1(VCC_net), .CO(n31434));
    SB_LUT4 rem_4_add_2298_7_lut (.I0(n45149), .I1(n2_adj_4938), .I2(n3454), 
            .I3(n30668), .O(color_23__N_164[5])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_36_i971_3_lut_3_lut (.I0(n1436), .I1(n6934), .I2(n377), 
            .I3(GND_net), .O(n1538));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i971_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_782_7_lut (.I0(GND_net), .I1(n1154), .I2(GND_net), 
            .I3(n31432), .O(n1221)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i966_3_lut_3_lut (.I0(n1436), .I1(n6929), .I2(n1416), 
            .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i966_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i965_3_lut_3_lut (.I0(n1436), .I1(n6928), .I2(n1415), 
            .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i965_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_553_2_lut (.I0(duty[0]), .I1(n45865), .I2(n25), .I3(VCC_net), 
            .O(pwm_setpoint_22__N_57[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_553_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_7 (.CI(n30668), .I0(n2_adj_4938), .I1(n3454), 
            .CO(n30669));
    SB_CARRY rem_4_add_782_7 (.CI(n31432), .I0(n1154), .I1(GND_net), .CO(n31433));
    SB_LUT4 rem_4_add_782_6_lut (.I0(GND_net), .I1(n1155), .I2(GND_net), 
            .I3(n31431), .O(n1222)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_6 (.CI(n31431), .I0(n1155), .I1(GND_net), .CO(n31432));
    SB_LUT4 rem_4_add_2298_6_lut (.I0(n45152), .I1(n2_adj_4938), .I2(n3455), 
            .I3(n30667), .O(color_23__N_164[4])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_6 (.CI(n30667), .I0(n2_adj_4938), .I1(n3455), 
            .CO(n30668));
    SB_LUT4 rem_4_add_2298_5_lut (.I0(n45155), .I1(n2_adj_4938), .I2(n3456), 
            .I3(n30666), .O(color_23__N_164[3])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_5 (.CI(n30666), .I0(n2_adj_4938), .I1(n3456), 
            .CO(n30667));
    SB_LUT4 div_36_i962_3_lut_3_lut (.I0(n1436), .I1(n6925), .I2(n1412), 
            .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i962_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_2298_4_lut (.I0(n45158), .I1(n2_adj_4938), .I2(n3457), 
            .I3(n30665), .O(color_23__N_164[2])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_782_5_lut (.I0(GND_net), .I1(n1156), .I2(VCC_net), 
            .I3(n31430), .O(n1223)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2298_4 (.CI(n30665), .I0(n2_adj_4938), .I1(n3457), 
            .CO(n30666));
    SB_CARRY rem_4_add_782_5 (.CI(n31430), .I0(n1156), .I1(VCC_net), .CO(n31431));
    SB_LUT4 rem_4_add_2298_3_lut (.I0(communication_counter[1]), .I1(n2_adj_4938), 
            .I2(n3458), .I3(n30664), .O(color_23__N_164[1])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_3 (.CI(n30664), .I0(n2_adj_4938), .I1(n3458), 
            .CO(n30665));
    SB_LUT4 rem_4_add_782_4_lut (.I0(GND_net), .I1(n1157), .I2(VCC_net), 
            .I3(n31429), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_4 (.CI(n31429), .I0(n1157), .I1(VCC_net), .CO(n31430));
    SB_LUT4 rem_4_add_782_3_lut (.I0(GND_net), .I1(n1158), .I2(GND_net), 
            .I3(n31428), .O(n1225)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_3 (.CI(n31428), .I0(n1158), .I1(GND_net), .CO(n31429));
    SB_LUT4 rem_4_add_2298_2_lut (.I0(communication_counter[0]), .I1(n2_adj_4938), 
            .I2(n3459), .I3(VCC_net), .O(color_23__N_164[0])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_2 (.CI(VCC_net), .I0(n2_adj_4938), .I1(n3459), 
            .CO(n30664));
    SB_LUT4 add_3154_12_lut (.I0(GND_net), .I1(n1529), .I2(n90), .I3(n30663), 
            .O(n6938)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3154_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3154_11_lut (.I0(GND_net), .I1(n1530), .I2(n91), .I3(n30662), 
            .O(n6939)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3154_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3154_11 (.CI(n30662), .I0(n1530), .I1(n91), .CO(n30663));
    SB_CARRY add_553_2 (.CI(VCC_net), .I0(n45865), .I1(n25), .CO(n30433));
    SB_CARRY rem_4_add_782_2 (.CI(VCC_net), .I0(n1258), .I1(VCC_net), 
            .CO(n31428));
    SB_LUT4 add_3154_10_lut (.I0(GND_net), .I1(n1531), .I2(n92), .I3(n30661), 
            .O(n6940)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3154_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_849_11_lut (.I0(n1283), .I1(n1250), .I2(VCC_net), 
            .I3(n31427), .O(n1349)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_849_10_lut (.I0(GND_net), .I1(n1251), .I2(VCC_net), 
            .I3(n31426), .O(n1318)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3154_10 (.CI(n30661), .I0(n1531), .I1(n92), .CO(n30662));
    SB_LUT4 add_3154_9_lut (.I0(GND_net), .I1(n1532), .I2(n93), .I3(n30660), 
            .O(n6941)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3154_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_10 (.CI(n31426), .I0(n1251), .I1(VCC_net), 
            .CO(n31427));
    SB_CARRY add_3154_9 (.CI(n30660), .I0(n1532), .I1(n93), .CO(n30661));
    SB_LUT4 add_3154_8_lut (.I0(GND_net), .I1(n1533), .I2(n94), .I3(n30659), 
            .O(n6942)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3154_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3154_8 (.CI(n30659), .I0(n1533), .I1(n94), .CO(n30660));
    SB_LUT4 add_3154_7_lut (.I0(GND_net), .I1(n1534), .I2(n95_adj_4360), 
            .I3(n30658), .O(n6943)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3154_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3154_7 (.CI(n30658), .I0(n1534), .I1(n95_adj_4360), .CO(n30659));
    SB_LUT4 rem_4_add_849_9_lut (.I0(GND_net), .I1(n1252), .I2(VCC_net), 
            .I3(n31425), .O(n1319)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3154_6_lut (.I0(GND_net), .I1(n1535), .I2(n96), .I3(n30657), 
            .O(n6944)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3154_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3154_6 (.CI(n30657), .I0(n1535), .I1(n96), .CO(n30658));
    SB_LUT4 add_3154_5_lut (.I0(GND_net), .I1(n1536), .I2(n97), .I3(n30656), 
            .O(n6945)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3154_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36004_3_lut_4_lut (.I0(n1418), .I1(n97), .I2(n98), .I3(n1419), 
            .O(n43128));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36004_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_36_LessThan_906_i34_3_lut_3_lut (.I0(n1418), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n34_adj_4621));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_906_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_CARRY add_3154_5 (.CI(n30656), .I0(n1536), .I1(n97), .CO(n30657));
    SB_LUT4 add_3154_4_lut (.I0(GND_net), .I1(n1537), .I2(n98), .I3(n30655), 
            .O(n6946)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3154_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_9 (.CI(n31425), .I0(n1252), .I1(VCC_net), .CO(n31426));
    SB_CARRY add_3154_4 (.CI(n30655), .I0(n1537), .I1(n98), .CO(n30656));
    SB_LUT4 rem_4_add_849_8_lut (.I0(GND_net), .I1(n1253), .I2(VCC_net), 
            .I3(n31424), .O(n1320)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3154_3_lut (.I0(GND_net), .I1(n1538), .I2(n99), .I3(n30654), 
            .O(n6947)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3154_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_8 (.CI(n31424), .I0(n1253), .I1(VCC_net), .CO(n31425));
    SB_CARRY add_3154_3 (.CI(n30654), .I0(n1538), .I1(n99), .CO(n30655));
    SB_LUT4 add_3154_2_lut (.I0(GND_net), .I1(n378), .I2(n558), .I3(VCC_net), 
            .O(n6948)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3154_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3154_2 (.CI(VCC_net), .I0(n378), .I1(n558), .CO(n30654));
    SB_LUT4 add_3152_11_lut (.I0(GND_net), .I1(n1412), .I2(n91), .I3(n30653), 
            .O(n6925)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3152_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3152_10_lut (.I0(GND_net), .I1(n1413), .I2(n92), .I3(n30652), 
            .O(n6926)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3152_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_849_7_lut (.I0(GND_net), .I1(n1254), .I2(GND_net), 
            .I3(n31423), .O(n1321)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3152_10 (.CI(n30652), .I0(n1413), .I1(n92), .CO(n30653));
    SB_LUT4 add_3152_9_lut (.I0(GND_net), .I1(n1414), .I2(n93), .I3(n30651), 
            .O(n6927)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3152_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3152_9 (.CI(n30651), .I0(n1414), .I1(n93), .CO(n30652));
    SB_LUT4 add_3152_8_lut (.I0(GND_net), .I1(n1415), .I2(n94), .I3(n30650), 
            .O(n6928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3152_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3152_8 (.CI(n30650), .I0(n1415), .I1(n94), .CO(n30651));
    SB_LUT4 add_3152_7_lut (.I0(GND_net), .I1(n1416), .I2(n95_adj_4360), 
            .I3(n30649), .O(n6929)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3152_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3152_7 (.CI(n30649), .I0(n1416), .I1(n95_adj_4360), .CO(n30650));
    SB_LUT4 add_3152_6_lut (.I0(GND_net), .I1(n1417), .I2(n96), .I3(n30648), 
            .O(n6930)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3152_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3152_6 (.CI(n30648), .I0(n1417), .I1(n96), .CO(n30649));
    SB_LUT4 add_3152_5_lut (.I0(GND_net), .I1(n1418), .I2(n97), .I3(n30647), 
            .O(n6931)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3152_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3152_5 (.CI(n30647), .I0(n1418), .I1(n97), .CO(n30648));
    SB_LUT4 add_3152_4_lut (.I0(GND_net), .I1(n1419), .I2(n98), .I3(n30646), 
            .O(n6932)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3152_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_7 (.CI(n31423), .I0(n1254), .I1(GND_net), .CO(n31424));
    SB_LUT4 rem_4_add_849_6_lut (.I0(GND_net), .I1(n1255), .I2(GND_net), 
            .I3(n31422), .O(n1322)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3152_4 (.CI(n30646), .I0(n1419), .I1(n98), .CO(n30647));
    SB_CARRY rem_4_add_849_6 (.CI(n31422), .I0(n1255), .I1(GND_net), .CO(n31423));
    SB_LUT4 add_3152_3_lut (.I0(GND_net), .I1(n1420), .I2(n99), .I3(n30645), 
            .O(n6933)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3152_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3152_3 (.CI(n30645), .I0(n1420), .I1(n99), .CO(n30646));
    SB_LUT4 add_3152_2_lut (.I0(GND_net), .I1(n377), .I2(n558), .I3(VCC_net), 
            .O(n6934)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3152_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3152_2 (.CI(VCC_net), .I0(n377), .I1(n558), .CO(n30645));
    SB_LUT4 add_3151_10_lut (.I0(GND_net), .I1(n1292), .I2(n92), .I3(n30644), 
            .O(n6914)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3151_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_849_5_lut (.I0(GND_net), .I1(n1256), .I2(VCC_net), 
            .I3(n31421), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3151_9_lut (.I0(GND_net), .I1(n1293), .I2(n93), .I3(n30643), 
            .O(n6915)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3151_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_5 (.CI(n31421), .I0(n1256), .I1(VCC_net), .CO(n31422));
    SB_LUT4 rem_4_add_849_4_lut (.I0(GND_net), .I1(n1257), .I2(VCC_net), 
            .I3(n31420), .O(n1324)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_4 (.CI(n31420), .I0(n1257), .I1(VCC_net), .CO(n31421));
    SB_CARRY add_3151_9 (.CI(n30643), .I0(n1293), .I1(n93), .CO(n30644));
    SB_LUT4 add_3151_8_lut (.I0(GND_net), .I1(n1294), .I2(n94), .I3(n30642), 
            .O(n6916)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3151_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3151_8 (.CI(n30642), .I0(n1294), .I1(n94), .CO(n30643));
    SB_LUT4 add_3151_7_lut (.I0(GND_net), .I1(n1295), .I2(n95_adj_4360), 
            .I3(n30641), .O(n6917)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3151_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_849_3_lut (.I0(GND_net), .I1(n1258), .I2(GND_net), 
            .I3(n31419), .O(n1325)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3151_7 (.CI(n30641), .I0(n1295), .I1(n95_adj_4360), .CO(n30642));
    SB_CARRY rem_4_add_849_3 (.CI(n31419), .I0(n1258), .I1(GND_net), .CO(n31420));
    SB_LUT4 add_3151_6_lut (.I0(GND_net), .I1(n1296), .I2(n96), .I3(n30640), 
            .O(n6918)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3151_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3151_6 (.CI(n30640), .I0(n1296), .I1(n96), .CO(n30641));
    SB_LUT4 div_36_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4559));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3151_5_lut (.I0(GND_net), .I1(n1297), .I2(n97), .I3(n30639), 
            .O(n6919)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3151_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_2 (.CI(VCC_net), .I0(n1358), .I1(VCC_net), 
            .CO(n31419));
    SB_CARRY add_3151_5 (.CI(n30639), .I0(n1297), .I1(n97), .CO(n30640));
    SB_LUT4 add_3151_4_lut (.I0(GND_net), .I1(n1298), .I2(n98), .I3(n30638), 
            .O(n6920)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3151_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3151_4 (.CI(n30638), .I0(n1298), .I1(n98), .CO(n30639));
    SB_LUT4 add_3151_3_lut (.I0(GND_net), .I1(n1299), .I2(n99), .I3(n30637), 
            .O(n6921)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3151_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3151_3 (.CI(n30637), .I0(n1299), .I1(n99), .CO(n30638));
    SB_LUT4 add_3151_2_lut (.I0(GND_net), .I1(n376), .I2(n558), .I3(VCC_net), 
            .O(n6922)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3151_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_916_12_lut (.I0(n1382), .I1(n1349), .I2(VCC_net), 
            .I3(n31418), .O(n1448)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_12_lut.LUT_INIT = 16'h8228;
    GND i1 (.Y(GND_net));
    SB_CARRY add_3151_2 (.CI(VCC_net), .I0(n376), .I1(n558), .CO(n30637));
    SB_LUT4 add_3150_9_lut (.I0(GND_net), .I1(n1169), .I2(n93), .I3(n30636), 
            .O(n6904)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3150_8_lut (.I0(GND_net), .I1(n1170), .I2(n94), .I3(n30635), 
            .O(n6905)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_916_11_lut (.I0(GND_net), .I1(n1350), .I2(VCC_net), 
            .I3(n31417), .O(n1417_adj_4496)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3150_8 (.CI(n30635), .I0(n1170), .I1(n94), .CO(n30636));
    SB_CARRY rem_4_add_916_11 (.CI(n31417), .I0(n1350), .I1(VCC_net), 
            .CO(n31418));
    SB_LUT4 add_3150_7_lut (.I0(GND_net), .I1(n1171), .I2(n95_adj_4360), 
            .I3(n30634), .O(n6906)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3150_7 (.CI(n30634), .I0(n1171), .I1(n95_adj_4360), .CO(n30635));
    SB_LUT4 add_3150_6_lut (.I0(GND_net), .I1(n1172), .I2(n96), .I3(n30633), 
            .O(n6907)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3150_6 (.CI(n30633), .I0(n1172), .I1(n96), .CO(n30634));
    SB_LUT4 add_3150_5_lut (.I0(GND_net), .I1(n1173), .I2(n97), .I3(n30632), 
            .O(n6908)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3150_5 (.CI(n30632), .I0(n1173), .I1(n97), .CO(n30633));
    SB_LUT4 add_3150_4_lut (.I0(GND_net), .I1(n1174), .I2(n98), .I3(n30631), 
            .O(n6909)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i1047_3_lut_3_lut (.I0(n1553), .I1(n6946), .I2(n1537), 
            .I3(GND_net), .O(n1651));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1047_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1045_3_lut_3_lut (.I0(n1553), .I1(n6944), .I2(n1535), 
            .I3(GND_net), .O(n1649));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1045_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3150_4 (.CI(n30631), .I0(n1174), .I1(n98), .CO(n30632));
    SB_LUT4 add_3150_3_lut (.I0(GND_net), .I1(n1175), .I2(n99), .I3(n30630), 
            .O(n6910)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3150_3 (.CI(n30630), .I0(n1175), .I1(n99), .CO(n30631));
    SB_LUT4 add_3150_2_lut (.I0(GND_net), .I1(n375), .I2(n558), .I3(VCC_net), 
            .O(n6911)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3150_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3150_2 (.CI(VCC_net), .I0(n375), .I1(n558), .CO(n30630));
    SB_LUT4 add_3149_8_lut (.I0(GND_net), .I1(n1043), .I2(n94), .I3(n30629), 
            .O(n6895)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3149_7_lut (.I0(GND_net), .I1(n1044), .I2(n95_adj_4360), 
            .I3(n30628), .O(n6896)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_916_10_lut (.I0(GND_net), .I1(n1351), .I2(VCC_net), 
            .I3(n31416), .O(n1418_adj_4497)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_7 (.CI(n30628), .I0(n1044), .I1(n95_adj_4360), .CO(n30629));
    SB_CARRY rem_4_add_916_10 (.CI(n31416), .I0(n1351), .I1(VCC_net), 
            .CO(n31417));
    SB_LUT4 add_3149_6_lut (.I0(GND_net), .I1(n1045), .I2(n96), .I3(n30627), 
            .O(n6897)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i1048_3_lut_3_lut (.I0(n1553), .I1(n6947), .I2(n1538), 
            .I3(GND_net), .O(n1652));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1048_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1042_3_lut_3_lut (.I0(n1553), .I1(n6941), .I2(n1532), 
            .I3(GND_net), .O(n1646));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1042_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3149_6 (.CI(n30627), .I0(n1045), .I1(n96), .CO(n30628));
    SB_LUT4 rem_4_add_916_9_lut (.I0(GND_net), .I1(n1352), .I2(VCC_net), 
            .I3(n31415), .O(n1419_adj_4498)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i1041_3_lut_3_lut (.I0(n1553), .I1(n6940), .I2(n1531), 
            .I3(GND_net), .O(n1645));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1041_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_3149_5_lut (.I0(GND_net), .I1(n1046), .I2(n97), .I3(n30626), 
            .O(n6898)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_5 (.CI(n30626), .I0(n1046), .I1(n97), .CO(n30627));
    SB_CARRY rem_4_add_916_9 (.CI(n31415), .I0(n1352), .I1(VCC_net), .CO(n31416));
    SB_LUT4 add_3149_4_lut (.I0(GND_net), .I1(n1047), .I2(n98), .I3(n30625), 
            .O(n6899)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i1049_3_lut_3_lut (.I0(n1553), .I1(n6948), .I2(n378), 
            .I3(GND_net), .O(n1653));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1049_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY add_3149_4 (.CI(n30625), .I0(n1047), .I1(n98), .CO(n30626));
    SB_LUT4 add_3149_3_lut (.I0(GND_net), .I1(n1048), .I2(n99), .I3(n30624), 
            .O(n6900)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_916_8_lut (.I0(GND_net), .I1(n1353), .I2(VCC_net), 
            .I3(n31414), .O(n1420_adj_4499)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_3 (.CI(n30624), .I0(n1048), .I1(n99), .CO(n30625));
    SB_LUT4 add_3149_2_lut (.I0(GND_net), .I1(n374), .I2(n558), .I3(VCC_net), 
            .O(n6901)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3149_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3149_2 (.CI(VCC_net), .I0(n374), .I1(n558), .CO(n30624));
    SB_LUT4 add_3148_7_lut (.I0(GND_net), .I1(n914), .I2(n95_adj_4360), 
            .I3(n30623), .O(n6887)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3148_6_lut (.I0(GND_net), .I1(n915), .I2(n96), .I3(n30622), 
            .O(n6888)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_8 (.CI(n31414), .I0(n1353), .I1(VCC_net), .CO(n31415));
    SB_CARRY add_3148_6 (.CI(n30622), .I0(n915), .I1(n96), .CO(n30623));
    SB_LUT4 add_3148_5_lut (.I0(GND_net), .I1(n916), .I2(n97), .I3(n30621), 
            .O(n6889)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_5 (.CI(n30621), .I0(n916), .I1(n97), .CO(n30622));
    SB_LUT4 add_3148_4_lut (.I0(GND_net), .I1(n917), .I2(n98), .I3(n30620), 
            .O(n6890)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_4 (.CI(n30620), .I0(n917), .I1(n98), .CO(n30621));
    SB_LUT4 rem_4_add_916_7_lut (.I0(GND_net), .I1(n1354), .I2(GND_net), 
            .I3(n31413), .O(n1421)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3148_3_lut (.I0(GND_net), .I1(n918), .I2(n99), .I3(n30619), 
            .O(n6891)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_3 (.CI(n30619), .I0(n918), .I1(n99), .CO(n30620));
    SB_CARRY rem_4_add_916_7 (.CI(n31413), .I0(n1354), .I1(GND_net), .CO(n31414));
    SB_LUT4 add_3148_2_lut (.I0(GND_net), .I1(n373), .I2(n558), .I3(VCC_net), 
            .O(n6892)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3148_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3148_2 (.CI(VCC_net), .I0(n373), .I1(n558), .CO(n30619));
    SB_LUT4 i24978_3_lut (.I0(n783), .I1(n97), .I2(n6_adj_4348), .I3(GND_net), 
            .O(n8_adj_4346));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i24978_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_36_i1044_3_lut_3_lut (.I0(n1553), .I1(n6943), .I2(n1534), 
            .I3(GND_net), .O(n1648));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1044_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1043_3_lut_3_lut (.I0(n1553), .I1(n6942), .I2(n1533), 
            .I3(GND_net), .O(n1647));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1043_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_6507_7_lut (.I0(GND_net), .I1(n3353), .I2(VCC_net), .I3(n30618), 
            .O(n11300)) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i1040_3_lut_3_lut (.I0(n1553), .I1(n6939), .I2(n1530), 
            .I3(GND_net), .O(n1644));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1040_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1039_3_lut_3_lut (.I0(n1553), .I1(n6938), .I2(n1529), 
            .I3(GND_net), .O(n1643));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1039_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 add_6507_6_lut (.I0(GND_net), .I1(n3354), .I2(GND_net), .I3(n30617), 
            .O(n11301)) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_916_6_lut (.I0(GND_net), .I1(n1355), .I2(GND_net), 
            .I3(n31412), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6507_6 (.CI(n30617), .I0(n3354), .I1(GND_net), .CO(n30618));
    SB_LUT4 i24970_3_lut (.I0(n784), .I1(n98), .I2(n4_adj_4349), .I3(GND_net), 
            .O(n6_adj_4348));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i24970_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 add_6507_5_lut (.I0(GND_net), .I1(n3355), .I2(GND_net), .I3(n30616), 
            .O(n11302)) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6507_5 (.CI(n30616), .I0(n3355), .I1(GND_net), .CO(n30617));
    SB_LUT4 i1_2_lut_adj_1713 (.I0(n2656), .I1(n2658), .I2(GND_net), .I3(GND_net), 
            .O(n40693));
    defparam i1_2_lut_adj_1713.LUT_INIT = 16'heeee;
    SB_LUT4 add_6507_4_lut (.I0(GND_net), .I1(n3356), .I2(VCC_net), .I3(n30615), 
            .O(n11303)) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6507_4 (.CI(n30615), .I0(n3356), .I1(VCC_net), .CO(n30616));
    SB_LUT4 add_6507_3_lut (.I0(GND_net), .I1(n3357), .I2(VCC_net), .I3(n30614), 
            .O(n11304)) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i1046_3_lut_3_lut (.I0(n1553), .I1(n6945), .I2(n1536), 
            .I3(GND_net), .O(n1650));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1046_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_916_6 (.CI(n31412), .I0(n1355), .I1(GND_net), .CO(n31413));
    SB_LUT4 rem_4_add_916_5_lut (.I0(GND_net), .I1(n1356), .I2(VCC_net), 
            .I3(n31411), .O(n1423)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6507_3 (.CI(n30614), .I0(n3357), .I1(VCC_net), .CO(n30615));
    SB_LUT4 add_6507_2_lut (.I0(GND_net), .I1(n3358), .I2(GND_net), .I3(VCC_net), 
            .O(n11305)) /* synthesis syn_instantiated=1 */ ;
    defparam add_6507_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6507_2 (.CI(VCC_net), .I0(n3358), .I1(GND_net), .CO(n30614));
    SB_CARRY rem_4_add_916_5 (.CI(n31411), .I0(n1356), .I1(VCC_net), .CO(n31412));
    SB_LUT4 rem_4_add_916_4_lut (.I0(GND_net), .I1(n1357), .I2(VCC_net), 
            .I3(n31410), .O(n1424)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_4 (.CI(n31410), .I0(n1357), .I1(VCC_net), .CO(n31411));
    SB_LUT4 i3_4_lut_adj_1714 (.I0(n3761), .I1(n6_adj_4626), .I2(n17264), 
            .I3(n46559), .O(n8_adj_4916));   // verilog/coms.v(126[12] 289[6])
    defparam i3_4_lut_adj_1714.LUT_INIT = 16'hcfce;
    SB_LUT4 rem_4_add_916_3_lut (.I0(GND_net), .I1(n1358), .I2(GND_net), 
            .I3(n31409), .O(n1425)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut_adj_1715 (.I0(n20639), .I1(n8_adj_4916), .I2(n17200), 
            .I3(n5_adj_4989), .O(n46050));   // verilog/coms.v(126[12] 289[6])
    defparam i4_4_lut_adj_1715.LUT_INIT = 16'hefcf;
    SB_CARRY rem_4_add_916_3 (.CI(n31409), .I0(n1358), .I1(GND_net), .CO(n31410));
    SB_CARRY rem_4_add_916_2 (.CI(VCC_net), .I0(n1458), .I1(VCC_net), 
            .CO(n31409));
    SB_LUT4 rem_4_add_983_13_lut (.I0(n1481), .I1(n1448), .I2(VCC_net), 
            .I3(n31408), .O(n1547)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_983_12_lut (.I0(GND_net), .I1(n1449), .I2(VCC_net), 
            .I3(n31407), .O(n1516)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_12 (.CI(n31407), .I0(n1449), .I1(VCC_net), 
            .CO(n31408));
    SB_LUT4 rem_4_add_983_11_lut (.I0(GND_net), .I1(n1450), .I2(VCC_net), 
            .I3(n31406), .O(n1517)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_11 (.CI(n31406), .I0(n1450), .I1(VCC_net), 
            .CO(n31407));
    SB_LUT4 div_36_LessThan_570_i45_2_lut (.I0(n915), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_570_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_983_10_lut (.I0(GND_net), .I1(n1451), .I2(VCC_net), 
            .I3(n31405), .O(n1518)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_10 (.CI(n31405), .I0(n1451), .I1(VCC_net), 
            .CO(n31406));
    SB_LUT4 rem_4_add_983_9_lut (.I0(GND_net), .I1(n1452), .I2(VCC_net), 
            .I3(n31404), .O(n1519)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_9 (.CI(n31404), .I0(n1452), .I1(VCC_net), .CO(n31405));
    SB_LUT4 rem_4_add_983_8_lut (.I0(GND_net), .I1(n1453), .I2(VCC_net), 
            .I3(n31403), .O(n1520)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_8 (.CI(n31403), .I0(n1453), .I1(VCC_net), .CO(n31404));
    SB_LUT4 rem_4_add_983_7_lut (.I0(GND_net), .I1(n1454), .I2(GND_net), 
            .I3(n31402), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_7 (.CI(n31402), .I0(n1454), .I1(GND_net), .CO(n31403));
    SB_LUT4 rem_4_add_983_6_lut (.I0(GND_net), .I1(n1455), .I2(GND_net), 
            .I3(n31401), .O(n1522)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_6 (.CI(n31401), .I0(n1455), .I1(GND_net), .CO(n31402));
    SB_LUT4 div_36_i1124_3_lut_3_lut (.I0(n1667), .I1(n6961), .I2(n1653), 
            .I3(GND_net), .O(n1764));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1124_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1123_3_lut_3_lut (.I0(n1667), .I1(n6960), .I2(n1652), 
            .I3(GND_net), .O(n1763));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1123_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_mux_3_i19_3_lut (.I0(encoder0_position[18]), .I1(n7_adj_4432), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n373));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1122_3_lut_3_lut (.I0(n1667), .I1(n6959), .I2(n1651), 
            .I3(GND_net), .O(n1762));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1122_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_983_5_lut (.I0(GND_net), .I1(n1456), .I2(VCC_net), 
            .I3(n31400), .O(n1523)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_5 (.CI(n31400), .I0(n1456), .I1(VCC_net), .CO(n31401));
    SB_LUT4 rem_4_add_983_4_lut (.I0(GND_net), .I1(n1457), .I2(VCC_net), 
            .I3(n31399), .O(n1524)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1716 (.I0(n2654), .I1(n40693), .I2(n2655), .I3(n2657), 
            .O(n38389));
    defparam i1_4_lut_adj_1716.LUT_INIT = 16'ha080;
    SB_CARRY rem_4_add_983_4 (.CI(n31399), .I0(n1457), .I1(VCC_net), .CO(n31400));
    SB_LUT4 div_36_i1121_3_lut_3_lut (.I0(n1667), .I1(n6958), .I2(n1650), 
            .I3(GND_net), .O(n1761));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1121_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1118_3_lut_3_lut (.I0(n1667), .I1(n6955), .I2(n1647), 
            .I3(GND_net), .O(n1758));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1118_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_983_3_lut (.I0(GND_net), .I1(n1458), .I2(GND_net), 
            .I3(n31398), .O(n1525)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_3 (.CI(n31398), .I0(n1458), .I1(GND_net), .CO(n31399));
    SB_CARRY rem_4_add_983_2 (.CI(VCC_net), .I0(n1558), .I1(VCC_net), 
            .CO(n31398));
    SB_LUT4 rem_4_add_1050_14_lut (.I0(n1580), .I1(n1547), .I2(VCC_net), 
            .I3(n31397), .O(n1646_adj_4481)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1050_13_lut (.I0(GND_net), .I1(n1548), .I2(VCC_net), 
            .I3(n31396), .O(n1615)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i1117_3_lut_3_lut (.I0(n1667), .I1(n6954), .I2(n1646), 
            .I3(GND_net), .O(n1757));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1117_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1125_3_lut_3_lut (.I0(n1667), .I1(n6962), .I2(n379), 
            .I3(GND_net), .O(n1765));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1125_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1050_13 (.CI(n31396), .I0(n1548), .I1(VCC_net), 
            .CO(n31397));
    SB_LUT4 rem_4_add_1050_12_lut (.I0(GND_net), .I1(n1549), .I2(VCC_net), 
            .I3(n31395), .O(n1616)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i24954_2_lut (.I0(n372), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_4434));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i24954_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY rem_4_add_1050_12 (.CI(n31395), .I0(n1549), .I1(VCC_net), 
            .CO(n31396));
    SB_LUT4 div_36_i1120_3_lut_3_lut (.I0(n1667), .I1(n6957), .I2(n1649), 
            .I3(GND_net), .O(n1760));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1120_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1050_11_lut (.I0(GND_net), .I1(n1550), .I2(VCC_net), 
            .I3(n31394), .O(n1617)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_36_i1119_3_lut_3_lut (.I0(n1667), .I1(n6956), .I2(n1648), 
            .I3(GND_net), .O(n1759));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1119_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1050_11 (.CI(n31394), .I0(n1550), .I1(VCC_net), 
            .CO(n31395));
    SB_DFF blink_43 (.Q(blink), .C(LED_c), .D(blink_N_255));   // verilog/TinyFPGA_B.v(48[8] 62[4])
    SB_LUT4 div_36_i572_1_lut (.I0(n938), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i572_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_570_i40_4_lut (.I0(n373), .I1(n99), .I2(n918), 
            .I3(n558), .O(n40_adj_4593));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_570_i40_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_36_LessThan_570_i44_3_lut (.I0(n42_adj_4594), .I1(n96), 
            .I2(n45), .I3(GND_net), .O(n44_adj_4595));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_570_i44_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i15_4_lut_adj_1717 (.I0(n2653), .I1(n30), .I2(n2637_adj_4492), 
            .I3(n2636_adj_4495), .O(n34));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i15_4_lut_adj_1717.LUT_INIT = 16'hfffe;
    SB_LUT4 i37258_4_lut (.I0(n44_adj_4595), .I1(n40_adj_4593), .I2(n45), 
            .I3(n43224), .O(n44383));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37258_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1718 (.I0(n44383), .I1(n17281), .I2(n95_adj_4360), 
            .I3(n914), .O(n938));
    defparam i1_4_lut_adj_1718.LUT_INIT = 16'hceef;
    SB_LUT4 div_36_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4558));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24938_3_lut (.I0(n648), .I1(n98), .I2(n4_adj_4443), .I3(GND_net), 
            .O(n6_adj_4438));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i24938_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_36_i1115_3_lut_3_lut (.I0(n1667), .I1(n6952), .I2(n1644), 
            .I3(GND_net), .O(n1755));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1115_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14345_3_lut (.I0(encoder0_position[23]), .I1(n2866), .I2(count_enable), 
            .I3(GND_net), .O(n19377));   // quad.v(35[10] 41[6])
    defparam i14345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1116_3_lut_3_lut (.I0(n1667), .I1(n6953), .I2(n1645), 
            .I3(GND_net), .O(n1756));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1116_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_mux_3_i20_3_lut (.I0(encoder0_position[19]), .I1(n6_adj_4431), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n372));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24922_2_lut (.I0(n371), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_4907));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i24922_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_36_i483_1_lut (.I0(n806), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i483_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_481_i42_4_lut (.I0(n372), .I1(n99), .I2(n785), 
            .I3(n558), .O(n42_adj_4592));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_481_i42_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i37524_3_lut (.I0(n42_adj_4592), .I1(n98), .I2(n784), .I3(GND_net), 
            .O(n44649));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37524_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i37525_3_lut (.I0(n44649), .I1(n97), .I2(n783), .I3(GND_net), 
            .O(n44650));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37525_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1719 (.I0(n44650), .I1(n17278), .I2(n96), .I3(n38026), 
            .O(n806));
    defparam i1_4_lut_adj_1719.LUT_INIT = 16'hefce;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i1_1_lut (.I0(communication_counter[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n33_adj_4969));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24898_2_lut (.I0(n370), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_4601));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i24898_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_36_mux_3_i21_3_lut (.I0(encoder0_position[20]), .I1(n5_adj_4358), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n371));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i392_1_lut (.I0(n671), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n672));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i392_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_390_i44_4_lut (.I0(n371), .I1(n99), .I2(n649), 
            .I3(n558), .O(n44));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_390_i44_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i37502_3_lut (.I0(n44), .I1(n98), .I2(n648), .I3(GND_net), 
            .O(n44627));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37502_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1720 (.I0(n44627), .I1(n17275), .I2(n97), .I3(n38024), 
            .O(n671));
    defparam i1_4_lut_adj_1720.LUT_INIT = 16'hefce;
    SB_LUT4 div_36_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4557));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24882_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i24882_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_36_mux_3_i22_3_lut (.I0(encoder0_position[21]), .I1(n4_adj_4326), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n370));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i299_1_lut (.I0(n533), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n534));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i299_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_297_i46_4_lut (.I0(n370), .I1(n99), .I2(n510), 
            .I3(n558), .O(n46));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_297_i46_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i1_4_lut_adj_1721 (.I0(n46), .I1(n17272), .I2(n98), .I3(n38022), 
            .O(n533));
    defparam i1_4_lut_adj_1721.LUT_INIT = 16'hefce;
    SB_LUT4 i1_4_lut_adj_1722 (.I0(n224), .I1(n99), .I2(n17269), .I3(n558), 
            .O(n5_adj_4915));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i1_4_lut_adj_1722.LUT_INIT = 16'h555d;
    SB_LUT4 div_36_mux_3_i23_3_lut (.I0(encoder0_position[22]), .I1(n3), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n369));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i204_1_lut (.I0(n392), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i204_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_i1114_3_lut_3_lut (.I0(n1667), .I1(n6951), .I2(n1643), 
            .I3(GND_net), .O(n1754));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1114_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i36070_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n42871));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36070_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_4_lut_adj_1723 (.I0(n42871), .I1(n17269), .I2(n99), .I3(n5_adj_4915), 
            .O(n392));
    defparam i1_4_lut_adj_1723.LUT_INIT = 16'hefce;
    SB_LUT4 div_36_i1197_3_lut_3_lut (.I0(n1778), .I1(n6975), .I2(n1764), 
            .I3(GND_net), .O(n1872));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1197_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_mux_5_i23_3_lut (.I0(gearBoxRatio[22]), .I1(n53), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n78));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1724 (.I0(n78), .I1(n77), .I2(GND_net), .I3(GND_net), 
            .O(n17244));
    defparam i1_2_lut_adj_1724.LUT_INIT = 16'hdddd;
    SB_LUT4 div_36_i1187_3_lut_3_lut (.I0(n1778), .I1(n6965), .I2(n1754), 
            .I3(GND_net), .O(n1862));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1187_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_mux_5_i22_3_lut (.I0(gearBoxRatio[21]), .I1(n54), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n79));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_36_mux_5_i21_3_lut (.I0(gearBoxRatio[20]), .I1(n55), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n80));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_36_mux_5_i20_3_lut (.I0(gearBoxRatio[19]), .I1(n56), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n81));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1725 (.I0(n81), .I1(n17236), .I2(GND_net), .I3(GND_net), 
            .O(n17311));
    defparam i1_2_lut_adj_1725.LUT_INIT = 16'hdddd;
    SB_LUT4 div_36_mux_5_i19_3_lut (.I0(gearBoxRatio[18]), .I1(n57), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n82));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_36_mux_5_i18_3_lut (.I0(gearBoxRatio[17]), .I1(n58), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n83));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_36_mux_5_i17_3_lut (.I0(gearBoxRatio[16]), .I1(n59), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n84));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i13_4_lut_adj_1726 (.I0(n2645), .I1(n2651), .I2(n2649), .I3(n2646), 
            .O(n32));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i13_4_lut_adj_1726.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1727 (.I0(n84), .I1(n17231), .I2(GND_net), .I3(GND_net), 
            .O(n17305));
    defparam i1_2_lut_adj_1727.LUT_INIT = 16'hdddd;
    SB_LUT4 div_36_i1196_3_lut_3_lut (.I0(n1778), .I1(n6974), .I2(n1763), 
            .I3(GND_net), .O(n1871));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1196_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_mux_5_i16_3_lut (.I0(gearBoxRatio[15]), .I1(n60), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n85));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_36_mux_5_i15_3_lut (.I0(gearBoxRatio[14]), .I1(n61), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n86));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i14344_3_lut (.I0(encoder0_position[22]), .I1(n2867), .I2(count_enable), 
            .I3(GND_net), .O(n19376));   // quad.v(35[10] 41[6])
    defparam i14344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14343_3_lut (.I0(encoder0_position[21]), .I1(n2868), .I2(count_enable), 
            .I3(GND_net), .O(n19375));   // quad.v(35[10] 41[6])
    defparam i14343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14342_3_lut (.I0(encoder0_position[20]), .I1(n2869), .I2(count_enable), 
            .I3(GND_net), .O(n19374));   // quad.v(35[10] 41[6])
    defparam i14342_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_mux_5_i14_3_lut (.I0(gearBoxRatio[13]), .I1(n62), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n87));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1728 (.I0(n87), .I1(n17225), .I2(GND_net), .I3(GND_net), 
            .O(n17299));
    defparam i1_2_lut_adj_1728.LUT_INIT = 16'hdddd;
    SB_LUT4 div_36_mux_5_i13_3_lut (.I0(gearBoxRatio[12]), .I1(n63), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n88));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_36_mux_5_i12_3_lut (.I0(gearBoxRatio[11]), .I1(n64), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n89));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_36_i1195_3_lut_3_lut (.I0(n1778), .I1(n6973), .I2(n1762), 
            .I3(GND_net), .O(n1870));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1195_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_mux_5_i11_3_lut (.I0(gearBoxRatio[10]), .I1(n65), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n90));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1729 (.I0(n90), .I1(n17293), .I2(GND_net), .I3(GND_net), 
            .O(n17211));
    defparam i1_2_lut_adj_1729.LUT_INIT = 16'hdddd;
    SB_LUT4 div_36_mux_5_i10_3_lut (.I0(gearBoxRatio[9]), .I1(n66), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n91));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_36_mux_5_i9_3_lut (.I0(gearBoxRatio[8]), .I1(n67), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n92));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_36_mux_5_i8_3_lut (.I0(gearBoxRatio[7]), .I1(n68), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n93));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1730 (.I0(n93), .I1(n17287), .I2(GND_net), .I3(GND_net), 
            .O(n17284));
    defparam i1_2_lut_adj_1730.LUT_INIT = 16'hdddd;
    SB_LUT4 div_36_mux_5_i7_3_lut (.I0(gearBoxRatio[6]), .I1(n69), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n94));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_36_mux_5_i6_3_lut (.I0(gearBoxRatio[5]), .I1(n70), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n95_adj_4360));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_36_mux_5_i5_3_lut (.I0(gearBoxRatio[4]), .I1(n71), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n96));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1731 (.I0(n96), .I1(n17278), .I2(GND_net), .I3(GND_net), 
            .O(n17275));
    defparam i1_2_lut_adj_1731.LUT_INIT = 16'hdddd;
    SB_LUT4 div_36_mux_5_i4_3_lut (.I0(gearBoxRatio[3]), .I1(n72), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n97));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_36_mux_5_i3_3_lut (.I0(gearBoxRatio[2]), .I1(n73), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n98));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_36_mux_5_i2_3_lut (.I0(gearBoxRatio[1]), .I1(n74), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n99));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_36_mux_5_i1_3_lut (.I0(gearBoxRatio[0]), .I1(n75), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n558));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_5_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i2_4_lut_adj_1732 (.I0(n558), .I1(n99), .I2(n224), .I3(n17269), 
            .O(n248));
    defparam i2_4_lut_adj_1732.LUT_INIT = 16'hff37;
    SB_LUT4 div_36_i1198_3_lut_3_lut (.I0(n1778), .I1(n6976), .I2(n1765), 
            .I3(GND_net), .O(n1873));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1198_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i38739_2_lut (.I0(encoder0_position[23]), .I1(gearBoxRatio[23]), 
            .I2(GND_net), .I3(GND_net), .O(n45862));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i38739_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i2_1_lut (.I0(communication_counter[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_4968));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4556));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i3_1_lut (.I0(communication_counter[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_4967));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4555));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i4_1_lut (.I0(communication_counter[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_4966));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4554));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i5_1_lut (.I0(communication_counter[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_4965));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4553));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i6_1_lut (.I0(communication_counter[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_4964));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_i1194_3_lut_3_lut (.I0(n1778), .I1(n6972), .I2(n1761), 
            .I3(GND_net), .O(n1869));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1194_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4552));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i7_1_lut (.I0(communication_counter[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_4963));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4551));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i8_1_lut (.I0(communication_counter[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_4962));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i9_1_lut (.I0(communication_counter[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4961));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4550));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i10_1_lut (.I0(communication_counter[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4960));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4549));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i11_1_lut (.I0(communication_counter[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4959));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4548));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13823_4_lut (.I0(n18584), .I1(state[1]), .I2(state_3__N_362[1]), 
            .I3(n18416), .O(n18855));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13823_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i13824_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n39307), .I3(GND_net), .O(n18856));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13824_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13825_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n39307), .I3(GND_net), .O(n18857));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13825_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14_4_lut_adj_1733 (.I0(n2652), .I1(n2650), .I2(n2647), .I3(n2648), 
            .O(n33));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i14_4_lut_adj_1733.LUT_INIT = 16'hfffe;
    SB_LUT4 i13826_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n39307), .I3(GND_net), .O(n18858));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13826_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13827_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n39307), .I3(GND_net), .O(n18859));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13827_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14354_3_lut (.I0(encoder1_position[8]), .I1(n2831), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19386));   // quad.v(35[10] 41[6])
    defparam i14354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14353_3_lut (.I0(encoder1_position[7]), .I1(n2832), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19385));   // quad.v(35[10] 41[6])
    defparam i14353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1734 (.I0(n2642_adj_4490), .I1(n2644), .I2(n2643_adj_4489), 
            .I3(n38389), .O(n31));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i12_4_lut_adj_1734.LUT_INIT = 16'hfffe;
    SB_LUT4 i13828_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n39307), .I3(GND_net), .O(n18860));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13828_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14352_3_lut (.I0(encoder1_position[6]), .I1(n2833), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19384));   // quad.v(35[10] 41[6])
    defparam i14352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13829_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n39307), .I3(GND_net), .O(n18861));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13829_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13830_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n39307), .I3(GND_net), .O(n18862));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13830_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14351_3_lut (.I0(encoder1_position[5]), .I1(n2834), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19383));   // quad.v(35[10] 41[6])
    defparam i14351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18_4_lut_adj_1735 (.I0(n31), .I1(n33), .I2(n32), .I3(n34), 
            .O(n2669));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i18_4_lut_adj_1735.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i12_1_lut (.I0(communication_counter[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4958));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4547));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13831_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n39307), .I3(GND_net), .O(n18863));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13831_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13832_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n39307), .I3(GND_net), .O(n18864));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13832_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13833_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n39307), .I3(GND_net), .O(n18865));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13833_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13834_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n39307), .I3(GND_net), .O(n18866));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13834_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13835_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n39307), .I3(GND_net), .O(n18867));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13835_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13836_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n39307), .I3(GND_net), .O(n18868));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13837_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n39307), .I3(GND_net), .O(n18869));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13838_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n39307), .I3(GND_net), .O(n18870));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13839_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n39307), .I3(GND_net), .O(n18871));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13840_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n39307), .I3(GND_net), .O(n18872));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13841_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n39307), .I3(GND_net), .O(n18873));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13842_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n39307), .I3(GND_net), .O(n18874));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_i1192_3_lut_3_lut (.I0(n1778), .I1(n6970), .I2(n1759), 
            .I3(GND_net), .O(n1867));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1192_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13843_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n39307), .I3(GND_net), .O(n18875));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13844_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n39307), .I3(GND_net), .O(n18876));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i13_1_lut (.I0(communication_counter[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4957));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13845_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n39307), .I3(GND_net), .O(n18877));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13846_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n39307), .I3(GND_net), .O(n18878));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13846_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13847_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n39307), .I3(GND_net), .O(n18879));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13847_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13848_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n39307), .I3(GND_net), .O(n18880));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13849_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n39307), .I3(GND_net), .O(n18881));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13850_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n39307), .I3(GND_net), .O(n18882));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13851_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n39307), .I3(GND_net), .O(n18883));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13851_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13852_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n39307), .I3(GND_net), .O(n18884));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13852_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13853_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n39307), .I3(GND_net), .O(n18885));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13853_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4546));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i14_1_lut (.I0(communication_counter[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4956));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4545));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i15_1_lut (.I0(communication_counter[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4955));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i16_1_lut (.I0(communication_counter[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4954));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i17_1_lut (.I0(communication_counter[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4953));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i18_1_lut (.I0(communication_counter[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4952));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i19_1_lut (.I0(communication_counter[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4951));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i20_1_lut (.I0(communication_counter[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4950));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_i1193_3_lut_3_lut (.I0(n1778), .I1(n6971), .I2(n1760), 
            .I3(GND_net), .O(n1868));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1193_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1199_3_lut_3_lut (.I0(n1778), .I1(n6977), .I2(n380), 
            .I3(GND_net), .O(n1874));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1199_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13854_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n39307), .I3(GND_net), .O(n18886));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13854_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_i1191_3_lut_3_lut (.I0(n1778), .I1(n6969), .I2(n1758), 
            .I3(GND_net), .O(n1866));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1191_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13866_2_lut (.I0(n18897), .I1(n18896), .I2(GND_net), .I3(GND_net), 
            .O(n18898));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13866_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24_3_lut (.I0(n42939), .I1(bit_ctr[27]), .I2(n4754), .I3(GND_net), 
            .O(n35915));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1190_3_lut_3_lut (.I0(n1778), .I1(n6968), .I2(n1757), 
            .I3(GND_net), .O(n1865));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1190_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_mux_3_i10_3_lut (.I0(communication_counter[9]), .I1(n24_adj_4386), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2658));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1934_3_lut (.I0(n2845), .I1(n2912), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2944));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1937_3_lut (.I0(n2848), .I1(n2915), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2947));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1937_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1939_3_lut (.I0(n2850), .I1(n2917), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2949));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1941_3_lut (.I0(n2852), .I1(n2919), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2951));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1938_3_lut (.I0(n2849), .I1(n2916), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2948));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1940_3_lut (.I0(n2851), .I1(n2918), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2950));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1936_3_lut (.I0(n2847), .I1(n2914), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2946));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1936_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1189_3_lut_3_lut (.I0(n1778), .I1(n6967), .I2(n1756), 
            .I3(GND_net), .O(n1864));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1189_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1943_3_lut (.I0(n2854), .I1(n2921), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2953));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1935_3_lut (.I0(n2846), .I1(n2913), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2945));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1942_3_lut (.I0(n2853), .I1(n2920), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2952));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1188_3_lut_3_lut (.I0(n1778), .I1(n6966), .I2(n1755), 
            .I3(GND_net), .O(n1863));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1188_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1933_3_lut (.I0(n2844), .I1(n2911), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2943));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1932_3_lut (.I0(n2843), .I1(n2910), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2942));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1926_3_lut (.I0(n2837_adj_4448), .I1(n2904), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2936));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1925_3_lut (.I0(n2836_adj_4449), .I1(n2903), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2935));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1924_3_lut (.I0(n2835_adj_4450), .I1(n2902), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2934));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1930_3_lut (.I0(n2841), .I1(n2908), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2940));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1928_3_lut (.I0(n2839_adj_4446), .I1(n2906), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2938));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1929_3_lut (.I0(n2840), .I1(n2907), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2939));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1927_3_lut (.I0(n2838_adj_4447), .I1(n2905), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2937));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1945_3_lut (.I0(n2856), .I1(n2923), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2955));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1944_3_lut (.I0(n2855), .I1(n2922), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2954));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1931_3_lut (.I0(n2842), .I1(n2909), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2941));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i7_3_lut (.I0(communication_counter[6]), .I1(n27_adj_4381), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2958));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1947_3_lut (.I0(n2858), .I1(n2925), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2957));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1946_3_lut (.I0(n2857_adj_4442), .I1(n2924), .I2(n2867_adj_4441), 
            .I3(GND_net), .O(n2956));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1736 (.I0(n2956), .I1(n2957), .I2(n2958), .I3(GND_net), 
            .O(n38343));
    defparam i1_3_lut_adj_1736.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_4_lut_adj_1737 (.I0(n2941), .I1(n2954), .I2(n38343), .I3(n2955), 
            .O(n27));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i5_4_lut_adj_1737.LUT_INIT = 16'heaaa;
    SB_LUT4 div_36_i1270_3_lut_3_lut (.I0(n1886), .I1(n6992), .I2(n1874), 
            .I3(GND_net), .O(n1979));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1270_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13_4_lut_adj_1738 (.I0(n2937), .I1(n2939), .I2(n2938), .I3(n2940), 
            .O(n35));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i13_4_lut_adj_1738.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1739 (.I0(n2934), .I1(n2935), .I2(n2933), .I3(n2936), 
            .O(n34_adj_4347));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i12_4_lut_adj_1739.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1740 (.I0(n35), .I1(n27), .I2(n2942), .I3(n2943), 
            .O(n40));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i18_4_lut_adj_1740.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1741 (.I0(n2952), .I1(n2945), .I2(n2953), .I3(n2946), 
            .O(n38));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i16_4_lut_adj_1741.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2950), .I1(n34_adj_4347), .I2(n2948), .I3(GND_net), 
            .O(n39));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1742 (.I0(n2951), .I1(n2949), .I2(n2947), .I3(n2944), 
            .O(n37));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i15_4_lut_adj_1742.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(n37), .I1(n39), .I2(n38), .I3(n40), .O(n2966));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14362_3_lut (.I0(encoder1_position[16]), .I1(n2823), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19394));   // quad.v(35[10] 41[6])
    defparam i14362_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1260_3_lut_3_lut (.I0(n1886), .I1(n6982), .I2(n1864), 
            .I3(GND_net), .O(n1969));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1260_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14361_3_lut (.I0(encoder1_position[15]), .I1(n2824), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19393));   // quad.v(35[10] 41[6])
    defparam i14361_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1743 (.I0(bit_ctr[0]), .I1(n42940), .I2(n4754), 
            .I3(GND_net), .O(n35917));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1743.LUT_INIT = 16'hacac;
    SB_LUT4 i24_3_lut_adj_1744 (.I0(n42936), .I1(bit_ctr[26]), .I2(n4754), 
            .I3(GND_net), .O(n35913));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1744.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i21_1_lut (.I0(communication_counter[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4949));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i22_1_lut (.I0(communication_counter[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4948));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i23_1_lut (.I0(communication_counter[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4947));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i24_1_lut (.I0(communication_counter[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4946));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_i1259_3_lut_3_lut (.I0(n1886), .I1(n6981), .I2(n1863), 
            .I3(GND_net), .O(n1968));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1259_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1258_3_lut_3_lut (.I0(n1886), .I1(n6980), .I2(n1862), 
            .I3(GND_net), .O(n1967));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1258_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i25_1_lut (.I0(communication_counter[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4945));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13906_3_lut (.I0(color[17]), .I1(n23_adj_4362), .I2(n15_adj_4367), 
            .I3(GND_net), .O(n18938));   // verilog/TinyFPGA_B.v(48[8] 62[4])
    defparam i13906_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13907_3_lut (.I0(color[20]), .I1(n23_adj_4362), .I2(n15_adj_4367), 
            .I3(GND_net), .O(n18939));   // verilog/TinyFPGA_B.v(48[8] 62[4])
    defparam i13907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i26_1_lut (.I0(communication_counter[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4944));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_2_lut_adj_1745 (.I0(color_23__N_164[3]), .I1(color_23__N_164[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4341));   // verilog/TinyFPGA_B.v(51[6:36])
    defparam i3_2_lut_adj_1745.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1746 (.I0(color_23__N_164[4]), .I1(color_23__N_164[6]), 
            .I2(color_23__N_164[2]), .I3(color_23__N_164[0]), .O(n13_adj_4340));   // verilog/TinyFPGA_B.v(51[6:36])
    defparam i1_4_lut_adj_1746.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1747 (.I0(color_23__N_164[7]), .I1(n13_adj_4340), 
            .I2(n11_adj_4341), .I3(color_23__N_164[1]), .O(n15_adj_4367));   // verilog/TinyFPGA_B.v(51[6:36])
    defparam i1_4_lut_adj_1747.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1748 (.I0(color_23__N_164[1]), .I1(blink), .I2(GND_net), 
            .I3(GND_net), .O(n40281));   // verilog/TinyFPGA_B.v(51[6:36])
    defparam i1_2_lut_adj_1748.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1749 (.I0(color_23__N_164[7]), .I1(n13_adj_4340), 
            .I2(n11_adj_4341), .I3(n40281), .O(n23_adj_4362));   // verilog/TinyFPGA_B.v(51[6:36])
    defparam i1_4_lut_adj_1749.LUT_INIT = 16'hfffe;
    SB_LUT4 i13908_3_lut (.I0(color[21]), .I1(n23_adj_4362), .I2(n15_adj_4367), 
            .I3(GND_net), .O(n18940));   // verilog/TinyFPGA_B.v(48[8] 62[4])
    defparam i13908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13911_3_lut (.I0(n18602), .I1(r_Bit_Index[0]), .I2(n18467), 
            .I3(GND_net), .O(n18943));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13911_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 div_36_i1269_3_lut_3_lut (.I0(n1886), .I1(n6991), .I2(n1873), 
            .I3(GND_net), .O(n1978));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1269_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1267_3_lut_3_lut (.I0(n1886), .I1(n6989), .I2(n1871), 
            .I3(GND_net), .O(n1976));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1267_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_LessThan_1722_i12_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2631), 
            .I3(GND_net), .O(n12_adj_4833));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i27_1_lut (.I0(communication_counter[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4943));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_1722_i10_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2636), 
            .I3(GND_net), .O(n10_adj_4831));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_36_LessThan_1722_i14_3_lut_3_lut (.I0(n95_adj_4360), .I1(n94), 
            .I2(n2633), .I3(GND_net), .O(n14_adj_4835));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_36_i1268_3_lut_3_lut (.I0(n1886), .I1(n6990), .I2(n1872), 
            .I3(GND_net), .O(n1977));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1268_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35942_2_lut_4_lut (.I0(n2623), .I1(n84), .I2(n2632), .I3(n93), 
            .O(n43066));
    defparam i35942_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_36_LessThan_1722_i16_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2623), 
            .I3(GND_net), .O(n16_adj_4837));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i35977_2_lut_4_lut (.I0(n2631), .I1(n92), .I2(n2635), .I3(n96), 
            .O(n43101));
    defparam i35977_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_36_LessThan_1777_i8_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2718), 
            .I3(GND_net), .O(n8_adj_4857));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i8_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_36_i1265_3_lut_3_lut (.I0(n1886), .I1(n6987), .I2(n1869), 
            .I3(GND_net), .O(n1974));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1265_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1266_3_lut_3_lut (.I0(n1886), .I1(n6988), .I2(n1870), 
            .I3(GND_net), .O(n1975));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1266_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1264_3_lut_3_lut (.I0(n1886), .I1(n6986), .I2(n1868), 
            .I3(GND_net), .O(n1973));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1264_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1271_3_lut_3_lut (.I0(n1886), .I1(n6993), .I2(n381), 
            .I3(GND_net), .O(n1980));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1271_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1263_3_lut_3_lut (.I0(n1886), .I1(n6985), .I2(n1867), 
            .I3(GND_net), .O(n1972));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1263_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1262_3_lut_3_lut (.I0(n1886), .I1(n6984), .I2(n1866), 
            .I3(GND_net), .O(n1971));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1262_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14374_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n39036), 
            .I3(GND_net), .O(n19406));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i14374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1750 (.I0(bit_ctr[22]), .I1(n42944), .I2(n4754), 
            .I3(GND_net), .O(n35929));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1750.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_i1261_3_lut_3_lut (.I0(n1886), .I1(n6983), .I2(n1865), 
            .I3(GND_net), .O(n1970));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1261_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1340_3_lut_3_lut (.I0(n1991), .I1(n7009), .I2(n1980), 
            .I3(GND_net), .O(n2082));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1340_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1332_3_lut_3_lut (.I0(n1991), .I1(n7001), .I2(n1972), 
            .I3(GND_net), .O(n2074));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1332_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1331_3_lut_3_lut (.I0(n1991), .I1(n7000), .I2(n1971), 
            .I3(GND_net), .O(n2073));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1331_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1330_3_lut_3_lut (.I0(n1991), .I1(n6999), .I2(n1970), 
            .I3(GND_net), .O(n2072));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1330_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1328_3_lut_3_lut (.I0(n1991), .I1(n6997), .I2(n1968), 
            .I3(GND_net), .O(n2070));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1328_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_LessThan_1777_i12_3_lut_3_lut (.I0(n95_adj_4360), .I1(n94), 
            .I2(n2715), .I3(GND_net), .O(n12_adj_4861));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i36593_2_lut_4_lut (.I0(n2705), .I1(n84), .I2(n2714), .I3(n93), 
            .O(n43718));
    defparam i36593_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_36_i1329_3_lut_3_lut (.I0(n1991), .I1(n6998), .I2(n1969), 
            .I3(GND_net), .O(n2071));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1329_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_LessThan_1777_i14_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2705), 
            .I3(GND_net), .O(n14_adj_4863));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_36_i1327_3_lut_3_lut (.I0(n1991), .I1(n6996), .I2(n1967), 
            .I3(GND_net), .O(n2069));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1327_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1338_3_lut_3_lut (.I0(n1991), .I1(n7007), .I2(n1978), 
            .I3(GND_net), .O(n2080));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1338_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_LessThan_1777_i10_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2713), 
            .I3(GND_net), .O(n10_adj_4859));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_36_i1339_3_lut_3_lut (.I0(n1991), .I1(n7008), .I2(n1979), 
            .I3(GND_net), .O(n2081));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1339_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13723_2_lut (.I0(n18897), .I1(n18753), .I2(GND_net), .I3(GND_net), 
            .O(n18755));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13723_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_36_i1337_3_lut_3_lut (.I0(n1991), .I1(n7006), .I2(n1977), 
            .I3(GND_net), .O(n2079));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1337_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35904_2_lut_4_lut (.I0(n2713), .I1(n92), .I2(n2717), .I3(n96), 
            .O(n43028));
    defparam i35904_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i22_3_lut_adj_1751 (.I0(bit_ctr[13]), .I1(n42964), .I2(n4754), 
            .I3(GND_net), .O(n35971));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1751.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_i1336_3_lut_3_lut (.I0(n1991), .I1(n7005), .I2(n1976), 
            .I3(GND_net), .O(n2078));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1336_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i38704_4_lut (.I0(r_SM_Main[2]), .I1(n42919), .I2(n42920), 
            .I3(r_SM_Main[1]), .O(n27445));
    defparam i38704_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 div_36_i1335_3_lut_3_lut (.I0(n1991), .I1(n7004), .I2(n1975), 
            .I3(GND_net), .O(n2077));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1335_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1334_3_lut_3_lut (.I0(n1991), .I1(n7003), .I2(n1974), 
            .I3(GND_net), .O(n2076));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1334_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i24_3_lut_adj_1752 (.I0(n42935), .I1(bit_ctr[25]), .I2(n4754), 
            .I3(GND_net), .O(n35911));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1752.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4423));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_i1341_3_lut_3_lut (.I0(n1991), .I1(n7010), .I2(n382), 
            .I3(GND_net), .O(n2083));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1341_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14382_3_lut (.I0(\half_duty[0] [1]), .I1(half_duty_new[1]), 
            .I2(n1111), .I3(GND_net), .O(n19414));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i14382_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i24_3_lut_adj_1753 (.I0(n42934), .I1(bit_ctr[24]), .I2(n4754), 
            .I3(GND_net), .O(n35909));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1753.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1333_3_lut_3_lut (.I0(n1991), .I1(n7002), .I2(n1973), 
            .I3(GND_net), .O(n2075));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1333_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i38017_1_lut_2_lut (.I0(n3362), .I1(n11300), .I2(GND_net), 
            .I3(GND_net), .O(n45142));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i38017_1_lut_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_36_i1407_3_lut_3_lut (.I0(n2093), .I1(n7026), .I2(n2082), 
            .I3(GND_net), .O(n2181));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1407_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1400_3_lut_3_lut (.I0(n2093), .I1(n7019), .I2(n2075), 
            .I3(GND_net), .O(n2174));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1400_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13995_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position[17]), 
            .I2(n14536), .I3(GND_net), .O(n19027));   // verilog/coms.v(126[12] 289[6])
    defparam i13995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13996_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position[18]), 
            .I2(n14536), .I3(GND_net), .O(n19028));   // verilog/coms.v(126[12] 289[6])
    defparam i13996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13997_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position[19]), 
            .I2(n14536), .I3(GND_net), .O(n19029));   // verilog/coms.v(126[12] 289[6])
    defparam i13997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13998_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position[20]), 
            .I2(n14536), .I3(GND_net), .O(n19030));   // verilog/coms.v(126[12] 289[6])
    defparam i13998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1409_3_lut_3_lut (.I0(n2093), .I1(n7028), .I2(n383), 
            .I3(GND_net), .O(n2183));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1409_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1397_3_lut_3_lut (.I0(n2093), .I1(n7016), .I2(n2072), 
            .I3(GND_net), .O(n2171));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1397_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1396_3_lut_3_lut (.I0(n2093), .I1(n7015), .I2(n2071), 
            .I3(GND_net), .O(n2170));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1396_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1395_3_lut_3_lut (.I0(n2093), .I1(n7014), .I2(n2070), 
            .I3(GND_net), .O(n2169));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1395_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 displacement_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4422));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_i1398_3_lut_3_lut (.I0(n2093), .I1(n7017), .I2(n2073), 
            .I3(GND_net), .O(n2172));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1398_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13999_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position[21]), 
            .I2(n14536), .I3(GND_net), .O(n19031));   // verilog/coms.v(126[12] 289[6])
    defparam i13999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14233_3_lut (.I0(\data_in_frame[15] [0]), .I1(rx_data[0]), 
            .I2(n37348), .I3(GND_net), .O(n19265));   // verilog/coms.v(126[12] 289[6])
    defparam i14233_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14000_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position[22]), 
            .I2(n14536), .I3(GND_net), .O(n19032));   // verilog/coms.v(126[12] 289[6])
    defparam i14000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14001_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position[23]), 
            .I2(n14536), .I3(GND_net), .O(n19033));   // verilog/coms.v(126[12] 289[6])
    defparam i14001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1394_3_lut_3_lut (.I0(n2093), .I1(n7013), .I2(n2069), 
            .I3(GND_net), .O(n2168));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1394_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14002_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position[8]), 
            .I2(n14536), .I3(GND_net), .O(n19034));   // verilog/coms.v(126[12] 289[6])
    defparam i14002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14003_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position[9]), 
            .I2(n14536), .I3(GND_net), .O(n19035));   // verilog/coms.v(126[12] 289[6])
    defparam i14003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14004_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position[10]), 
            .I2(n14536), .I3(GND_net), .O(n19036));   // verilog/coms.v(126[12] 289[6])
    defparam i14004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14393_3_lut (.I0(\half_duty[0] [7]), .I1(half_duty_new[7]), 
            .I2(n1111), .I3(GND_net), .O(n19425));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i14393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1406_3_lut_3_lut (.I0(n2093), .I1(n7025), .I2(n2081), 
            .I3(GND_net), .O(n2180));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1406_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14392_3_lut (.I0(\half_duty[0] [6]), .I1(half_duty_new[6]), 
            .I2(n1111), .I3(GND_net), .O(n19424));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i14392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1405_3_lut_3_lut (.I0(n2093), .I1(n7024), .I2(n2080), 
            .I3(GND_net), .O(n2179));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1405_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1404_3_lut_3_lut (.I0(n2093), .I1(n7023), .I2(n2079), 
            .I3(GND_net), .O(n2178));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1404_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1403_3_lut_3_lut (.I0(n2093), .I1(n7022), .I2(n2078), 
            .I3(GND_net), .O(n2177));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1403_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1402_3_lut_3_lut (.I0(n2093), .I1(n7021), .I2(n2077), 
            .I3(GND_net), .O(n2176));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1402_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1408_3_lut_3_lut (.I0(n2093), .I1(n7027), .I2(n2083), 
            .I3(GND_net), .O(n2182));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1408_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1401_3_lut_3_lut (.I0(n2093), .I1(n7020), .I2(n2076), 
            .I3(GND_net), .O(n2175));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1401_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14005_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position[11]), 
            .I2(n14536), .I3(GND_net), .O(n19037));   // verilog/coms.v(126[12] 289[6])
    defparam i14005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1399_3_lut_3_lut (.I0(n2093), .I1(n7018), .I2(n2074), 
            .I3(GND_net), .O(n2173));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1399_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14391_3_lut (.I0(\half_duty[0] [5]), .I1(half_duty_new[5]), 
            .I2(n1111), .I3(GND_net), .O(n19423));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i14391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1754 (.I0(blink), .I1(n15_adj_4367), .I2(GND_net), 
            .I3(GND_net), .O(blink_N_255));
    defparam i1_2_lut_adj_1754.LUT_INIT = 16'h9999;
    SB_LUT4 mux_61_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[0]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14234_3_lut (.I0(\data_in_frame[15] [1]), .I1(rx_data[1]), 
            .I2(n37348), .I3(GND_net), .O(n19266));   // verilog/coms.v(126[12] 289[6])
    defparam i14234_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14006_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position[12]), 
            .I2(n14536), .I3(GND_net), .O(n19038));   // verilog/coms.v(126[12] 289[6])
    defparam i14006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4421));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14390_3_lut (.I0(\half_duty[0] [4]), .I1(half_duty_new[4]), 
            .I2(n1111), .I3(GND_net), .O(n19422));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i14390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14389_3_lut (.I0(\half_duty[0] [3]), .I1(half_duty_new[3]), 
            .I2(n1111), .I3(GND_net), .O(n19421));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i14389_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_60_i1_3_lut (.I0(encoder0_position[0]), .I1(motor_state_23__N_106[0]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14007_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position[13]), 
            .I2(n14536), .I3(GND_net), .O(n19039));   // verilog/coms.v(126[12] 289[6])
    defparam i14007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14008_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position[14]), 
            .I2(n14536), .I3(GND_net), .O(n19040));   // verilog/coms.v(126[12] 289[6])
    defparam i14008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14388_3_lut (.I0(\half_duty[0] [2]), .I1(half_duty_new[2]), 
            .I2(n1111), .I3(GND_net), .O(n19420));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i14388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_61_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[1]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i2_3_lut (.I0(encoder0_position[1]), .I1(motor_state_23__N_106[1]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14009_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position[15]), 
            .I2(n14536), .I3(GND_net), .O(n19041));   // verilog/coms.v(126[12] 289[6])
    defparam i14009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14169_3_lut (.I0(\data_in_frame[7] [0]), .I1(rx_data[0]), .I2(n37368), 
            .I3(GND_net), .O(n19201));   // verilog/coms.v(126[12] 289[6])
    defparam i14169_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_61_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[2]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i3_3_lut (.I0(encoder0_position[2]), .I1(motor_state_23__N_106[2]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_61_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[3]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i4_3_lut (.I0(encoder0_position[3]), .I1(motor_state_23__N_106[3]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14010_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position[0]), 
            .I2(n14536), .I3(GND_net), .O(n19042));   // verilog/coms.v(126[12] 289[6])
    defparam i14010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_61_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[4]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 displacement_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4420));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_60_i5_3_lut (.I0(encoder0_position[4]), .I1(motor_state_23__N_106[4]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14235_3_lut (.I0(\data_in_frame[15] [2]), .I1(rx_data[2]), 
            .I2(n37348), .I3(GND_net), .O(n19267));   // verilog/coms.v(126[12] 289[6])
    defparam i14235_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14387_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4), .I3(n17255), 
            .O(n19419));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i14387_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14170_3_lut (.I0(\data_in_frame[7] [1]), .I1(rx_data[1]), .I2(n37368), 
            .I3(GND_net), .O(n19202));   // verilog/coms.v(126[12] 289[6])
    defparam i14170_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1755 (.I0(bit_ctr[16]), .I1(n42943), .I2(n4754), 
            .I3(GND_net), .O(n35927));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1755.LUT_INIT = 16'hacac;
    SB_LUT4 i13631_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n39307), .I3(GND_net), .O(n18663));   // verilog/neopixel.v(35[12] 117[6])
    defparam i13631_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i24_3_lut_adj_1756 (.I0(n42933), .I1(bit_ctr[23]), .I2(n4754), 
            .I3(GND_net), .O(n35907));   // verilog/neopixel.v(35[12] 117[6])
    defparam i24_3_lut_adj_1756.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_61_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[5]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i6_3_lut (.I0(encoder0_position[5]), .I1(motor_state_23__N_106[5]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_61_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[6]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i7_3_lut (.I0(encoder0_position[6]), .I1(motor_state_23__N_106[6]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4419));   // verilog/TinyFPGA_B.v(243[21:79])
    defparam displacement_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_61_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[7]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i8_3_lut (.I0(encoder0_position[7]), .I1(motor_state_23__N_106[7]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1669_3_lut (.I0(n2452_adj_4581), .I1(n2519), .I2(n2471_adj_4574), 
            .I3(GND_net), .O(n2551_adj_4511));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14401_3_lut (.I0(setpoint[7]), .I1(n4666), .I2(n39863), .I3(GND_net), 
            .O(n19433));   // verilog/coms.v(126[12] 289[6])
    defparam i14401_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_i107_1_lut_4_lut (.I0(n558), .I1(n99), .I2(n224), .I3(n17269), 
            .O(n249));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i107_1_lut_4_lut.LUT_INIT = 16'h00c8;
    SB_LUT4 i1_2_lut_4_lut (.I0(n98), .I1(n97), .I2(n96), .I3(n17278), 
            .O(n17269));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 mux_61_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[8]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i9_3_lut (.I0(encoder0_position[8]), .I1(motor_state_23__N_106[8]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14400_3_lut (.I0(setpoint[6]), .I1(n4665), .I2(n39863), .I3(GND_net), 
            .O(n19432));   // verilog/coms.v(126[12] 289[6])
    defparam i14400_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut_adj_1757 (.I0(n97), .I1(n96), .I2(n17278), 
            .I3(GND_net), .O(n17272));
    defparam i1_2_lut_3_lut_adj_1757.LUT_INIT = 16'hf7f7;
    SB_LUT4 mux_61_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[9]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i10_3_lut (.I0(encoder0_position[9]), .I1(motor_state_23__N_106[9]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i1_3_lut (.I0(communication_counter[0]), .I1(n33_adj_4376), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3459));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_61_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[10]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i11_3_lut (.I0(encoder0_position[10]), .I1(motor_state_23__N_106[10]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14411_3_lut (.I0(setpoint[17]), .I1(n4676), .I2(n39863), 
            .I3(GND_net), .O(n19443));   // verilog/coms.v(126[12] 289[6])
    defparam i14411_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_mux_3_i2_3_lut (.I0(communication_counter[1]), .I1(n32_adj_4377), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3458));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 mux_61_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[11]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i12_3_lut (.I0(encoder0_position[11]), .I1(motor_state_23__N_106[11]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38033_1_lut (.I0(n3457), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45158));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i38033_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2287_3_lut (.I0(n3358), .I1(n11305), .I2(n3362), .I3(GND_net), 
            .O(n3457));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2287_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i38030_1_lut (.I0(n3456), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45155));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i38030_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2286_3_lut (.I0(n3357), .I1(n11304), .I2(n3362), .I3(GND_net), 
            .O(n3456));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2286_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i38027_1_lut (.I0(n3455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45152));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i38027_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2285_3_lut (.I0(n3356), .I1(n11303), .I2(n3362), .I3(GND_net), 
            .O(n3455));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2285_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i25_4_lut (.I0(n27365), .I1(n38070), .I2(state[0]), .I3(n17195), 
            .O(n11_adj_4911));   // verilog/neopixel.v(35[12] 117[6])
    defparam i25_4_lut.LUT_INIT = 16'h303a;
    SB_LUT4 mux_61_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[12]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i13_3_lut (.I0(encoder0_position[12]), .I1(motor_state_23__N_106[12]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i38024_1_lut (.I0(n3454), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45149));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i38024_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2284_3_lut (.I0(n3355), .I1(n11302), .I2(n3362), .I3(GND_net), 
            .O(n3454));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2284_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i38021_1_lut (.I0(n3453), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45146));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i38021_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2283_3_lut (.I0(n3354), .I1(n11301), .I2(n3362), .I3(GND_net), 
            .O(n3453));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2283_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_i2215_3_lut (.I0(n3254), .I1(n3321), .I2(n3263), .I3(GND_net), 
            .O(n3353));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2219_3_lut (.I0(n3258), .I1(n3325), .I2(n3263), .I3(GND_net), 
            .O(n3357));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2217_3_lut (.I0(n3256), .I1(n3323), .I2(n3263), .I3(GND_net), 
            .O(n3355));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2216_3_lut (.I0(n3255), .I1(n3322), .I2(n3263), .I3(GND_net), 
            .O(n3354));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i3_3_lut (.I0(communication_counter[2]), .I1(n31_adj_4378), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3358));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2218_3_lut (.I0(n3257), .I1(n3324), .I2(n3263), .I3(GND_net), 
            .O(n3356));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2206_3_lut (.I0(n3245), .I1(n3312), .I2(n3263), .I3(GND_net), 
            .O(n3344));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2204_3_lut (.I0(n3243), .I1(n3310), .I2(n3263), .I3(GND_net), 
            .O(n3342));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1758 (.I0(n3246), .I1(n3342), .I2(n3313), .I3(n3263), 
            .O(n40301));
    defparam i1_4_lut_adj_1758.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_2_lut_adj_1759 (.I0(n3356), .I1(n3358), .I2(GND_net), .I3(GND_net), 
            .O(n40673));
    defparam i1_2_lut_adj_1759.LUT_INIT = 16'heeee;
    SB_LUT4 rem_4_i2208_3_lut (.I0(n3247), .I1(n3314), .I2(n3263), .I3(GND_net), 
            .O(n3346));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2213_3_lut (.I0(n3252), .I1(n3319), .I2(n3263), .I3(GND_net), 
            .O(n3351));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1760 (.I0(n3249), .I1(n3351), .I2(n3316), .I3(n3263), 
            .O(n40377));
    defparam i1_4_lut_adj_1760.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1761 (.I0(n40377), .I1(n3251), .I2(n3318), .I3(n3263), 
            .O(n40379));
    defparam i1_4_lut_adj_1761.LUT_INIT = 16'hfaee;
    SB_LUT4 i1_4_lut_adj_1762 (.I0(n3242), .I1(n40379), .I2(n3309), .I3(n3263), 
            .O(n40381));
    defparam i1_4_lut_adj_1762.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1763 (.I0(n3240), .I1(n40381), .I2(n3307), .I3(n3263), 
            .O(n40383));
    defparam i1_4_lut_adj_1763.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1764 (.I0(n3239), .I1(n40383), .I2(n3306), .I3(n3263), 
            .O(n40385));
    defparam i1_4_lut_adj_1764.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1765 (.I0(n3244), .I1(n3344), .I2(n3311), .I3(n3263), 
            .O(n40299));
    defparam i1_4_lut_adj_1765.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1766 (.I0(n40301), .I1(n3253), .I2(n3320), .I3(n3263), 
            .O(n40303));
    defparam i1_4_lut_adj_1766.LUT_INIT = 16'hfaee;
    SB_LUT4 i1_4_lut_adj_1767 (.I0(n3354), .I1(n40673), .I2(n3355), .I3(n3357), 
            .O(n38358));
    defparam i1_4_lut_adj_1767.LUT_INIT = 16'ha080;
    SB_LUT4 rem_4_i2202_3_lut (.I0(n3241), .I1(n3308), .I2(n3263), .I3(GND_net), 
            .O(n3340));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14410_3_lut (.I0(setpoint[16]), .I1(n4675), .I2(n39863), 
            .I3(GND_net), .O(n19442));   // verilog/coms.v(126[12] 289[6])
    defparam i14410_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1768 (.I0(n3340), .I1(n38358), .I2(n40303), .I3(n40299), 
            .O(n40309));
    defparam i1_4_lut_adj_1768.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1769 (.I0(n3237), .I1(n40309), .I2(n3304), .I3(n3263), 
            .O(n40311));
    defparam i1_4_lut_adj_1769.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1770 (.I0(n3236), .I1(n40385), .I2(n3303), .I3(n3263), 
            .O(n40387));
    defparam i1_4_lut_adj_1770.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1771 (.I0(n3353), .I1(n3250), .I2(n3317), .I3(n3263), 
            .O(n40397));
    defparam i1_4_lut_adj_1771.LUT_INIT = 16'hfaee;
    SB_LUT4 i3_4_lut_adj_1772 (.I0(n3248), .I1(n3346), .I2(n3315), .I3(n3263), 
            .O(n28_adj_5005));
    defparam i3_4_lut_adj_1772.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1773 (.I0(n40387), .I1(n3235), .I2(n3302), .I3(n3263), 
            .O(n46_adj_5004));
    defparam i1_4_lut_adj_1773.LUT_INIT = 16'hfaee;
    SB_LUT4 i1_4_lut_adj_1774 (.I0(n40311), .I1(n3233), .I2(n3300), .I3(n3263), 
            .O(n47_adj_5003));
    defparam i1_4_lut_adj_1774.LUT_INIT = 16'hfaee;
    SB_LUT4 rem_4_i2199_3_lut (.I0(n3238), .I1(n3305), .I2(n3263), .I3(GND_net), 
            .O(n3337));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1775 (.I0(n3234), .I1(n3337), .I2(n3301), .I3(n3263), 
            .O(n40019));
    defparam i1_4_lut_adj_1775.LUT_INIT = 16'hfcee;
    SB_LUT4 rem_4_i2192_3_lut (.I0(n3231), .I1(n3298), .I2(n3263), .I3(GND_net), 
            .O(n3330));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1776 (.I0(n47_adj_5003), .I1(n46_adj_5004), .I2(n28_adj_5005), 
            .I3(n40397), .O(n40403));
    defparam i1_4_lut_adj_1776.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1777 (.I0(n3232), .I1(n40019), .I2(n3299), .I3(n3263), 
            .O(n40021));
    defparam i1_4_lut_adj_1777.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1778 (.I0(n40712), .I1(n40021), .I2(n40403), 
            .I3(n3330), .O(n3362));
    defparam i1_4_lut_adj_1778.LUT_INIT = 16'hfffe;
    SB_LUT4 i38020_2_lut (.I0(n3362), .I1(n11300), .I2(GND_net), .I3(GND_net), 
            .O(n3452));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i38020_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i14409_3_lut (.I0(setpoint[15]), .I1(n4674), .I2(n39863), 
            .I3(GND_net), .O(n19441));   // verilog/coms.v(126[12] 289[6])
    defparam i14409_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_i1468_3_lut_3_lut (.I0(n2192), .I1(n7040), .I2(n2177), 
            .I3(GND_net), .O(n2273));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1468_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut_adj_1779 (.I0(n95_adj_4360), .I1(n94), .I2(n93), 
            .I3(n17287), .O(n17278));
    defparam i1_2_lut_4_lut_adj_1779.LUT_INIT = 16'hff7f;
    SB_LUT4 div_36_i1459_3_lut_3_lut (.I0(n2192), .I1(n7031), .I2(n2168), 
            .I3(GND_net), .O(n2264));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1459_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut_adj_1780 (.I0(n94), .I1(n93), .I2(n17287), 
            .I3(GND_net), .O(n17281));
    defparam i1_2_lut_3_lut_adj_1780.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_36_i1469_3_lut_3_lut (.I0(n2192), .I1(n7041), .I2(n2178), 
            .I3(GND_net), .O(n2274));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1469_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut_adj_1781 (.I0(n92), .I1(n91), .I2(n90), .I3(n17293), 
            .O(n17287));
    defparam i1_2_lut_4_lut_adj_1781.LUT_INIT = 16'hff7f;
    SB_LUT4 i14341_3_lut (.I0(encoder0_position[19]), .I1(n2870), .I2(count_enable), 
            .I3(GND_net), .O(n19373));   // quad.v(35[10] 41[6])
    defparam i14341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1473_3_lut_3_lut (.I0(n2192), .I1(n7045), .I2(n2182), 
            .I3(GND_net), .O(n2278));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1473_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut_adj_1782 (.I0(n91), .I1(n90), .I2(n17293), 
            .I3(GND_net), .O(n17290));
    defparam i1_2_lut_3_lut_adj_1782.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1783 (.I0(n89), .I1(n88), .I2(n87), .I3(n17225), 
            .O(n17293));
    defparam i1_2_lut_4_lut_adj_1783.LUT_INIT = 16'hff7f;
    SB_LUT4 div_36_i1472_3_lut_3_lut (.I0(n2192), .I1(n7044), .I2(n2181), 
            .I3(GND_net), .O(n2277));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1472_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 unary_minus_18_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24_adj_4338));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_i1475_3_lut_3_lut (.I0(n2192), .I1(n7047), .I2(n384), 
            .I3(GND_net), .O(n2280));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1475_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_61_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[13]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i14_3_lut (.I0(encoder0_position[13]), .I1(motor_state_23__N_106[13]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1463_3_lut_3_lut (.I0(n2192), .I1(n7035), .I2(n2172), 
            .I3(GND_net), .O(n2268));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1463_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 unary_minus_18_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4337));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14340_3_lut (.I0(encoder0_position[18]), .I1(n2871), .I2(count_enable), 
            .I3(GND_net), .O(n19372));   // quad.v(35[10] 41[6])
    defparam i14340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14413_3_lut (.I0(setpoint[19]), .I1(n4678), .I2(n39863), 
            .I3(GND_net), .O(n19445));   // verilog/coms.v(126[12] 289[6])
    defparam i14413_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_i1462_3_lut_3_lut (.I0(n2192), .I1(n7034), .I2(n2171), 
            .I3(GND_net), .O(n2267));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1462_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut_adj_1784 (.I0(n88), .I1(n87), .I2(n17225), 
            .I3(GND_net), .O(n17296));
    defparam i1_2_lut_3_lut_adj_1784.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1785 (.I0(n86), .I1(n85), .I2(n84), .I3(n17231), 
            .O(n17225));
    defparam i1_2_lut_4_lut_adj_1785.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1786 (.I0(n85), .I1(n84), .I2(n17231), 
            .I3(GND_net), .O(n17302));
    defparam i1_2_lut_3_lut_adj_1786.LUT_INIT = 16'hf7f7;
    SB_LUT4 i14412_3_lut (.I0(setpoint[18]), .I1(n4677), .I2(n39863), 
            .I3(GND_net), .O(n19444));   // verilog/coms.v(126[12] 289[6])
    defparam i14412_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_i1461_3_lut_3_lut (.I0(n2192), .I1(n7033), .I2(n2170), 
            .I3(GND_net), .O(n2266));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1461_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 unary_minus_18_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22_adj_4336));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_61_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[14]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i15_3_lut (.I0(encoder0_position[14]), .I1(motor_state_23__N_106[14]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1464_3_lut_3_lut (.I0(n2192), .I1(n7036), .I2(n2173), 
            .I3(GND_net), .O(n2269));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1464_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1460_3_lut_3_lut (.I0(n2192), .I1(n7032), .I2(n2169), 
            .I3(GND_net), .O(n2265));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1460_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut_adj_1787 (.I0(n83), .I1(n82), .I2(n81), .I3(n17236), 
            .O(n17231));
    defparam i1_2_lut_4_lut_adj_1787.LUT_INIT = 16'hff7f;
    SB_LUT4 unary_minus_18_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4335));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_61_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[15]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i16_3_lut (.I0(encoder0_position[15]), .I1(motor_state_23__N_106[15]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1470_3_lut_3_lut (.I0(n2192), .I1(n7042), .I2(n2179), 
            .I3(GND_net), .O(n2275));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1470_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut_adj_1788 (.I0(n82), .I1(n81), .I2(n17236), 
            .I3(GND_net), .O(n17308));
    defparam i1_2_lut_3_lut_adj_1788.LUT_INIT = 16'hf7f7;
    SB_LUT4 mux_61_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[16]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i17_3_lut (.I0(encoder0_position[16]), .I1(motor_state_23__N_106[16]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14415_3_lut (.I0(setpoint[21]), .I1(n4680), .I2(n39863), 
            .I3(GND_net), .O(n19447));   // verilog/coms.v(126[12] 289[6])
    defparam i14415_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_i1471_3_lut_3_lut (.I0(n2192), .I1(n7043), .I2(n2180), 
            .I3(GND_net), .O(n2276));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1471_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1474_3_lut_3_lut (.I0(n2192), .I1(n7046), .I2(n2183), 
            .I3(GND_net), .O(n2279));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1474_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_61_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[17]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 div_36_i1467_3_lut_3_lut (.I0(n2192), .I1(n7039), .I2(n2176), 
            .I3(GND_net), .O(n2272));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1467_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_60_i18_3_lut (.I0(encoder0_position[17]), .I1(motor_state_23__N_106[17]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1465_3_lut_3_lut (.I0(n2192), .I1(n7037), .I2(n2174), 
            .I3(GND_net), .O(n2270));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1465_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut_adj_1789 (.I0(n80), .I1(n79), .I2(n78), .I3(n77), 
            .O(n17236));
    defparam i1_2_lut_4_lut_adj_1789.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1790 (.I0(n79), .I1(n78), .I2(n77), .I3(GND_net), 
            .O(n17241));
    defparam i1_2_lut_3_lut_adj_1790.LUT_INIT = 16'hf7f7;
    SB_LUT4 i24906_3_lut_4_lut (.I0(n510), .I1(n99), .I2(n370), .I3(n558), 
            .O(n4_adj_4339));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i24906_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i24930_3_lut_4_lut (.I0(n649), .I1(n99), .I2(n371), .I3(n558), 
            .O(n4_adj_4443));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i24930_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i24962_3_lut_4_lut (.I0(n785), .I1(n99), .I2(n372), .I3(n558), 
            .O(n4_adj_4349));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i24962_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 div_36_i1466_3_lut_3_lut (.I0(n2192), .I1(n7038), .I2(n2175), 
            .I3(GND_net), .O(n2271));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1466_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_LessThan_985_i32_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1536), 
            .I3(GND_net), .O(n32_adj_4630));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_985_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i14414_3_lut (.I0(setpoint[20]), .I1(n4679), .I2(n39863), 
            .I3(GND_net), .O(n19446));   // verilog/coms.v(126[12] 289[6])
    defparam i14414_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35946_2_lut_4_lut (.I0(n1531), .I1(n92), .I2(n1535), .I3(n96), 
            .O(n43070));
    defparam i35946_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i14417_3_lut (.I0(setpoint[23]), .I1(n4682), .I2(n39863), 
            .I3(GND_net), .O(n19449));   // verilog/coms.v(126[12] 289[6])
    defparam i14417_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_18_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18_adj_4334));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_985_i34_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1531), 
            .I3(GND_net), .O(n34_adj_4632));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_985_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 rem_4_i586_rep_55_3_lut_4_lut (.I0(n40223), .I1(n746), .I2(n12167), 
            .I3(n749), .O(n956));
    defparam rem_4_i586_rep_55_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mux_61_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[18]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i19_3_lut (.I0(encoder0_position[18]), .I1(motor_state_23__N_106[18]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i587_3_lut_4_lut (.I0(n40223), .I1(n746), .I2(n12168), 
            .I3(n855), .O(n957));
    defparam rem_4_i587_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 rem_4_i585_3_lut_4_lut (.I0(n40223), .I1(n746), .I2(n12166), 
            .I3(n748), .O(n955));
    defparam rem_4_i585_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mux_61_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[19]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i20_3_lut (.I0(encoder0_position[19]), .I1(motor_state_23__N_106[19]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i584_3_lut_4_lut (.I0(n40223), .I1(n746), .I2(n12165), 
            .I3(n852), .O(n954));
    defparam rem_4_i584_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i14416_3_lut (.I0(setpoint[22]), .I1(n4681), .I2(n39863), 
            .I3(GND_net), .O(n19448));   // verilog/coms.v(126[12] 289[6])
    defparam i14416_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_i1530_3_lut_3_lut (.I0(n2288), .I1(n7058), .I2(n2272), 
            .I3(GND_net), .O(n2365));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1530_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 unary_minus_18_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4333));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_61_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[20]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i22_3_lut_adj_1791 (.I0(bit_ctr[21]), .I1(n42942), .I2(n4754), 
            .I3(GND_net), .O(n35925));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1791.LUT_INIT = 16'hacac;
    SB_LUT4 mux_60_i21_3_lut (.I0(encoder0_position[20]), .I1(motor_state_23__N_106[20]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1522_3_lut_3_lut (.I0(n2288), .I1(n7050), .I2(n2264), 
            .I3(GND_net), .O(n2357));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1522_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1525_3_lut_3_lut (.I0(n2288), .I1(n7053), .I2(n2267), 
            .I3(GND_net), .O(n2360));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1525_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1523_3_lut_3_lut (.I0(n2288), .I1(n7051), .I2(n2265), 
            .I3(GND_net), .O(n2358));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1523_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1526_3_lut_3_lut (.I0(n2288), .I1(n7054), .I2(n2268), 
            .I3(GND_net), .O(n2361));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1526_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14418_3_lut (.I0(quadA_debounced_adj_4372), .I1(reg_B_adj_5057[1]), 
            .I2(n39886), .I3(GND_net), .O(n19450));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i14418_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2141_3_lut (.I0(n3148), .I1(n3215), .I2(n3164), .I3(GND_net), 
            .O(n3247));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2140_3_lut (.I0(n3147), .I1(n3214), .I2(n3164), .I3(GND_net), 
            .O(n3246));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2135_3_lut (.I0(n3142), .I1(n3209), .I2(n3164), .I3(GND_net), 
            .O(n3241));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2134_3_lut (.I0(n3141), .I1(n3208), .I2(n3164), .I3(GND_net), 
            .O(n3240));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1062_i30_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1651), 
            .I3(GND_net), .O(n30_adj_4642));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1062_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 rem_4_i2129_3_lut (.I0(n3136), .I1(n3203), .I2(n3164), .I3(GND_net), 
            .O(n3235));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2127_3_lut (.I0(n3134), .I1(n3201), .I2(n3164), .I3(GND_net), 
            .O(n3233));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1532_3_lut_3_lut (.I0(n2288), .I1(n7060), .I2(n2274), 
            .I3(GND_net), .O(n2367));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1532_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i2128_3_lut (.I0(n3135), .I1(n3202), .I2(n3164), .I3(GND_net), 
            .O(n3234));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2126_3_lut (.I0(n3133), .I1(n3200), .I2(n3164), .I3(GND_net), 
            .O(n3232));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2138_3_lut (.I0(n3145), .I1(n3212), .I2(n3164), .I3(GND_net), 
            .O(n3244));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35920_2_lut_4_lut (.I0(n1646), .I1(n92), .I2(n1650), .I3(n96), 
            .O(n43044));
    defparam i35920_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 rem_4_i2144_3_lut (.I0(n3151), .I1(n3218), .I2(n3164), .I3(GND_net), 
            .O(n3250));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2147_3_lut (.I0(n3154), .I1(n3221), .I2(n3164), .I3(GND_net), 
            .O(n3253));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2142_3_lut (.I0(n3149), .I1(n3216), .I2(n3164), .I3(GND_net), 
            .O(n3248));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2133_3_lut (.I0(n3140), .I1(n3207), .I2(n3164), .I3(GND_net), 
            .O(n3239));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1062_i32_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1646), 
            .I3(GND_net), .O(n32_adj_4644));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1062_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i14360_3_lut (.I0(encoder1_position[14]), .I1(n2825), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19392));   // quad.v(35[10] 41[6])
    defparam i14360_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1538_3_lut_3_lut (.I0(n2288), .I1(n7066), .I2(n2280), 
            .I3(GND_net), .O(n2373));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1538_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14359_3_lut (.I0(encoder1_position[13]), .I1(n2826), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19391));   // quad.v(35[10] 41[6])
    defparam i14359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2131_3_lut (.I0(n3138), .I1(n3205), .I2(n3164), .I3(GND_net), 
            .O(n3237));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1537_3_lut_3_lut (.I0(n2288), .I1(n7065), .I2(n2279), 
            .I3(GND_net), .O(n2372));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1537_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i2132_3_lut (.I0(n3139), .I1(n3206), .I2(n3164), .I3(GND_net), 
            .O(n3238));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2130_3_lut (.I0(n3137), .I1(n3204), .I2(n3164), .I3(GND_net), 
            .O(n3236));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2125_3_lut (.I0(n3132), .I1(n3199), .I2(n3164), .I3(GND_net), 
            .O(n3231));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2139_3_lut (.I0(n3146), .I1(n3213), .I2(n3164), .I3(GND_net), 
            .O(n3245));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2145_3_lut (.I0(n3152), .I1(n3219), .I2(n3164), .I3(GND_net), 
            .O(n3251));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2137_3_lut (.I0(n3144), .I1(n3211), .I2(n3164), .I3(GND_net), 
            .O(n3243));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1536_3_lut_3_lut (.I0(n2288), .I1(n7064), .I2(n2278), 
            .I3(GND_net), .O(n2371));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1536_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i2143_3_lut (.I0(n3150), .I1(n3217), .I2(n3164), .I3(GND_net), 
            .O(n3249));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2146_3_lut (.I0(n3153), .I1(n3220), .I2(n3164), .I3(GND_net), 
            .O(n3252));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2149_3_lut (.I0(n3156), .I1(n3223), .I2(n3164), .I3(GND_net), 
            .O(n3255));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14358_3_lut (.I0(encoder1_position[12]), .I1(n2827), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19390));   // quad.v(35[10] 41[6])
    defparam i14358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2136_3_lut (.I0(n3143), .I1(n3210), .I2(n3164), .I3(GND_net), 
            .O(n3242));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2148_3_lut (.I0(n3155), .I1(n3222), .I2(n3164), .I3(GND_net), 
            .O(n3254));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i4_3_lut (.I0(communication_counter[3]), .I1(n30_adj_4379), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3258));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2151_3_lut (.I0(n3158), .I1(n3225), .I2(n3164), .I3(GND_net), 
            .O(n3257));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14357_3_lut (.I0(encoder1_position[11]), .I1(n2828), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19389));   // quad.v(35[10] 41[6])
    defparam i14357_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2150_3_lut (.I0(n3157), .I1(n3224), .I2(n3164), .I3(GND_net), 
            .O(n3256));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14356_3_lut (.I0(encoder1_position[10]), .I1(n2829), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19388));   // quad.v(35[10] 41[6])
    defparam i14356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1792 (.I0(n3256), .I1(n3257), .I2(n3258), .I3(GND_net), 
            .O(n38410));
    defparam i1_3_lut_adj_1792.LUT_INIT = 16'hfefe;
    SB_LUT4 i7_4_lut_adj_1793 (.I0(n3254), .I1(n3242), .I2(n38410), .I3(n3255), 
            .O(n32_adj_4982));
    defparam i7_4_lut_adj_1793.LUT_INIT = 16'heccc;
    SB_LUT4 i14355_3_lut (.I0(encoder1_position[9]), .I1(n2830), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19387));   // quad.v(35[10] 41[6])
    defparam i14355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17_4_lut_adj_1794 (.I0(n3252), .I1(n3249), .I2(n3243), .I3(n3251), 
            .O(n42_adj_4978));
    defparam i17_4_lut_adj_1794.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n3245), .I1(n3231), .I2(n3230), .I3(GND_net), 
            .O(n38_adj_4981));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut_adj_1795 (.I0(n3248), .I1(n3253), .I2(n3250), .I3(n3244), 
            .O(n43_adj_4977));
    defparam i18_4_lut_adj_1795.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1796 (.I0(n3236), .I1(n3238), .I2(n3237), .I3(n3239), 
            .O(n40_adj_4979));
    defparam i15_4_lut_adj_1796.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1797 (.I0(n3240), .I1(n42_adj_4978), .I2(n32_adj_4982), 
            .I3(n3241), .O(n46_adj_4976));
    defparam i21_4_lut_adj_1797.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1798 (.I0(n3232), .I1(n3234), .I2(n3233), .I3(n3235), 
            .O(n39_adj_4980));
    defparam i14_4_lut_adj_1798.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n43_adj_4977), .I1(n3246), .I2(n38_adj_4981), 
            .I3(n3247), .O(n47));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n47), .I1(n39_adj_4980), .I2(n46_adj_4976), 
            .I3(n40_adj_4979), .O(n3263));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_36_i1529_3_lut_3_lut (.I0(n2288), .I1(n7057), .I2(n2271), 
            .I3(GND_net), .O(n2364));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1529_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 unary_minus_18_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_i1528_3_lut_3_lut (.I0(n2288), .I1(n7056), .I2(n2270), 
            .I3(GND_net), .O(n2363));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1528_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 unary_minus_18_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4332));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_i1524_3_lut_3_lut (.I0(n2288), .I1(n7052), .I2(n2266), 
            .I3(GND_net), .O(n2359));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1524_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1539_3_lut_3_lut (.I0(n2288), .I1(n7067), .I2(n385), 
            .I3(GND_net), .O(n2374));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1539_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_LessThan_1137_i28_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1763), 
            .I3(GND_net), .O(n28_adj_4654));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1137_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(35[10] 38[2])
    SB_LUT4 i22_3_lut_adj_1799 (.I0(bit_ctr[28]), .I1(n42945), .I2(n4754), 
            .I3(GND_net), .O(n35931));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1799.LUT_INIT = 16'hacac;
    coms setpoint_23__I_0 (.rx_data({rx_data}), .PWMLimit({PWMLimit}), .clk32MHz(clk32MHz), 
         .GND_net(GND_net), .n19434(n19434), .setpoint({setpoint}), .n19435(n19435), 
         .n19436(n19436), .n19437(n19437), .n19438(n19438), .n19439(n19439), 
         .n19440(n19440), .n19427(n19427), .n19428(n19428), .n19429(n19429), 
         .n19430(n19430), .n19431(n19431), .control_mode({control_mode}), 
         .VCC_net(VCC_net), .n19448(n19448), .n19449(n19449), .n19446(n19446), 
         .n19447(n19447), .n19444(n19444), .n19445(n19445), .n19441(n19441), 
         .n19442(n19442), .n19443(n19443), .n19432(n19432), .n19433(n19433), 
         .n46050(n46050), .n19145(n19145), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .n19144(n19144), .n19143(n19143), .n19142(n19142), .n19141(n19141), 
         .n19140(n19140), .n19139(n19139), .n19138(n19138), .n19137(n19137), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .n19136(n19136), 
         .n19135(n19135), .n19134(n19134), .n19133(n19133), .n19132(n19132), 
         .n19131(n19131), .n19130(n19130), .n19129(n19129), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .n19128(n19128), .n19127(n19127), .n19126(n19126), .n17199(n17199), 
         .\data_out_frame[5] ({\data_out_frame[5] }), .\data_out_frame[7] ({\data_out_frame[7] }), 
         .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), 
         .n63(n63_adj_4439), .n17268(n17268), .n2857(n2857), .n38098(n38098), 
         .n17200(n17200), .n17202(n17202), .n19125(n19125), .n19124(n19124), 
         .n19123(n19123), .n19122(n19122), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .n19121(n19121), 
         .\data_out_frame[17] ({\data_out_frame[17] }), .n19120(n19120), 
         .n19119(n19119), .n19118(n19118), .n19117(n19117), .n19116(n19116), 
         .n19115(n19115), .n19114(n19114), .n19113(n19113), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .n4661(n4661), .n19112(n19112), .n19111(n19111), .n19110(n19110), 
         .n4659(n4659), .\data_out_frame[12] ({\data_out_frame[12] }), .n19109(n19109), 
         .n19108(n19108), .n19107(n19107), .n19106(n19106), .n19105(n19105), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .n19104(n19104), 
         .n18435(n18435), .n6119(n6119), .ID0(ID0), .n19103(n19103), 
         .n19102(n19102), .rx_data_ready(rx_data_ready), .ID2(ID2), .\data_out_frame[14] ({\data_out_frame[14] }), 
         .n19101(n19101), .n19272(n19272), .\data_in_frame[15] ({\data_in_frame[15] }), 
         .n19271(n19271), .n19270(n19270), .n19100(n19100), .n19099(n19099), 
         .n19098(n19098), .n19097(n19097), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .\data_out_frame[6] ({\data_out_frame[6] }), .n19096(n19096), .n19095(n19095), 
         .\data_out_frame[4][0] (\data_out_frame[4] [0]), .n19094(n19094), 
         .\data_out_frame[4][2] (\data_out_frame[4] [2]), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .\data_out_frame[9] ({\data_out_frame[9] }), .n19093(n19093), .n19092(n19092), 
         .n19091(n19091), .n19090(n19090), .n19089(n19089), .n19088(n19088), 
         .n19087(n19087), .n19086(n19086), .n19085(n19085), .n19084(n19084), 
         .n19083(n19083), .n19082(n19082), .n19081(n19081), .n19080(n19080), 
         .n19079(n19079), .n19078(n19078), .n19077(n19077), .n19076(n19076), 
         .n19075(n19075), .n19074(n19074), .n19073(n19073), .n19072(n19072), 
         .n19071(n19071), .n19070(n19070), .n19069(n19069), .n19068(n19068), 
         .n19067(n19067), .n19066(n19066), .n19065(n19065), .n19269(n19269), 
         .n19064(n19064), .n19268(n19268), .n19063(n19063), .n19062(n19062), 
         .n19061(n19061), .n19060(n19060), .n19059(n19059), .n19058(n19058), 
         .n19057(n19057), .n19056(n19056), .n19055(n19055), .n19054(n19054), 
         .n19053(n19053), .n19052(n19052), .n19051(n19051), .n19050(n19050), 
         .n19049(n19049), .n19048(n19048), .n19047(n19047), .n19046(n19046), 
         .n19045(n19045), .n19044(n19044), .n19043(n19043), .n19267(n19267), 
         .n19042(n19042), .n19041(n19041), .n19040(n19040), .n19039(n19039), 
         .n19038(n19038), .n19266(n19266), .n19037(n19037), .n19036(n19036), 
         .n19035(n19035), .n19034(n19034), .n19033(n19033), .n19032(n19032), 
         .n19265(n19265), .n19031(n19031), .n19030(n19030), .n19029(n19029), 
         .n19028(n19028), .n19027(n19027), .ID1(ID1), .n14536(n14536), 
         .n4660(n4660), .n19026(n19026), .n19025(n19025), .n19024(n19024), 
         .n19023(n19023), .n19022(n19022), .n4673(n4673), .n19021(n19021), 
         .n19020(n19020), .n4672(n4672), .n4671(n4671), .n4670(n4670), 
         .n4669(n4669), .n4668(n4668), .n19019(n19019), .n19018(n19018), 
         .n19017(n19017), .n19014(n19014), .n19013(n19013), .\data_out_frame[0][4] (\data_out_frame[0] [4]), 
         .n19012(n19012), .\data_out_frame[0][3] (\data_out_frame[0] [3]), 
         .n19011(n19011), .\data_in[3] ({\data_in[3] }), .n19010(n19010), 
         .n19009(n19009), .n19008(n19008), .n19007(n19007), .n19006(n19006), 
         .n19005(n19005), .n19004(n19004), .n19003(n19003), .\data_in[2] ({\data_in[2] }), 
         .n19002(n19002), .n19001(n19001), .n19000(n19000), .n18999(n18999), 
         .n18998(n18998), .n18997(n18997), .n18996(n18996), .n18995(n18995), 
         .\data_in[1] ({\data_in[1] }), .n18994(n18994), .n18993(n18993), 
         .n18992(n18992), .n18991(n18991), .n18990(n18990), .n18989(n18989), 
         .n18988(n18988), .n18987(n18987), .\data_in[0] ({\data_in[0] }), 
         .n18986(n18986), .n18985(n18985), .n18984(n18984), .n18983(n18983), 
         .n18982(n18982), .n18981(n18981), .\Ki[7] (Ki[7]), .\Ki[6] (Ki[6]), 
         .\Ki[5] (Ki[5]), .\Ki[4] (Ki[4]), .\Ki[3] (Ki[3]), .\Ki[2] (Ki[2]), 
         .\Ki[1] (Ki[1]), .\Kp[7] (Kp[7]), .\Kp[6] (Kp[6]), .\Kp[5] (Kp[5]), 
         .\Kp[4] (Kp[4]), .\Kp[3] (Kp[3]), .\Kp[2] (Kp[2]), .\Kp[1] (Kp[1]), 
         .gearBoxRatio({gearBoxRatio}), .IntegralLimit({IntegralLimit}), 
         .\Kp[0] (Kp[0]), .\Ki[0] (Ki[0]), .\data_in_frame[7] ({\data_in_frame[7] }), 
         .n37368(n37368), .n17264(n17264), .n37348(n37348), .n18829(n18829), 
         .n19208(n19208), .n3761(n3761), .n740(n740), .n19207(n19207), 
         .n19206(n19206), .n19205(n19205), .n19204(n19204), .n2664(n2664), 
         .n36597(n36597), .n19203(n19203), .n18798(n18798), .LED_c(LED_c), 
         .n20639(n20639), .n5(n5_adj_4440), .n46559(n46559), .n5_adj_3(n5_adj_4989), 
         .n19202(n19202), .n19201(n19201), .n37376(n37376), .n40(n40_adj_4988), 
         .n4666(n4666), .n4665(n4665), .n4676(n4676), .n4675(n4675), 
         .n4674(n4674), .n4678(n4678), .n4677(n4677), .n4680(n4680), 
         .n4679(n4679), .n4682(n4682), .n4681(n4681), .n39863(n39863), 
         .n4667(n4667), .n4664(n4664), .n4663(n4663), .n4662(n4662), 
         .n18758(n18758), .n18755(n18755), .n18752(n18752), .n18749(n18749), 
         .n19426(n19426), .r_SM_Main({r_SM_Main_adj_5046}), .n18746(n18746), 
         .n18767(n18767), .n18764(n18764), .n18761(n18761), .n18744(n18744), 
         .n18747(n18747), .\r_SM_Main_2__N_3320[1] (r_SM_Main_2__N_3320[1]), 
         .n18750(n18750), .n18753(n18753), .n18756(n18756), .n18759(n18759), 
         .n18762(n18762), .n18765(n18765), .n18896(n18896), .n18898(n18898), 
         .n18816(n18816), .n18815(n18815), .tx_active(tx_active), .n18814(n18814), 
         .tx_o(tx_o), .n45935(n45935), .tx_enable(tx_enable), .n18402(n18402), 
         .n12501(n12501), .n18897(n18897), .n36985(n36985), .\r_Clock_Count[2] (r_Clock_Count[2]), 
         .n36987(n36987), .\r_Clock_Count[3] (r_Clock_Count[3]), .n36989(n36989), 
         .\r_Clock_Count[4] (r_Clock_Count[4]), .n36919(n36919), .\r_Clock_Count[5] (r_Clock_Count[5]), 
         .n36743(n36743), .\r_Clock_Count[6] (r_Clock_Count[6]), .n36695(n36695), 
         .\r_Clock_Count[7] (r_Clock_Count[7]), .n36983(n36983), .\r_Clock_Count[1] (r_Clock_Count[1]), 
         .n18780(n18780), .r_Bit_Index({r_Bit_Index}), .n18777(n18777), 
         .n19419(n19419), .n27445(n27445), .\r_SM_Main[1]_adj_4 (r_SM_Main[1]), 
         .n95(n95), .n16(n16_adj_4990), .\r_SM_Main[2]_adj_5 (r_SM_Main[2]), 
         .r_Rx_Data(r_Rx_Data), .PIN_13_N_105(PIN_13_N_105), .n37215(n37215), 
         .n37220(n37220), .n37217(n37217), .n37216(n37216), .n37218(n37218), 
         .n37219(n37219), .n37214(n37214), .n18943(n18943), .n18806(n18806), 
         .n18793(n18793), .n18786(n18786), .n18785(n18785), .n18784(n18784), 
         .n18783(n18783), .n18782(n18782), .n18781(n18781), .n42920(n42920), 
         .n20874(n20874), .n42919(n42919), .n17255(n17255), .n4(n4), 
         .n26349(n26349), .n4_adj_6(n4_adj_4365), .n4_adj_7(n4_adj_4412), 
         .n17250(n17250), .n4926(n4926), .n18467(n18467), .n20896(n20896), 
         .n18602(n18602)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(195[8] 216[4])
    SB_LUT4 mux_61_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[21]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i22_3_lut (.I0(encoder0_position[21]), .I1(motor_state_23__N_106[21]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1531_3_lut_3_lut (.I0(n2288), .I1(n7059), .I2(n2273), 
            .I3(GND_net), .O(n2366));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1531_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1534_3_lut_3_lut (.I0(n2288), .I1(n7062), .I2(n2276), 
            .I3(GND_net), .O(n2369));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1534_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13749_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n26349), 
            .I3(n17250), .O(n18781));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13749_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i35898_2_lut_4_lut (.I0(n1758), .I1(n92), .I2(n1762), .I3(n96), 
            .O(n43022));
    defparam i35898_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i14402_3_lut (.I0(setpoint[8]), .I1(n4667), .I2(n39863), .I3(GND_net), 
            .O(n19434));   // verilog/coms.v(126[12] 289[6])
    defparam i14402_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_LessThan_1137_i30_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1758), 
            .I3(GND_net), .O(n30_adj_4656));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1137_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i13750_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n26349), 
            .I3(n17255), .O(n18782));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13750_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 div_36_i1535_3_lut_3_lut (.I0(n2288), .I1(n7063), .I2(n2277), 
            .I3(GND_net), .O(n2370));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1535_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13751_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_4365), 
            .I3(n17250), .O(n18783));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13751_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13752_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_4365), 
            .I3(n17255), .O(n18784));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13752_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13753_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_4412), 
            .I3(n17250), .O(n18785));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13753_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13754_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_4412), 
            .I3(n17255), .O(n18786));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13754_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_36_i1533_3_lut_3_lut (.I0(n2288), .I1(n7061), .I2(n2275), 
            .I3(GND_net), .O(n2368));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1533_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1527_3_lut_3_lut (.I0(n2288), .I1(n7055), .I2(n2269), 
            .I3(GND_net), .O(n2362));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1527_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13761_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4), .I3(n17250), 
            .O(n18793));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13761_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_36_LessThan_1210_i26_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1872), 
            .I3(GND_net), .O(n26_adj_4666));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1210_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i36602_2_lut_4_lut (.I0(n1867), .I1(n92), .I2(n1871), .I3(n96), 
            .O(n43727));
    defparam i36602_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_36_LessThan_1210_i28_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1867), 
            .I3(GND_net), .O(n28_adj_4668));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1210_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i13766_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n18798));   // verilog/coms.v(126[12] 289[6])
    defparam i13766_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31034_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(GND_net), .I3(GND_net), .O(n38094));
    defparam i31034_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i35878_2_lut_4_lut (.I0(n1869), .I1(n94), .I2(n1870), .I3(n95_adj_4360), 
            .O(n43002));
    defparam i35878_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i36495_2_lut (.I0(start), .I1(n27453), .I2(GND_net), .I3(GND_net), 
            .O(n42970));   // verilog/neopixel.v(35[12] 117[6])
    defparam i36495_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i31_4_lut (.I0(n42970), .I1(n42968), .I2(state[1]), .I3(\neo_pixel_transmitter.done ), 
            .O(n35977));   // verilog/neopixel.v(35[12] 117[6])
    defparam i31_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 unary_minus_18_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4331));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_61_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[22]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_60_i23_3_lut (.I0(encoder0_position[22]), .I1(motor_state_23__N_106[22]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1210_i30_3_lut_3_lut (.I0(n95_adj_4360), .I1(n94), 
            .I2(n1869), .I3(GND_net), .O(n30_adj_4670));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1210_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 unary_minus_18_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14171_3_lut (.I0(\data_in_frame[7] [2]), .I1(rx_data[2]), .I2(n37368), 
            .I3(GND_net), .O(n19203));   // verilog/coms.v(126[12] 289[6])
    defparam i14171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2069_rep_56_3_lut (.I0(n3044), .I1(n3111), .I2(n3065), 
            .I3(GND_net), .O(n3143));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2069_rep_56_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1281_i24_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1978), 
            .I3(GND_net), .O(n24_adj_4684));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1281_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i36551_2_lut_4_lut (.I0(n1973), .I1(n92), .I2(n1977), .I3(n96), 
            .O(n43676));
    defparam i36551_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 rem_4_i2072_3_lut (.I0(n3047), .I1(n3114), .I2(n3065), .I3(GND_net), 
            .O(n3146));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2077_3_lut (.I0(n3052), .I1(n3119), .I2(n3065), .I3(GND_net), 
            .O(n3151));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2076_3_lut (.I0(n3051), .I1(n3118), .I2(n3065), .I3(GND_net), 
            .O(n3150));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2058_3_lut (.I0(n3033), .I1(n3100), .I2(n3065), .I3(GND_net), 
            .O(n3132));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2074_3_lut (.I0(n3049), .I1(n3116), .I2(n3065), .I3(GND_net), 
            .O(n3148));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2078_3_lut (.I0(n3053), .I1(n3120), .I2(n3065), .I3(GND_net), 
            .O(n3152));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2075_3_lut (.I0(n3050), .I1(n3117), .I2(n3065), .I3(GND_net), 
            .O(n3149));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2070_3_lut (.I0(n3045), .I1(n3112), .I2(n3065), .I3(GND_net), 
            .O(n3144));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2066_3_lut (.I0(n3041), .I1(n3108), .I2(n3065), .I3(GND_net), 
            .O(n3140));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2065_3_lut (.I0(n3040), .I1(n3107), .I2(n3065), .I3(GND_net), 
            .O(n3139));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2064_3_lut (.I0(n3039), .I1(n3106), .I2(n3065), .I3(GND_net), 
            .O(n3138));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2062_3_lut (.I0(n3037), .I1(n3104), .I2(n3065), .I3(GND_net), 
            .O(n3136));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2063_3_lut (.I0(n3038), .I1(n3105), .I2(n3065), .I3(GND_net), 
            .O(n3137));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2061_3_lut (.I0(n3036), .I1(n3103), .I2(n3065), .I3(GND_net), 
            .O(n3135));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2060_3_lut (.I0(n3035), .I1(n3102), .I2(n3065), .I3(GND_net), 
            .O(n3134));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2059_3_lut (.I0(n3034), .I1(n3101), .I2(n3065), .I3(GND_net), 
            .O(n3133));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2073_3_lut (.I0(n3048), .I1(n3115), .I2(n3065), .I3(GND_net), 
            .O(n3147));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2079_3_lut (.I0(n3054), .I1(n3121), .I2(n3065), .I3(GND_net), 
            .O(n3153));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2071_3_lut (.I0(n3046), .I1(n3113), .I2(n3065), .I3(GND_net), 
            .O(n3145));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1281_i26_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1973), 
            .I3(GND_net), .O(n26_adj_4686));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1281_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 rem_4_i2068_3_lut (.I0(n3043), .I1(n3110), .I2(n3065), .I3(GND_net), 
            .O(n3142));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2081_3_lut (.I0(n3056), .I1(n3123), .I2(n3065), .I3(GND_net), 
            .O(n3155));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2067_3_lut (.I0(n3042), .I1(n3109), .I2(n3065), .I3(GND_net), 
            .O(n3141));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2080_3_lut (.I0(n3055), .I1(n3122), .I2(n3065), .I3(GND_net), 
            .O(n3154));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i5_3_lut (.I0(communication_counter[4]), .I1(n29_adj_4380), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3158));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2083_3_lut (.I0(n3058), .I1(n3125), .I2(n3065), .I3(GND_net), 
            .O(n3157));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36555_2_lut_4_lut (.I0(n1975), .I1(n94), .I2(n1976), .I3(n95_adj_4360), 
            .O(n43680));
    defparam i36555_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 rem_4_i2082_3_lut (.I0(n3057), .I1(n3124), .I2(n3065), .I3(GND_net), 
            .O(n3156));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1800 (.I0(n3156), .I1(n3157), .I2(n3158), .I3(GND_net), 
            .O(n38353));
    defparam i1_3_lut_adj_1800.LUT_INIT = 16'hfefe;
    SB_LUT4 div_36_LessThan_1281_i28_3_lut_3_lut (.I0(n95_adj_4360), .I1(n94), 
            .I2(n1975), .I3(GND_net), .O(n28_adj_4688));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1281_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i6_4_lut_adj_1801 (.I0(n3154), .I1(n3141), .I2(n38353), .I3(n3155), 
            .O(n30_adj_4997));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i6_4_lut_adj_1801.LUT_INIT = 16'heccc;
    SB_LUT4 i16_4_lut_adj_1802 (.I0(n3142), .I1(n3145), .I2(n3153), .I3(n3147), 
            .O(n40_adj_4995));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i16_4_lut_adj_1802.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(n3133), .I1(n3134), .I2(GND_net), .I3(GND_net), 
            .O(n26_adj_4998));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i14_4_lut_adj_1803 (.I0(n3135), .I1(n3137), .I2(n3136), .I3(n3138), 
            .O(n38_adj_4996));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i14_4_lut_adj_1803.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1804 (.I0(n3139), .I1(n40_adj_4995), .I2(n30_adj_4997), 
            .I3(n3140), .O(n44_adj_4991));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i20_4_lut_adj_1804.LUT_INIT = 16'hfffe;
    SB_LUT4 i14369_3_lut (.I0(encoder1_position[23]), .I1(n2816), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19401));   // quad.v(35[10] 41[6])
    defparam i14369_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18_4_lut_adj_1805 (.I0(n3144), .I1(n3149), .I2(n3152), .I3(n3148), 
            .O(n42_adj_4993));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i18_4_lut_adj_1805.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1806 (.I0(n3132), .I1(n38_adj_4996), .I2(n26_adj_4998), 
            .I3(n3131), .O(n43_adj_4992));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i19_4_lut_adj_1806.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1807 (.I0(n3150), .I1(n3151), .I2(n3146), .I3(n3143), 
            .O(n41_adj_4994));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i17_4_lut_adj_1807.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(n41_adj_4994), .I1(n43_adj_4992), .I2(n42_adj_4993), 
            .I3(n44_adj_4991), .O(n3164));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14368_3_lut (.I0(encoder1_position[22]), .I1(n2817), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19400));   // quad.v(35[10] 41[6])
    defparam i14368_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14367_3_lut (.I0(encoder1_position[21]), .I1(n2818), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19399));   // quad.v(35[10] 41[6])
    defparam i14367_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1350_i22_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2081), 
            .I3(GND_net), .O(n22_adj_4702));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1350_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i36488_2_lut_4_lut (.I0(n2076), .I1(n92), .I2(n2080), .I3(n96), 
            .O(n43613));
    defparam i36488_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i4_4_lut_adj_1808 (.I0(control_mode[3]), .I1(control_mode[7]), 
            .I2(control_mode[4]), .I3(control_mode[5]), .O(n10_adj_4433));   // verilog/TinyFPGA_B.v(221[5:22])
    defparam i4_4_lut_adj_1808.LUT_INIT = 16'hfffe;
    SB_LUT4 i14366_3_lut (.I0(encoder1_position[20]), .I1(n2819), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19398));   // quad.v(35[10] 41[6])
    defparam i14366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_adj_1809 (.I0(control_mode[6]), .I1(n10_adj_4433), 
            .I2(control_mode[2]), .I3(GND_net), .O(n17189));   // verilog/TinyFPGA_B.v(221[5:22])
    defparam i5_3_lut_adj_1809.LUT_INIT = 16'hfefe;
    SB_LUT4 div_36_LessThan_1350_i24_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2076), 
            .I3(GND_net), .O(n24_adj_4704));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1350_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i2_3_lut (.I0(control_mode[0]), .I1(control_mode[1]), .I2(n17189), 
            .I3(GND_net), .O(n15_adj_4359));   // verilog/TinyFPGA_B.v(222[5:22])
    defparam i2_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i14365_3_lut (.I0(encoder1_position[19]), .I1(n2820), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19397));   // quad.v(35[10] 41[6])
    defparam i14365_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_61_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15_adj_4359), .I3(n15_adj_4361), .O(motor_state_23__N_106[23]));   // verilog/TinyFPGA_B.v(222[5] 225[10])
    defparam mux_61_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14364_3_lut (.I0(encoder1_position[18]), .I1(n2821), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19396));   // quad.v(35[10] 41[6])
    defparam i14364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_60_i24_3_lut (.I0(encoder0_position[23]), .I1(motor_state_23__N_106[23]), 
            .I2(n15_adj_4368), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(221[5] 225[10])
    defparam mux_60_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36500_2_lut_4_lut (.I0(n2078), .I1(n94), .I2(n2079), .I3(n95_adj_4360), 
            .O(n43625));
    defparam i36500_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_36_LessThan_1350_i26_3_lut_3_lut (.I0(n95_adj_4360), .I1(n94), 
            .I2(n2078), .I3(GND_net), .O(n26_adj_4706));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1350_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i14363_3_lut (.I0(encoder1_position[17]), .I1(n2822), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n19395));   // quad.v(35[10] 41[6])
    defparam i14363_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13770_3_lut (.I0(encoder0_position[0]), .I1(n2889), .I2(count_enable), 
            .I3(GND_net), .O(n18802));   // quad.v(35[10] 41[6])
    defparam i13770_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33740_4_lut (.I0(n17202), .I1(n17268), .I2(n740), .I3(n2857), 
            .O(n40805));
    defparam i33740_4_lut.LUT_INIT = 16'hfac8;
    SB_LUT4 i13745_4_lut (.I0(n18602), .I1(r_Bit_Index[2]), .I2(n4926), 
            .I3(n18467), .O(n18777));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13745_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i1_4_lut_adj_1810 (.I0(n38098), .I1(n40_adj_4988), .I2(n40805), 
            .I3(n37376), .O(n41_adj_4987));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1810.LUT_INIT = 16'hcc4c;
    SB_LUT4 i1_4_lut_adj_1811 (.I0(n17199), .I1(n41_adj_4987), .I2(\FRAME_MATCHER.state [3]), 
            .I3(\FRAME_MATCHER.state [0]), .O(n36597));   // verilog/coms.v(126[12] 289[6])
    defparam i1_4_lut_adj_1811.LUT_INIT = 16'hccdc;
    SB_LUT4 i13772_3_lut (.I0(encoder1_position[0]), .I1(n2839), .I2(count_enable_adj_4374), 
            .I3(GND_net), .O(n18804));   // quad.v(35[10] 41[6])
    defparam i13772_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13773_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n39036), 
            .I3(GND_net), .O(n18805));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13774_4_lut (.I0(r_SM_Main[2]), .I1(n20874), .I2(n20896), 
            .I3(r_SM_Main[1]), .O(n18806));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13774_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 unary_minus_18_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4330));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_4_inv_0_i1_1_lut (.I0(gearBoxRatio[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4544));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13778_3_lut (.I0(\half_duty[0] [0]), .I1(half_duty_new[0]), 
            .I2(n1111), .I3(GND_net), .O(n18810));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13778_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14172_3_lut (.I0(\data_in_frame[7] [3]), .I1(rx_data[3]), .I2(n37368), 
            .I3(GND_net), .O(n19204));   // verilog/coms.v(126[12] 289[6])
    defparam i14172_3_lut.LUT_INIT = 16'hacac;
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.n19372(n19372), .encoder0_position({encoder0_position}), 
            .clk32MHz(clk32MHz), .n19373(n19373), .n19374(n19374), .n19375(n19375), 
            .n19376(n19376), .n19377(n19377), .n19368(n19368), .n19369(n19369), 
            .n19370(n19370), .n19371(n19371), .n19366(n19366), .n19367(n19367), 
            .n19364(n19364), .n19365(n19365), .n19362(n19362), .n19363(n19363), 
            .n19360(n19360), .n19361(n19361), .n19358(n19358), .n19359(n19359), 
            .n19355(n19355), .n19356(n19356), .n19357(n19357), .data_o({quadA_debounced, 
            quadB_debounced}), .n2865({n2866, n2867, n2868, n2869, 
            n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, 
            n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, 
            n2886, n2887, n2888, n2889}), .GND_net(GND_net), .n18802(n18802), 
            .count_enable(count_enable), .n19406(n19406), .reg_B({reg_B}), 
            .PIN_2_c_0(PIN_2_c_0), .n18805(n18805), .PIN_1_c_1(PIN_1_c_1), 
            .n39036(n39036)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(247[15] 252[4])
    SB_LUT4 i14173_3_lut (.I0(\data_in_frame[7] [4]), .I1(rx_data[4]), .I2(n37368), 
            .I3(GND_net), .O(n19205));   // verilog/coms.v(126[12] 289[6])
    defparam i14173_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14174_3_lut (.I0(\data_in_frame[7] [5]), .I1(rx_data[5]), .I2(n37368), 
            .I3(GND_net), .O(n19206));   // verilog/coms.v(126[12] 289[6])
    defparam i14174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14175_3_lut (.I0(\data_in_frame[7] [6]), .I1(rx_data[6]), .I2(n37368), 
            .I3(GND_net), .O(n19207));   // verilog/coms.v(126[12] 289[6])
    defparam i14175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i19654_3_lut (.I0(r_SM_Main_adj_5046[0]), .I1(n45935), .I2(r_SM_Main_adj_5046[1]), 
            .I3(GND_net), .O(n24672));   // verilog/uart_tx.v(31[16:25])
    defparam i19654_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i19655_3_lut (.I0(tx_o), .I1(n24672), .I2(r_SM_Main_adj_5046[2]), 
            .I3(GND_net), .O(n18814));
    defparam i19655_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_unary_minus_4_inv_0_i2_1_lut (.I0(gearBoxRatio[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_4543));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_4_inv_0_i3_1_lut (.I0(gearBoxRatio[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4542));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_4_inv_0_i4_1_lut (.I0(gearBoxRatio[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_4541));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13748_4_lut (.I0(n18602), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(n18467), .O(n18780));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13748_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i22_3_lut_adj_1812 (.I0(bit_ctr[31]), .I1(n42951), .I2(n4754), 
            .I3(GND_net), .O(n35943));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1812.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1813 (.I0(bit_ctr[30]), .I1(n42950), .I2(n4754), 
            .I3(GND_net), .O(n35941));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1813.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1814 (.I0(bit_ctr[19]), .I1(n42949), .I2(n4754), 
            .I3(GND_net), .O(n35939));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1814.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1815 (.I0(bit_ctr[18]), .I1(n42948), .I2(n4754), 
            .I3(GND_net), .O(n35937));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1815.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1816 (.I0(bit_ctr[17]), .I1(n42947), .I2(n4754), 
            .I3(GND_net), .O(n35935));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1816.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1817 (.I0(bit_ctr[29]), .I1(n42946), .I2(n4754), 
            .I3(GND_net), .O(n35933));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1817.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_unary_minus_4_inv_0_i5_1_lut (.I0(gearBoxRatio[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4540));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13729_2_lut (.I0(n18897), .I1(n18759), .I2(GND_net), .I3(GND_net), 
            .O(n18761));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13729_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13732_2_lut (.I0(n18897), .I1(n18762), .I2(GND_net), .I3(GND_net), 
            .O(n18764));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13732_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_18_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_4_inv_0_i6_1_lut (.I0(gearBoxRatio[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4539));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13735_2_lut (.I0(n18897), .I1(n18765), .I2(GND_net), .I3(GND_net), 
            .O(n18767));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13735_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_36_unary_minus_4_inv_0_i7_1_lut (.I0(gearBoxRatio[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4538));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_4_inv_0_i8_1_lut (.I0(gearBoxRatio[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4537));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_4_inv_0_i9_1_lut (.I0(gearBoxRatio[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4536));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_4_inv_0_i10_1_lut (.I0(gearBoxRatio[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4535));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19659_3_lut (.I0(n18402), .I1(r_SM_Main_adj_5046[1]), .I2(tx_active), 
            .I3(GND_net), .O(n18815));   // verilog/uart_tx.v(31[16:25])
    defparam i19659_3_lut.LUT_INIT = 16'h7272;
    SB_LUT4 div_36_unary_minus_4_inv_0_i11_1_lut (.I0(gearBoxRatio[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4534));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13784_4_lut (.I0(r_SM_Main_adj_5046[2]), .I1(n12501), .I2(r_SM_Main_2__N_3320[1]), 
            .I3(r_SM_Main_adj_5046[0]), .O(n18816));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13784_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i1_3_lut_adj_1818 (.I0(n37214), .I1(r_Clock_Count[1]), .I2(n16_adj_4990), 
            .I3(GND_net), .O(n36983));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_1818.LUT_INIT = 16'heaea;
    SB_LUT4 i13714_2_lut (.I0(n18897), .I1(n18744), .I2(GND_net), .I3(GND_net), 
            .O(n18746));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13714_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22_3_lut_adj_1819 (.I0(bit_ctr[2]), .I1(n42953), .I2(n4754), 
            .I3(GND_net), .O(n35949));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1819.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1820 (.I0(bit_ctr[1]), .I1(n42952), .I2(n4754), 
            .I3(GND_net), .O(n35947));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1820.LUT_INIT = 16'hacac;
    SB_LUT4 i1_3_lut_adj_1821 (.I0(n37215), .I1(r_Clock_Count[7]), .I2(n16_adj_4990), 
            .I3(GND_net), .O(n36695));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_adj_1821.LUT_INIT = 16'heaea;
    SB_LUT4 i22_3_lut_adj_1822 (.I0(bit_ctr[4]), .I1(n42955), .I2(n4754), 
            .I3(GND_net), .O(n35953));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1822.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1823 (.I0(bit_ctr[3]), .I1(n42954), .I2(n4754), 
            .I3(GND_net), .O(n35951));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1823.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2003_3_lut (.I0(n2946), .I1(n3013), .I2(n2966), .I3(GND_net), 
            .O(n3045));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2009_3_lut (.I0(n2952), .I1(n3019), .I2(n2966), .I3(GND_net), 
            .O(n3051));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2005_3_lut (.I0(n2948), .I1(n3015), .I2(n2966), .I3(GND_net), 
            .O(n3047));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1824 (.I0(bit_ctr[6]), .I1(n42957), .I2(n4754), 
            .I3(GND_net), .O(n35957));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1824.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1825 (.I0(bit_ctr[5]), .I1(n42956), .I2(n4754), 
            .I3(GND_net), .O(n35955));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1825.LUT_INIT = 16'hacac;
    SB_LUT4 i22_3_lut_adj_1826 (.I0(bit_ctr[8]), .I1(n42959), .I2(n4754), 
            .I3(GND_net), .O(n35961));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1826.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2002_3_lut (.I0(n2945), .I1(n3012), .I2(n2966), .I3(GND_net), 
            .O(n3044));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1991_3_lut (.I0(n2934), .I1(n3001), .I2(n2966), .I3(GND_net), 
            .O(n3033));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2007_3_lut (.I0(n2950), .I1(n3017), .I2(n2966), .I3(GND_net), 
            .O(n3049));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2006_3_lut (.I0(n2949), .I1(n3016), .I2(n2966), .I3(GND_net), 
            .O(n3048));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2011_3_lut (.I0(n2954), .I1(n3021), .I2(n2966), .I3(GND_net), 
            .O(n3053));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1827 (.I0(bit_ctr[7]), .I1(n42958), .I2(n4754), 
            .I3(GND_net), .O(n35959));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1827.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2008_3_lut (.I0(n2951), .I1(n3018), .I2(n2966), .I3(GND_net), 
            .O(n3050));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2004_3_lut (.I0(n2947), .I1(n3014), .I2(n2966), .I3(GND_net), 
            .O(n3046));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2004_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2010_3_lut (.I0(n2953), .I1(n3020), .I2(n2966), .I3(GND_net), 
            .O(n3052));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2001_3_lut (.I0(n2944), .I1(n3011), .I2(n2966), .I3(GND_net), 
            .O(n3043));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1995_3_lut (.I0(n2938), .I1(n3005), .I2(n2966), .I3(GND_net), 
            .O(n3037));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1993_3_lut (.I0(n2936), .I1(n3003), .I2(n2966), .I3(GND_net), 
            .O(n3035));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1994_3_lut (.I0(n2937), .I1(n3004), .I2(n2966), .I3(GND_net), 
            .O(n3036));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1992_3_lut (.I0(n2935), .I1(n3002), .I2(n2966), .I3(GND_net), 
            .O(n3034));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1999_3_lut (.I0(n2942), .I1(n3009), .I2(n2966), .I3(GND_net), 
            .O(n3041));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1997_3_lut (.I0(n2940), .I1(n3007), .I2(n2966), .I3(GND_net), 
            .O(n3039));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1828 (.I0(bit_ctr[10]), .I1(n42961), .I2(n4754), 
            .I3(GND_net), .O(n35965));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1828.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_i1598_3_lut_3_lut (.I0(n2381), .I1(n7085), .I2(n2372), 
            .I3(GND_net), .O(n2462));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1598_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1583_3_lut_3_lut (.I0(n2381), .I1(n7070), .I2(n2357), 
            .I3(GND_net), .O(n2447));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1583_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1998_3_lut (.I0(n2941), .I1(n3008), .I2(n2966), .I3(GND_net), 
            .O(n3040));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1996_3_lut (.I0(n2939), .I1(n3006), .I2(n2966), .I3(GND_net), 
            .O(n3038));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i1996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2013_3_lut (.I0(n2956), .I1(n3023), .I2(n2966), .I3(GND_net), 
            .O(n3055));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2012_3_lut (.I0(n2955), .I1(n3022), .I2(n2966), .I3(GND_net), 
            .O(n3054));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2000_3_lut (.I0(n2943), .I1(n3010), .I2(n2966), .I3(GND_net), 
            .O(n3042));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i6_3_lut (.I0(communication_counter[5]), .I1(n28), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3058));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22_3_lut_adj_1829 (.I0(bit_ctr[9]), .I1(n42960), .I2(n4754), 
            .I3(GND_net), .O(n35963));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1829.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2015_3_lut (.I0(n2958), .I1(n3025), .I2(n2966), .I3(GND_net), 
            .O(n3057));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2014_3_lut (.I0(n2957), .I1(n3024), .I2(n2966), .I3(GND_net), 
            .O(n3056));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam rem_4_i2014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1830 (.I0(n3056), .I1(n3057), .I2(n3058), .I3(GND_net), 
            .O(n38405));
    defparam i1_3_lut_adj_1830.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1831 (.I0(n3042), .I1(n3054), .I2(n38405), .I3(n3055), 
            .O(n29));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i6_4_lut_adj_1831.LUT_INIT = 16'heaaa;
    SB_LUT4 i14_4_lut_adj_1832 (.I0(n3038), .I1(n3040), .I2(n3039), .I3(n3041), 
            .O(n37_adj_4353));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i14_4_lut_adj_1832.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1833 (.I0(n3034), .I1(n3036), .I2(n3035), .I3(n3037), 
            .O(n36));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i13_4_lut_adj_1833.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1834 (.I0(n37_adj_4353), .I1(n29), .I2(n3043), 
            .I3(n3052), .O(n42));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i19_4_lut_adj_1834.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1835 (.I0(n3046), .I1(n3050), .I2(n3053), .I3(n3048), 
            .O(n40_adj_4351));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i17_4_lut_adj_1835.LUT_INIT = 16'hfffe;
    SB_LUT4 div_36_i1584_3_lut_3_lut (.I0(n2381), .I1(n7071), .I2(n2358), 
            .I3(GND_net), .O(n2448));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1584_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1587_3_lut_3_lut (.I0(n2381), .I1(n7074), .I2(n2361), 
            .I3(GND_net), .O(n2451));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1587_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i22_3_lut_adj_1836 (.I0(bit_ctr[12]), .I1(n42963), .I2(n4754), 
            .I3(GND_net), .O(n35969));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1836.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_i1588_3_lut_3_lut (.I0(n2381), .I1(n7075), .I2(n2362), 
            .I3(GND_net), .O(n2452));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1588_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i22_3_lut_adj_1837 (.I0(bit_ctr[11]), .I1(n42962), .I2(n4754), 
            .I3(GND_net), .O(n35967));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1837.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_i1585_3_lut_3_lut (.I0(n2381), .I1(n7072), .I2(n2359), 
            .I3(GND_net), .O(n2449));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1585_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1586_3_lut_3_lut (.I0(n2381), .I1(n7073), .I2(n2360), 
            .I3(GND_net), .O(n2450));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1586_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i18_4_lut_adj_1838 (.I0(n3049), .I1(n36), .I2(n3033), .I3(n3032), 
            .O(n41));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i18_4_lut_adj_1838.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1839 (.I0(n3044), .I1(n3047), .I2(n3051), .I3(n3045), 
            .O(n39_adj_4352));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i16_4_lut_adj_1839.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1840 (.I0(n39_adj_4352), .I1(n41), .I2(n40_adj_4351), 
            .I3(n42), .O(n3065));   // verilog/TinyFPGA_B.v(51[6:33])
    defparam i22_4_lut_adj_1840.LUT_INIT = 16'hfffe;
    SB_LUT4 i14399_3_lut (.I0(setpoint[5]), .I1(n4664), .I2(n39863), .I3(GND_net), 
            .O(n19431));   // verilog/coms.v(126[12] 289[6])
    defparam i14399_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_i1594_3_lut_3_lut (.I0(n2381), .I1(n7081), .I2(n2368), 
            .I3(GND_net), .O(n2458));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1594_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1600_3_lut_3_lut (.I0(n2381), .I1(n7087), .I2(n2374), 
            .I3(GND_net), .O(n2464));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1600_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14398_3_lut (.I0(setpoint[4]), .I1(n4663), .I2(n39863), .I3(GND_net), 
            .O(n19430));   // verilog/coms.v(126[12] 289[6])
    defparam i14398_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14176_3_lut (.I0(\data_in_frame[7] [7]), .I1(rx_data[7]), .I2(n37368), 
            .I3(GND_net), .O(n19208));   // verilog/coms.v(126[12] 289[6])
    defparam i14176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_LessThan_1417_i20_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2181), 
            .I3(GND_net), .O(n20_adj_4720));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i36437_2_lut_4_lut (.I0(n2176), .I1(n92), .I2(n2180), .I3(n96), 
            .O(n43562));
    defparam i36437_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_36_LessThan_1417_i22_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2176), 
            .I3(GND_net), .O(n22_adj_4722));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_36_LessThan_1417_i24_3_lut_3_lut (.I0(n95_adj_4360), .I1(n94), 
            .I2(n2178), .I3(GND_net), .O(n24_adj_4724));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1417_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_36_i1589_3_lut_3_lut (.I0(n2381), .I1(n7076), .I2(n2363), 
            .I3(GND_net), .O(n2453));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1589_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1591_3_lut_3_lut (.I0(n2381), .I1(n7078), .I2(n2365), 
            .I3(GND_net), .O(n2455));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1591_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i36452_2_lut_4_lut (.I0(n2178), .I1(n94), .I2(n2179), .I3(n95_adj_4360), 
            .O(n43577));
    defparam i36452_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_36_LessThan_1482_i18_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2278), 
            .I3(GND_net), .O(n18_adj_4742));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_36_unary_minus_4_inv_0_i12_1_lut (.I0(gearBoxRatio[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4533));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36380_2_lut_4_lut (.I0(n2273), .I1(n92), .I2(n2277), .I3(n96), 
            .O(n43505));
    defparam i36380_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_36_unary_minus_4_inv_0_i13_1_lut (.I0(gearBoxRatio[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4532));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_1482_i20_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2273), 
            .I3(GND_net), .O(n20_adj_4744));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_36_i1590_3_lut_3_lut (.I0(n2381), .I1(n7077), .I2(n2364), 
            .I3(GND_net), .O(n2454));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1590_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_LessThan_1482_i22_3_lut_3_lut (.I0(n95_adj_4360), .I1(n94), 
            .I2(n2275), .I3(GND_net), .O(n22_adj_4746));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1482_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_36_unary_minus_4_inv_0_i14_1_lut (.I0(gearBoxRatio[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_4531));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_4_inv_0_i15_1_lut (.I0(gearBoxRatio[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4530));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_i1601_3_lut_3_lut (.I0(n2381), .I1(n7088), .I2(n386), 
            .I3(GND_net), .O(n2465));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1601_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_unary_minus_4_inv_0_i16_1_lut (.I0(gearBoxRatio[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4529));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4329));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_4_inv_0_i17_1_lut (.I0(gearBoxRatio[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4528));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_i1593_3_lut_3_lut (.I0(n2381), .I1(n7080), .I2(n2367), 
            .I3(GND_net), .O(n2457));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1593_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1592_3_lut_3_lut (.I0(n2381), .I1(n7079), .I2(n2366), 
            .I3(GND_net), .O(n2456));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1592_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i36384_2_lut_4_lut (.I0(n2275), .I1(n94), .I2(n2276), .I3(n95_adj_4360), 
            .O(n43509));
    defparam i36384_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_36_i1599_3_lut_3_lut (.I0(n2381), .I1(n7086), .I2(n2373), 
            .I3(GND_net), .O(n2463));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1599_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1597_3_lut_3_lut (.I0(n2381), .I1(n7084), .I2(n2371), 
            .I3(GND_net), .O(n2461));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1597_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_LessThan_1545_i16_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2372), 
            .I3(GND_net), .O(n16_adj_4760));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_36_i1596_3_lut_3_lut (.I0(n2381), .I1(n7083), .I2(n2370), 
            .I3(GND_net), .O(n2460));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1596_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1595_3_lut_3_lut (.I0(n2381), .I1(n7082), .I2(n2369), 
            .I3(GND_net), .O(n2459));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1595_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i36281_2_lut_4_lut (.I0(n2367), .I1(n92), .I2(n2371), .I3(n96), 
            .O(n43406));
    defparam i36281_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_36_LessThan_1545_i18_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2367), 
            .I3(GND_net), .O(n18_adj_4762));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i22_3_lut_adj_1841 (.I0(bit_ctr[15]), .I1(n42966), .I2(n4754), 
            .I3(GND_net), .O(n35975));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1841.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_LessThan_1545_i20_3_lut_3_lut (.I0(n95_adj_4360), .I1(n94), 
            .I2(n2369), .I3(GND_net), .O(n20_adj_4764));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 unary_minus_18_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36203_2_lut_4_lut (.I0(n2359), .I1(n84), .I2(n2368), .I3(n93), 
            .O(n43327));
    defparam i36203_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_36_LessThan_1545_i22_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2359), 
            .I3(GND_net), .O(n22_adj_4766));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1545_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_36_LessThan_1606_i14_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2463), 
            .I3(GND_net), .O(n14_adj_4787));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_36_unary_minus_4_inv_0_i18_1_lut (.I0(gearBoxRatio[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4527));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36183_2_lut_4_lut (.I0(n2458), .I1(n92), .I2(n2462), .I3(n96), 
            .O(n43307));
    defparam i36183_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_36_LessThan_1606_i16_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2458), 
            .I3(GND_net), .O(n16_adj_4789));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_36_unary_minus_4_inv_0_i19_1_lut (.I0(gearBoxRatio[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4526));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_1606_i18_3_lut_3_lut (.I0(n95_adj_4360), .I1(n94), 
            .I2(n2460), .I3(GND_net), .O(n18_adj_4791));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i36136_2_lut_4_lut (.I0(n2450), .I1(n84), .I2(n2459), .I3(n93), 
            .O(n43260));
    defparam i36136_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_36_unary_minus_4_inv_0_i20_1_lut (.I0(gearBoxRatio[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4525));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_1830_i41_4_lut (.I0(n2702), .I1(n80), .I2(n7163), 
            .I3(n2724), .O(n41_adj_4904));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i41_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_LessThan_1830_i39_4_lut (.I0(n2703), .I1(n81), .I2(n7164), 
            .I3(n2724), .O(n39_adj_4903));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i39_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_mux_3_i1_3_lut (.I0(encoder0_position[0]), .I1(n25_adj_4364), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n391));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1830_i45_4_lut (.I0(n2700), .I1(n78), .I2(n7161), 
            .I3(n2724), .O(n45_adj_4906));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i45_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_LessThan_1830_i43_4_lut (.I0(n2701), .I1(n79), .I2(n7162), 
            .I3(n2724), .O(n43_adj_4905));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i43_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_LessThan_1830_i37_4_lut (.I0(n2704), .I1(n82), .I2(n7165), 
            .I3(n2724), .O(n37_adj_4902));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i37_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_LessThan_1830_i29_4_lut (.I0(n2708), .I1(n86), .I2(n7169), 
            .I3(n2724), .O(n29_adj_4897));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i29_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_LessThan_1830_i31_4_lut (.I0(n2707), .I1(n85), .I2(n7168), 
            .I3(n2724), .O(n31_adj_4899));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i31_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_LessThan_1830_i21_4_lut (.I0(n2712), .I1(n90), .I2(n7173), 
            .I3(n2724), .O(n21_adj_4892));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i21_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_LessThan_1830_i23_4_lut (.I0(n2711), .I1(n89), .I2(n7172), 
            .I3(n2724), .O(n23_adj_4893));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i23_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_LessThan_1830_i25_4_lut (.I0(n2710), .I1(n88), .I2(n7171), 
            .I3(n2724), .O(n25_adj_4895));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i25_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_LessThan_1830_i17_4_lut (.I0(n2714), .I1(n92), .I2(n7175), 
            .I3(n2724), .O(n17_adj_4890));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i17_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 i22_3_lut_adj_1842 (.I0(bit_ctr[14]), .I1(n42965), .I2(n4754), 
            .I3(GND_net), .O(n35973));   // verilog/neopixel.v(35[12] 117[6])
    defparam i22_3_lut_adj_1842.LUT_INIT = 16'hacac;
    SB_LUT4 div_36_LessThan_1830_i19_4_lut (.I0(n2713), .I1(n91), .I2(n7174), 
            .I3(n2724), .O(n19_adj_4891));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i19_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_LessThan_1830_i9_4_lut (.I0(n2718), .I1(n96), .I2(n7179), 
            .I3(n2724), .O(n9_adj_4883));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i9_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_LessThan_1830_i7_4_lut (.I0(n2719), .I1(n97), .I2(n7180), 
            .I3(n2724), .O(n7_adj_4881));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i7_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_LessThan_1830_i35_4_lut (.I0(n2705), .I1(n83), .I2(n7166), 
            .I3(n2724), .O(n35_adj_4901));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i35_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_LessThan_1830_i33_4_lut (.I0(n2706), .I1(n84), .I2(n7167), 
            .I3(n2724), .O(n33_adj_4900));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i33_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_LessThan_1830_i11_4_lut (.I0(n2717), .I1(n95_adj_4360), 
            .I2(n7178), .I3(n2724), .O(n11_adj_4885));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i11_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_LessThan_1830_i13_4_lut (.I0(n2716), .I1(n94), .I2(n7177), 
            .I3(n2724), .O(n13_adj_4887));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i13_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_LessThan_1830_i15_4_lut (.I0(n2715), .I1(n93), .I2(n7176), 
            .I3(n2724), .O(n15_adj_4888));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i15_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_LessThan_1830_i27_4_lut (.I0(n2709), .I1(n87), .I2(n7170), 
            .I3(n2724), .O(n27_adj_4896));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i27_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_36_i1832_1_lut (.I0(n2801), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2802));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1832_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36476_4_lut (.I0(n27_adj_4896), .I1(n15_adj_4888), .I2(n13_adj_4887), 
            .I3(n11_adj_4885), .O(n43601));
    defparam i36476_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_36_LessThan_1830_i12_3_lut (.I0(n93), .I1(n84), .I2(n33_adj_4900), 
            .I3(GND_net), .O(n12_adj_4886));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i36458_2_lut (.I0(n33_adj_4900), .I1(n15_adj_4888), .I2(GND_net), 
            .I3(GND_net), .O(n43583));
    defparam i36458_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_36_LessThan_1830_i10_3_lut (.I0(n95_adj_4360), .I1(n94), 
            .I2(n13_adj_4887), .I3(GND_net), .O(n10_adj_4884));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_36_LessThan_1830_i30_3_lut (.I0(n12_adj_4886), .I1(n83), 
            .I2(n35_adj_4901), .I3(GND_net), .O(n30_adj_4898));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_36_i1828_3_lut (.I0(n2720), .I1(n7181), .I2(n2724), .I3(GND_net), 
            .O(n2798));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36539_3_lut (.I0(n7_adj_4881), .I1(n2798), .I2(n98), .I3(GND_net), 
            .O(n43664));
    defparam i36539_3_lut.LUT_INIT = 16'hebeb;
    SB_LUT4 i37130_4_lut (.I0(n13_adj_4887), .I1(n11_adj_4885), .I2(n9_adj_4883), 
            .I3(n43664), .O(n44255));
    defparam i37130_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i37116_4_lut (.I0(n19_adj_4891), .I1(n17_adj_4890), .I2(n15_adj_4888), 
            .I3(n44255), .O(n44241));
    defparam i37116_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_36_i1646_3_lut_3_lut (.I0(n2471), .I1(n7095), .I2(n2451), 
            .I3(GND_net), .O(n2538));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1646_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i37809_4_lut (.I0(n25_adj_4895), .I1(n23_adj_4893), .I2(n21_adj_4892), 
            .I3(n44241), .O(n44934));
    defparam i37809_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i37390_4_lut (.I0(n31_adj_4899), .I1(n29_adj_4897), .I2(n27_adj_4896), 
            .I3(n44934), .O(n44515));
    defparam i37390_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i37895_4_lut (.I0(n37_adj_4902), .I1(n35_adj_4901), .I2(n33_adj_4900), 
            .I3(n44515), .O(n45020));
    defparam i37895_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_36_LessThan_1830_i16_3_lut (.I0(n91), .I1(n79), .I2(n43_adj_4905), 
            .I3(GND_net), .O(n16_adj_4889));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_36_LessThan_1830_i6_3_lut (.I0(n98), .I1(n97), .I2(n7_adj_4881), 
            .I3(GND_net), .O(n6_adj_4880));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i37454_3_lut (.I0(n6_adj_4880), .I1(n90), .I2(n21_adj_4892), 
            .I3(GND_net), .O(n44579));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37454_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37455_3_lut (.I0(n44579), .I1(n89), .I2(n23_adj_4893), .I3(GND_net), 
            .O(n44580));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37455_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36497_4_lut (.I0(n21_adj_4892), .I1(n19_adj_4891), .I2(n17_adj_4890), 
            .I3(n9_adj_4883), .O(n43622));
    defparam i36497_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36412_2_lut (.I0(n43_adj_4905), .I1(n19_adj_4891), .I2(GND_net), 
            .I3(GND_net), .O(n43537));
    defparam i36412_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_36_i1643_3_lut_3_lut (.I0(n2471), .I1(n7092), .I2(n2448), 
            .I3(GND_net), .O(n2535));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1643_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1642_3_lut_3_lut (.I0(n2471), .I1(n7091), .I2(n2447), 
            .I3(GND_net), .O(n2534));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1642_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1644_3_lut_3_lut (.I0(n2471), .I1(n7093), .I2(n2449), 
            .I3(GND_net), .O(n2536));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1644_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1645_3_lut_3_lut (.I0(n2471), .I1(n7094), .I2(n2450), 
            .I3(GND_net), .O(n2537));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1645_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_LessThan_1830_i8_3_lut (.I0(n96), .I1(n92), .I2(n17_adj_4890), 
            .I3(GND_net), .O(n8_adj_4882));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_36_LessThan_1830_i24_3_lut (.I0(n16_adj_4889), .I1(n78), 
            .I2(n45_adj_4906), .I3(GND_net), .O(n24_adj_4894));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_36_i1661_3_lut_3_lut (.I0(n2471), .I1(n7110), .I2(n387), 
            .I3(GND_net), .O(n2553));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1661_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1650_3_lut_3_lut (.I0(n2471), .I1(n7099), .I2(n2455), 
            .I3(GND_net), .O(n2542));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1650_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i36414_4_lut (.I0(n43_adj_4905), .I1(n25_adj_4895), .I2(n23_adj_4893), 
            .I3(n43622), .O(n43539));
    defparam i36414_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_36_i1651_3_lut_3_lut (.I0(n2471), .I1(n7100), .I2(n2456), 
            .I3(GND_net), .O(n2543));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1651_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i37579_4_lut (.I0(n24_adj_4894), .I1(n8_adj_4882), .I2(n45_adj_4906), 
            .I3(n43537), .O(n44704));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37579_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36877_3_lut (.I0(n44580), .I1(n88), .I2(n25_adj_4895), .I3(GND_net), 
            .O(n44002));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36877_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_36_i1829_3_lut (.I0(n390), .I1(n7182), .I2(n2724), .I3(GND_net), 
            .O(n2799));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1830_i4_4_lut (.I0(n391), .I1(n99), .I2(n2799), 
            .I3(n558), .O(n4_adj_4879));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1830_i4_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_36_i1652_3_lut_3_lut (.I0(n2471), .I1(n7101), .I2(n2457), 
            .I3(GND_net), .O(n2544));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1652_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i37450_3_lut (.I0(n4_adj_4879), .I1(n87), .I2(n27_adj_4896), 
            .I3(GND_net), .O(n44575));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37450_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37451_3_lut (.I0(n44575), .I1(n86), .I2(n29_adj_4897), .I3(GND_net), 
            .O(n44576));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37451_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_36_i1653_3_lut_3_lut (.I0(n2471), .I1(n7102), .I2(n2458), 
            .I3(GND_net), .O(n2545));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1653_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1654_3_lut_3_lut (.I0(n2471), .I1(n7103), .I2(n2459), 
            .I3(GND_net), .O(n2546));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1654_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i36462_4_lut (.I0(n33_adj_4900), .I1(n31_adj_4899), .I2(n29_adj_4897), 
            .I3(n43601), .O(n43587));
    defparam i36462_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37793_4_lut (.I0(n30_adj_4898), .I1(n10_adj_4884), .I2(n35_adj_4901), 
            .I3(n43583), .O(n44918));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37793_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36879_3_lut (.I0(n44576), .I1(n85), .I2(n31_adj_4899), .I3(GND_net), 
            .O(n44004));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36879_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37969_4_lut (.I0(n44004), .I1(n44918), .I2(n35_adj_4901), 
            .I3(n43587), .O(n45094));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37969_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i37970_3_lut (.I0(n45094), .I1(n82), .I2(n37_adj_4902), .I3(GND_net), 
            .O(n45095));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37970_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37923_3_lut (.I0(n45095), .I1(n81), .I2(n39_adj_4903), .I3(GND_net), 
            .O(n45048));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37923_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36427_4_lut (.I0(n43_adj_4905), .I1(n41_adj_4904), .I2(n39_adj_4903), 
            .I3(n45020), .O(n43552));
    defparam i36427_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_36_i1648_3_lut_3_lut (.I0(n2471), .I1(n7097), .I2(n2453), 
            .I3(GND_net), .O(n2540));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1648_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1656_3_lut_3_lut (.I0(n2471), .I1(n7105), .I2(n2461), 
            .I3(GND_net), .O(n2548));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1656_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i37883_4_lut (.I0(n44002), .I1(n44704), .I2(n45_adj_4906), 
            .I3(n43539), .O(n45008));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37883_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36885_3_lut (.I0(n45048), .I1(n80), .I2(n41_adj_4904), .I3(GND_net), 
            .O(n44010));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i36885_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_36_i1807_3_lut (.I0(n2699), .I1(n7160), .I2(n2724), .I3(GND_net), 
            .O(n2777));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1649_3_lut_3_lut (.I0(n2471), .I1(n7098), .I2(n2454), 
            .I3(GND_net), .O(n2541));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1649_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i37885_4_lut (.I0(n44010), .I1(n45008), .I2(n45_adj_4906), 
            .I3(n43552), .O(n45010));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37885_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i37886_3_lut (.I0(n45010), .I1(n77), .I2(n2777), .I3(GND_net), 
            .O(n2801));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37886_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 div_36_i1660_3_lut_3_lut (.I0(n2471), .I1(n7109), .I2(n2465), 
            .I3(GND_net), .O(n2552));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1660_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_LessThan_1606_i20_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2450), 
            .I3(GND_net), .O(n20_adj_4793));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1606_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_36_i1659_3_lut_3_lut (.I0(n2471), .I1(n7108), .I2(n2464), 
            .I3(GND_net), .O(n2551));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1659_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_LessThan_1777_i33_2_lut (.I0(n2706), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4876));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1777_i31_2_lut (.I0(n2707), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4874));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1777_i37_2_lut (.I0(n2704), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4878));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1777_i35_2_lut (.I0(n2705), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4877));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_mux_3_i2_3_lut (.I0(encoder0_position[1]), .I1(n24), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n390));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_i1658_3_lut_3_lut (.I0(n2471), .I1(n7107), .I2(n2463), 
            .I3(GND_net), .O(n2550));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1658_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1647_3_lut_3_lut (.I0(n2471), .I1(n7096), .I2(n2452), 
            .I3(GND_net), .O(n2539));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1647_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_i1655_3_lut_3_lut (.I0(n2471), .I1(n7104), .I2(n2460), 
            .I3(GND_net), .O(n2547));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1655_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_LessThan_1777_i25_2_lut (.I0(n2710), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4870));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_i1657_3_lut_3_lut (.I0(n2471), .I1(n7106), .I2(n2462), 
            .I3(GND_net), .O(n2549));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1657_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_36_LessThan_1777_i27_2_lut (.I0(n2709), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4871));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1777_i21_2_lut (.I0(n2712), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4867));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1777_i23_2_lut (.I0(n2711), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4868));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1777_i9_2_lut (.I0(n2718), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_4858));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i9_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1665_i12_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2551), 
            .I3(GND_net), .O(n12_adj_4809));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i36081_2_lut_4_lut (.I0(n2546), .I1(n92), .I2(n2550), .I3(n96), 
            .O(n43205));
    defparam i36081_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_36_LessThan_1665_i14_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2546), 
            .I3(GND_net), .O(n14_adj_4811));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_36_LessThan_1777_i13_2_lut (.I0(n2716), .I1(n95_adj_4360), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4862));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1777_i15_2_lut (.I0(n2715), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4864));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1777_i17_2_lut (.I0(n2714), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4865));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1777_i29_2_lut (.I0(n2708), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4872));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1665_i16_3_lut_3_lut (.I0(n95_adj_4360), .I1(n94), 
            .I2(n2548), .I3(GND_net), .O(n16_adj_4813));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_36_LessThan_1777_i11_2_lut (.I0(n2717), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4860));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1777_i19_2_lut (.I0(n2713), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4866));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_i1779_1_lut (.I0(n2723), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1779_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35886_4_lut (.I0(n29_adj_4872), .I1(n17_adj_4865), .I2(n15_adj_4864), 
            .I3(n13_adj_4862), .O(n43010));
    defparam i35886_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36652_4_lut (.I0(n11_adj_4860), .I1(n9_adj_4858), .I2(n2719), 
            .I3(n98), .O(n43777));
    defparam i36652_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i37200_4_lut (.I0(n17_adj_4865), .I1(n15_adj_4864), .I2(n13_adj_4862), 
            .I3(n43777), .O(n44325));
    defparam i37200_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i37196_4_lut (.I0(n23_adj_4868), .I1(n21_adj_4867), .I2(n19_adj_4866), 
            .I3(n44325), .O(n44321));
    defparam i37196_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35888_4_lut (.I0(n29_adj_4872), .I1(n27_adj_4871), .I2(n25_adj_4870), 
            .I3(n44321), .O(n43012));
    defparam i35888_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_36_LessThan_1777_i6_4_lut (.I0(n390), .I1(n99), .I2(n2720), 
            .I3(n558), .O(n6_adj_4856));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i6_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i37683_3_lut (.I0(n6_adj_4856), .I1(n87), .I2(n29_adj_4872), 
            .I3(GND_net), .O(n44808));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37683_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_36_LessThan_1777_i32_3_lut (.I0(n14_adj_4863), .I1(n83), 
            .I2(n37_adj_4878), .I3(GND_net), .O(n32_adj_4875));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1777_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37684_3_lut (.I0(n44808), .I1(n86), .I2(n31_adj_4874), .I3(GND_net), 
            .O(n44809));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37684_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35876_4_lut (.I0(n35_adj_4877), .I1(n33_adj_4876), .I2(n31_adj_4874), 
            .I3(n43010), .O(n43000));
    defparam i35876_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37787_4_lut (.I0(n32_adj_4875), .I1(n12_adj_4861), .I2(n37_adj_4878), 
            .I3(n43718), .O(n44912));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37787_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i37578_3_lut (.I0(n44809), .I1(n85), .I2(n33_adj_4876), .I3(GND_net), 
            .O(n30_adj_4873));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37578_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37685_3_lut (.I0(n8_adj_4857), .I1(n90), .I2(n23_adj_4868), 
            .I3(GND_net), .O(n44810));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37685_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37686_3_lut (.I0(n44810), .I1(n89), .I2(n25_adj_4870), .I3(GND_net), 
            .O(n44811));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37686_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36628_4_lut (.I0(n25_adj_4870), .I1(n23_adj_4868), .I2(n21_adj_4867), 
            .I3(n43028), .O(n43753));
    defparam i36628_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i37575_3_lut (.I0(n10_adj_4859), .I1(n91), .I2(n21_adj_4867), 
            .I3(GND_net), .O(n44700));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37575_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37574_3_lut (.I0(n44811), .I1(n88), .I2(n27_adj_4871), .I3(GND_net), 
            .O(n24_adj_4869));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37574_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37432_4_lut (.I0(n35_adj_4877), .I1(n33_adj_4876), .I2(n31_adj_4874), 
            .I3(n43012), .O(n44557));
    defparam i37432_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i37905_4_lut (.I0(n30_adj_4873), .I1(n44912), .I2(n37_adj_4878), 
            .I3(n43000), .O(n45030));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37905_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i37671_4_lut (.I0(n24_adj_4869), .I1(n44700), .I2(n27_adj_4871), 
            .I3(n43753), .O(n44796));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37671_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i37999_4_lut (.I0(n44796), .I1(n45030), .I2(n37_adj_4878), 
            .I3(n44557), .O(n45124));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37999_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i38000_3_lut (.I0(n45124), .I1(n82), .I2(n2703), .I3(GND_net), 
            .O(n45125));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i38000_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i37996_3_lut (.I0(n45125), .I1(n81), .I2(n2702), .I3(GND_net), 
            .O(n45121));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37996_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i37849_3_lut (.I0(n45121), .I1(n80), .I2(n2701), .I3(GND_net), 
            .O(n44974));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37849_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i37850_3_lut (.I0(n44974), .I1(n79), .I2(n2700), .I3(GND_net), 
            .O(n44975));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37850_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1964_4_lut (.I0(n44975), .I1(n77), .I2(n78), .I3(n2699), 
            .O(n2723));
    defparam i1964_4_lut.LUT_INIT = 16'hceef;
    SB_LUT4 i36048_2_lut_4_lut (.I0(n2538), .I1(n84), .I2(n2547), .I3(n93), 
            .O(n43172));
    defparam i36048_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_36_unary_minus_4_inv_0_i21_1_lut (.I0(gearBoxRatio[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4524));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_4_inv_0_i22_1_lut (.I0(gearBoxRatio[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4523));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_LessThan_1665_i18_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2538), 
            .I3(GND_net), .O(n18_adj_4815));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1665_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i14394_3_lut_4_lut (.I0(r_SM_Main_adj_5046[2]), .I1(r_SM_Main_2__N_3320[1]), 
            .I2(r_SM_Main_adj_5046[0]), .I3(r_SM_Main_adj_5046[1]), .O(n19426));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i14394_3_lut_4_lut.LUT_INIT = 16'h1540;
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.n19395(n19395), .encoder1_position({encoder1_position}), 
            .clk32MHz(clk32MHz), .n19396(n19396), .n19397(n19397), .n19398(n19398), 
            .n19399(n19399), .n19400(n19400), .n19401(n19401), .n19387(n19387), 
            .n19388(n19388), .n19389(n19389), .n19390(n19390), .n19391(n19391), 
            .n19392(n19392), .n19393(n19393), .n19394(n19394), .n19383(n19383), 
            .n19384(n19384), .n19385(n19385), .n19386(n19386), .n19379(n19379), 
            .n19380(n19380), .n19381(n19381), .n19382(n19382), .data_o({quadA_debounced_adj_4372, 
            quadB_debounced_adj_4373}), .GND_net(GND_net), .n2815({n2816, 
            n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, 
            n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, 
            n2833, n2834, n2835, n2836, n2837, n2838, n2839}), 
            .n18804(n18804), .count_enable(count_enable_adj_4374), .n19450(n19450), 
            .PIN_6_c_0(PIN_6_c_0), .reg_B({reg_B_adj_5057}), .PIN_7_c_1(PIN_7_c_1), 
            .n18830(n18830), .n39886(n39886)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(255[15] 260[4])
    SB_LUT4 div_36_LessThan_1722_i45_2_lut (.I0(n2619), .I1(n80), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4855));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1722_i41_2_lut (.I0(n2621), .I1(n82), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4852));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1722_i43_2_lut (.I0(n2620), .I1(n81), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4853));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_mux_3_i3_3_lut (.I0(encoder0_position[2]), .I1(n23), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n389));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_36_LessThan_1722_i33_2_lut (.I0(n2625), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4847));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1722_i35_2_lut (.I0(n2624), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4849));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1722_i27_2_lut (.I0(n2628), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4844));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1722_i29_2_lut (.I0(n2627), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4845));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1722_i23_2_lut (.I0(n2630), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4842));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1722_i25_2_lut (.I0(n2629), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4843));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1722_i11_2_lut (.I0(n2636), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4832));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1722_i39_2_lut (.I0(n2622), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4851));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1722_i37_2_lut (.I0(n2623), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4850));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1722_i15_2_lut (.I0(n2634), .I1(n95_adj_4360), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4836));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1722_i17_2_lut (.I0(n2633), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4838));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1722_i19_2_lut (.I0(n2632), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_4839));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1722_i31_2_lut (.I0(n2626), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4846));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1722_i13_2_lut (.I0(n2635), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_4834));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_LessThan_1722_i21_2_lut (.I0(n2631), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_4841));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_36_i1724_1_lut (.I0(n2642), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2643));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_i1724_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35950_4_lut (.I0(n31_adj_4846), .I1(n19_adj_4839), .I2(n17_adj_4838), 
            .I3(n15_adj_4836), .O(n43074));
    defparam i35950_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_36_LessThan_1722_i34_3_lut (.I0(n16_adj_4837), .I1(n83), 
            .I2(n39_adj_4851), .I3(GND_net), .O(n34_adj_4848));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36714_4_lut (.I0(n13_adj_4834), .I1(n11_adj_4832), .I2(n2637), 
            .I3(n98), .O(n43839));
    defparam i36714_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i37228_4_lut (.I0(n19_adj_4839), .I1(n17_adj_4838), .I2(n15_adj_4836), 
            .I3(n43839), .O(n44353));
    defparam i37228_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i37222_4_lut (.I0(n25_adj_4843), .I1(n23_adj_4842), .I2(n21_adj_4841), 
            .I3(n44353), .O(n44347));
    defparam i37222_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35955_4_lut (.I0(n31_adj_4846), .I1(n29_adj_4845), .I2(n27_adj_4844), 
            .I3(n44347), .O(n43079));
    defparam i35955_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37444_4_lut (.I0(n37_adj_4850), .I1(n35_adj_4849), .I2(n33_adj_4847), 
            .I3(n43079), .O(n44569));
    defparam i37444_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i37757_3_lut (.I0(n10_adj_4831), .I1(n90), .I2(n25_adj_4843), 
            .I3(GND_net), .O(n44882));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37757_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37758_3_lut (.I0(n44882), .I1(n89), .I2(n27_adj_4844), .I3(GND_net), 
            .O(n44883));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37758_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36690_4_lut (.I0(n27_adj_4844), .I1(n25_adj_4843), .I2(n23_adj_4842), 
            .I3(n43101), .O(n43815));
    defparam i36690_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_36_LessThan_1722_i20_3_lut (.I0(n12_adj_4833), .I1(n91), 
            .I2(n23_adj_4842), .I3(GND_net), .O(n20_adj_4840));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37564_3_lut (.I0(n44883), .I1(n88), .I2(n29_adj_4845), .I3(GND_net), 
            .O(n44689));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37564_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_36_LessThan_1722_i8_4_lut (.I0(n389), .I1(n99), .I2(n2638), 
            .I3(n558), .O(n8_adj_4830));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_LessThan_1722_i8_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i37693_3_lut (.I0(n8_adj_4830), .I1(n87), .I2(n31_adj_4846), 
            .I3(GND_net), .O(n44818));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37693_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37694_3_lut (.I0(n44818), .I1(n86), .I2(n33_adj_4847), .I3(GND_net), 
            .O(n44819));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37694_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35944_4_lut (.I0(n37_adj_4850), .I1(n35_adj_4849), .I2(n33_adj_4847), 
            .I3(n43074), .O(n43068));
    defparam i35944_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37916_4_lut (.I0(n34_adj_4848), .I1(n14_adj_4835), .I2(n39_adj_4851), 
            .I3(n43066), .O(n45041));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37916_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i37566_3_lut (.I0(n44819), .I1(n85), .I2(n35_adj_4849), .I3(GND_net), 
            .O(n44691));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37566_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37987_4_lut (.I0(n44691), .I1(n45041), .I2(n39_adj_4851), 
            .I3(n43068), .O(n45112));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37987_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i37988_3_lut (.I0(n45112), .I1(n82), .I2(n41_adj_4852), .I3(GND_net), 
            .O(n45113));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37988_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37960_3_lut (.I0(n45113), .I1(n81), .I2(n43_adj_4853), .I3(GND_net), 
            .O(n45085));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37960_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37918_4_lut (.I0(n43_adj_4853), .I1(n41_adj_4852), .I2(n39_adj_4851), 
            .I3(n44569), .O(n45043));
    defparam i37918_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i37569_4_lut (.I0(n44689), .I1(n20_adj_4840), .I2(n29_adj_4845), 
            .I3(n43815), .O(n44694));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37569_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i37942_3_lut (.I0(n45085), .I1(n80), .I2(n45_adj_4855), .I3(GND_net), 
            .O(n44_adj_4854));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37942_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i37571_4_lut (.I0(n44_adj_4854), .I1(n44694), .I2(n45_adj_4855), 
            .I3(n45043), .O(n44696));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam i37571_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1843 (.I0(n44696), .I1(n17244), .I2(n79), .I3(n2618), 
            .O(n2642));
    defparam i1_4_lut_adj_1843.LUT_INIT = 16'hceef;
    SB_LUT4 unary_minus_18_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4328));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_4_inv_0_i23_1_lut (.I0(gearBoxRatio[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4522));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_18_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4327));   // verilog/TinyFPGA_B.v(137[23:28])
    defparam unary_minus_18_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_36_unary_minus_4_inv_0_i24_1_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2_adj_4521));   // verilog/TinyFPGA_B.v(243[21:53])
    defparam div_36_unary_minus_4_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    motorControl control (.\Kp[4] (Kp[4]), .\Kp[2] (Kp[2]), .GND_net(GND_net), 
            .\Kp[3] (Kp[3]), .\Kp[0] (Kp[0]), .\Kp[1] (Kp[1]), .\Kp[5] (Kp[5]), 
            .duty({duty}), .PWMLimit({PWMLimit}), .\Ki[7] (Ki[7]), .IntegralLimit({IntegralLimit}), 
            .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), .\Ki[1] (Ki[1]), .\Ki[0] (Ki[0]), 
            .\Ki[2] (Ki[2]), .\Ki[3] (Ki[3]), .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), 
            .\Ki[6] (Ki[6]), .clk32MHz(clk32MHz), .VCC_net(VCC_net), .n25(n25), 
            .motor_state({motor_state}), .setpoint({setpoint}), .n45865(n45865)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(227[16] 240[4])
    \pwm(32000000,20000,32000000,23,1)  PWM (.pwm_setpoint({pwm_setpoint}), 
            .GND_net(GND_net), .\half_duty_new[0] (half_duty_new[0]), .CLK_c(CLK_c), 
            .PIN_19_c_0(PIN_19_c_0), .n19420(n19420), .\half_duty[0][2] (\half_duty[0] [2]), 
            .n19421(n19421), .\half_duty[0][3] (\half_duty[0] [3]), .n19422(n19422), 
            .\half_duty[0][4] (\half_duty[0] [4]), .n19423(n19423), .\half_duty[0][5] (\half_duty[0] [5]), 
            .n19424(n19424), .\half_duty[0][6] (\half_duty[0] [6]), .n19425(n19425), 
            .\half_duty[0][7] (\half_duty[0] [7]), .n19414(n19414), .\half_duty[0][1] (\half_duty[0] [1]), 
            .n1111(n1111), .VCC_net(VCC_net), .\half_duty_new[1] (half_duty_new[1]), 
            .\half_duty[0][0] (\half_duty[0] [0]), .\half_duty_new[2] (half_duty_new[2]), 
            .\half_duty_new[3] (half_duty_new[3]), .\half_duty_new[4] (half_duty_new[4]), 
            .\half_duty_new[5] (half_duty_new[5]), .\half_duty_new[6] (half_duty_new[6]), 
            .\half_duty_new[7] (half_duty_new[7]), .n18810(n18810)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(119[43] 125[3])
    
endmodule
//
// Verilog Description of module neopixel
//

module neopixel (timer, GND_net, \neo_pixel_transmitter.done , clk32MHz, 
            n42947, bit_ctr, n19, n42956, n35971, n35973, n35975, 
            n35967, n35969, n35963, n35965, n35959, n35961, n35955, 
            n35957, n35951, n35953, n35947, n35949, n35933, n35935, 
            n35937, n35939, n35941, n35943, n35931, n35925, n35907, 
            VCC_net, n35927, n35909, n35911, n35929, \neo_pixel_transmitter.t0 , 
            \one_wire_N_513[11] , n42943, n10, n42966, \one_wire_N_513[7] , 
            n8, n42955, \one_wire_N_513[5] , n42965, n42964, n42954, 
            n38094, \state[1] , n42963, start, n42968, n42962, n35923, 
            n42953, n42961, \state_3__N_362[1] , n27365, n17195, n38070, 
            n35913, n35917, n35915, n18886, n18885, n18884, n18883, 
            n18882, n18881, n18880, n18879, n18878, n18877, n18876, 
            n18875, n18874, n18873, n18872, n18871, n18870, n18869, 
            n18868, n18867, n18866, n18865, n18864, n18863, n18862, 
            n18861, n18860, n18859, n18858, n18857, n18856, n18855, 
            \state[0] , n38192, n42960, n42952, n18416, n18584, 
            n42959, n42951, n42950, n35977, n42946, n42945, PIN_8_c, 
            n42939, n11, n42940, n42958, n42936, n42935, n18663, 
            n42934, n42957, n42933, n42944, n42942, n42941, n42949, 
            n42948, n1105, n4754, n27453, n39307, \color[20] , \color[21] , 
            \color[17] ) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [31:0]timer;
    input GND_net;
    output \neo_pixel_transmitter.done ;
    input clk32MHz;
    output n42947;
    output [31:0]bit_ctr;
    input n19;
    output n42956;
    input n35971;
    input n35973;
    input n35975;
    input n35967;
    input n35969;
    input n35963;
    input n35965;
    input n35959;
    input n35961;
    input n35955;
    input n35957;
    input n35951;
    input n35953;
    input n35947;
    input n35949;
    input n35933;
    input n35935;
    input n35937;
    input n35939;
    input n35941;
    input n35943;
    input n35931;
    input n35925;
    input n35907;
    input VCC_net;
    input n35927;
    input n35909;
    input n35911;
    input n35929;
    output [31:0]\neo_pixel_transmitter.t0 ;
    output \one_wire_N_513[11] ;
    output n42943;
    output n10;
    output n42966;
    output \one_wire_N_513[7] ;
    output n8;
    output n42955;
    output \one_wire_N_513[5] ;
    output n42965;
    output n42964;
    output n42954;
    input n38094;
    output \state[1] ;
    output n42963;
    output start;
    output n42968;
    output n42962;
    input n35923;
    output n42953;
    output n42961;
    output \state_3__N_362[1] ;
    output n27365;
    output n17195;
    output n38070;
    input n35913;
    input n35917;
    input n35915;
    input n18886;
    input n18885;
    input n18884;
    input n18883;
    input n18882;
    input n18881;
    input n18880;
    input n18879;
    input n18878;
    input n18877;
    input n18876;
    input n18875;
    input n18874;
    input n18873;
    input n18872;
    input n18871;
    input n18870;
    input n18869;
    input n18868;
    input n18867;
    input n18866;
    input n18865;
    input n18864;
    input n18863;
    input n18862;
    input n18861;
    input n18860;
    input n18859;
    input n18858;
    input n18857;
    input n18856;
    input n18855;
    output \state[0] ;
    input n38192;
    output n42960;
    output n42952;
    output n18416;
    output n18584;
    output n42959;
    output n42951;
    output n42950;
    input n35977;
    output n42946;
    output n42945;
    output PIN_8_c;
    output n42939;
    input n11;
    output n42940;
    output n42958;
    output n42936;
    output n42935;
    input n18663;
    output n42934;
    output n42957;
    output n42933;
    output n42944;
    output n42942;
    output n42941;
    output n42949;
    output n42948;
    output n1105;
    output n4754;
    output n27453;
    output n39307;
    input \color[20] ;
    input \color[21] ;
    input \color[17] ;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n2690, n2591, n2621, n31688, n30418;
    wire [31:0]n1;
    
    wire n30419;
    wire [31:0]n133;
    
    wire n31157, n31689, \neo_pixel_transmitter.done_N_570 , n39942, 
        n2691, n2592, n31687, n24, n30417;
    wire [31:0]one_wire_N_513;
    
    wire n31158, n2692, n2593, n31686, n2693, n2594, n31685, n2694, 
        n2595, n31684, n31156, n30275, n2695, n2596, n31683, n2696, 
        n2597, n31682, n31155, n6, n30416, n31154, n30263, n5, 
        n30415, n2697, n2598, n31681, n2698, n2599, n31680, n2699, 
        n2600, n31679, n2700, n2601, n31678, n2701, n2602, n31677, 
        n2702, n2603, n31676, n2703, n2604, n31675, n20, n30414, 
        n2704, n2605, n31674, n31153, n31152, n31151, n31150, 
        n2302, n2292, n2293, n2301, n30, n2309, n27219, n2294, 
        n2306, n2304, n34, n2291, n2303, n2305, n32, n2298, 
        n2295, n2296, n2300, n33, n2308, n2297, n2307, n2299, 
        n31, n2324, n31149, n31148, n2423, n45855, n31147, n2705, 
        n2606, n31673, n2403, n2409, n27, n2390, n2391, n2397, 
        n2394, n33_adj_4196, n2392, n2405, n2400, n2398, n32_adj_4197, 
        n2396, n2402, n2408, n2399, n31_adj_4198, n2393, n2406, 
        n2395, n2407, n35, n2404, n2401, n37, n31146, n31145, 
        n31144, n2522, n45854, n26, n30413, n18_adj_4200, n2706, 
        n2607, n31672, n30412, n30276, n2707, n2608, n31671, n30411, 
        n2708, n2609, n45853, n31670, n2709, n2588, n2489, n31669, 
        n30274, n2589, n2490, n31668, n2590, n2491, n31667, n30410, 
        n2492, n31666, n30409, n708, n2493, n31665, n2494, n31664, 
        n2495, n31663, n2496, n31662, n2497, n31661, n2498, n31660, 
        n30264, n30273, n15780, n38037, n60, n2499, n31659, n2009, 
        n27237, n838, n38039, n2000, n1999, n2007, n2003, n28_adj_4203, 
        n2500, n31658, n2501, n31657, n30408, n1996, n1994, n2006, 
        n26_adj_4204, n1997, n2001, n1995, n2008, n27_adj_4205, 
        n2502, n31656, n2004, n2002, n2005, n1998, n25_adj_4206, 
        n2027, n2503, n31655, n2504, n31654, n30407, n30262, n30406, 
        n2505, n31653, n2506, n31652, n2507, n31651, n2508, n31650, 
        n30272, n2509, n31649, n30405, n31648, n31647, n2126, 
        n45858, n31646, n31645, n31644, n31643, n31642, n30404, 
        n31641, n31640, n31639, n31638, n31637, n31636, n31635, 
        n30403, n31634, n31633, n31632, n31631, n31630, n31629, 
        n32659, n30402, n4, n31628, n31627, n31626, n31625, n31624, 
        n31623, n31622, n31621, n31620, n31619, n31618, n31617, 
        n31616, n30271, n31615, n31614, n31613, n31612, n31611, 
        n45856, n31610, n2192, n2225, n31609, n2193, n31608, n2194, 
        n31607, n2195, n31606, n2196, n31605, n2197, n31604, n2198, 
        n31603, n2199, n31602, n2200, n31601, n2201, n31600, n24_adj_4208, 
        n34_adj_4209, n22_adj_4210, n38, n30261, n36, n2202, n31599, 
        n2203, n31598, n37_adj_4211, n2204, n31597, n35_adj_4212, 
        n27335, n17206, n38456, n2205, n31596, n2206, n31595, 
        n2207, n31594, n30270, n2208, n31593, n2209, n45857, n31592, 
        n2093, n31591, n2094, n31590, n1108, n2095, n31589, n2096, 
        n31588, n2097, n31587, n2098, n31586, n2099, n31585, n2100, 
        n31584, n2101, n31583, n30269, n2102, n31582, n2103, n31581, 
        n2104, n31580, n2105, n31579, n27_adj_4213, n2106, n31578, 
        n30260, n2107, n31577, n2108, n31576, n30268, n2109, n31575, 
        n31574, n31573, n31572, n31571, n31570, n31569, n31568, 
        n31567, n17196, n4724, n27164, n29_adj_4214, n28_adj_4215, 
        n32476, n17064, n27172, n4_adj_4216, n14, n31566, n31565, 
        n18_adj_4217, n31564, n30_adj_4218, n31563, n28_adj_4219, 
        n29_adj_4220, n31562, n27_adj_4221, n31561, n31560, n45859, 
        n31559, n1895, n1928, n31558, n1896, n31557, n1897, n31556, 
        n1898, n31555, n1899, n31554, n1900, n31553, n1901, n31552, 
        n1902, n31551, n1903, n31550, n1904, n31549, n1905, n31548, 
        n1906, n31547, n1907, n31546, n1908, n31545, n1909, n45860, 
        n31544, n37332, n21_adj_4222, n22_adj_4223, n28_adj_4224, 
        n23_adj_4225, n25_adj_4226, n32_adj_4227, n19_adj_4228, n5_adj_4229, 
        n38086, n37374, n116, n26_adj_4230, n36_adj_4231, n34_adj_4232, 
        n40, n38_adj_4233, n39, n37_adj_4234, n1796, n1829, n31543, 
        n1797, n31542, n1798, n31541, n1799, n31540, n1800, n31539, 
        n1801, n31538, n1802, n31537, n30267, n1803, n31536, n1804, 
        n31535, n1805, n31534, n3182, n3083, n3116, n31816, n1806, 
        n31533, n3183, n3084, n31815, n1807, n31532, n3184, n3085, 
        n31814, n1808, n31531, n3185, n3086, n31813, n1809, n45861, 
        n31530, n3186, n3087, n31812, n3187, n3088, n31811, n1697, 
        n1730, n31529, n1698, n31528, n3188, n3089, n31810, n1699, 
        n31527, n3189, n3090, n31809, n1700, n31526, n3190, n3091, 
        n31808, n1701, n31525, n3191, n3092, n31807, n1702, n31524, 
        n3192, n3093, n31806, n1703, n31523, n3193, n3094, n31805, 
        n1704, n31522, n3194, n3095, n31804, n1705, n31521, n1706, 
        n31520, n3195, n3096, n31803, n3196, n3097, n31802, n1707, 
        n31519, n22_adj_4235, n1708, n20_adj_4236, n21_adj_4237, n1709, 
        n19_adj_4238, n3197, n3098, n31801, n31518, n45864, n31517, 
        n30259, n3198, n3099, n31800, n1598, n1631, n31516, n3199, 
        n3100, n31799, n1599, n31515, n1600, n31514, n3200, n3101, 
        n31798, n1601, n31513, n3201, n3102, n31797, n1602, n31512, 
        n3202, n3103, n31796, n1603, n31511, n3203, n3104, n31795, 
        n1604, n31510, n3204, n3105, n31794, n1605, n31509;
    wire [3:0]state_3__N_362;
    
    wire n1606, n31508, n3205, n3106, n31793, n1607, n31507, n3206, 
        n3107, n31792, n1608, n31506, n3207, n3108, n31791, n30266, 
        n1609, n45866, n31505, n3208, n3109, n45863, n31790, n1499, 
        n1532, n31504, n3209, n1500, n31503, n2984, n3017, n31789, 
        n30289, n2985, n31788, n1501, n31502, n1502, n31501, n2986, 
        n31787, n2987, n31786, n1503, n31500, n2988, n31785, n1504, 
        n31499, n2989, n31784, n1505, n31498, n2990, n31783, n1506, 
        n31497, n2991, n31782, n1507, n31496, n2992, n31781, n1508, 
        n31495, n2993, n31780, n1509, n45867, n31494, n2994, n31779, 
        n1400, n1433, n31493, n2995, n31778, n1401, n31492, n2996, 
        n31777, n1402, n31491, n30288, n1403, n31490, n2997, n31776, 
        n2998, n31775, n1404, n31489, n1405, n31488, n2999, n31774, 
        n3000, n31773, n1406, n31487, n3001, n31772, n1407, n31486, 
        n3002, n31771, n1408, n31485, n3003, n31770, n1409, n45869, 
        n31484, n3004, n31769, n3005, n31768, n3006, n31767, n1301, 
        n1334, n31483, n1302, n31482, n1303, n31481, n1304, n31480, 
        n3007, n31766, n1305, n31479, n3008, n31765, n3009, n45868, 
        n31764, n1306, n31478, n1307, n31477, n1308, n31476, n2885, 
        n2918, n31763, n2886, n31762, n2887, n31761, n1309, n45870, 
        n31475, n2888, n31760, n1202, n1235, n31474, n1203, n31473, 
        n1204, n31472, n2889, n31759, n2890, n31758, n1205, n31471, 
        n30287, n2891, n31757, n1206, n31470, n2892, n31756, n1207, 
        n31469, n1208, n31468, n2893, n31755, n1209, n45872, n31467, 
        n2894, n31754, n1103, n1136, n31466, n1104, n31465, n2895, 
        n31753, n1105_adj_4239, n31464, n30286, n2896, n31752, n1106, 
        n31463, n2897, n31751, n2898, n31750, n1107, n31462, n1108_adj_4240, 
        n31461, n2899, n31749, n2900, n31748, n1109, n45873, n31460, 
        n2901, n31747, n2902, n31746, n4_adj_4241, n1037, n31459, 
        n1005, n31458, n2903, n31745, n1006, n31457, n2904, n31744, 
        n2905, n31743, n1007, n31456, n2906, n31742, n1008, n31455, 
        n1009, n45874, n31454, n2907, n31741, n2908, n31740;
    wire [31:0]n971;
    
    wire n905, n31453, n2909, n45871, n31739, n906, n31452, n31451, 
        n18523, n31450, n2786, n2819, n31738, n2787, n31737, n15788, 
        n31449, n2788, n31736, n2789, n31735, n2790, n31734, n2791, 
        n31733, n2792, n31732, n2793, n31731, n2794, n31730, n2795, 
        n31729, \neo_pixel_transmitter.done_N_576 , n18367, n2796, n31728, 
        n2797, n31727, n31174, n31173, n31172, n2798, n31726, 
        n2799, n31725, n31171, n2800, n31724, n31170, n2801, n31723, 
        n31169, n2802, n31722, n31168, n2803, n31721, n31167, 
        n2804, n31720, n31166, n30285, n31165, n2805, n31719, 
        n2806, n31718, n31164, n31159, n2807, n31717, n2808, n31716, 
        n30432, n30431, n30430, n2809, n45875, n31715, n30265, 
        n30284, n30429, n2687, n2720, n31714, n2688, n31713, n2689, 
        n31712, n30428, n31711, n42, n31710, n30427, n46, n44, 
        n30283, n45, n43, n30426, n31709, n31708, n31707, n40_adj_4246, 
        n48, n52, n31706, n39_adj_4247, n31705, n31704, n30425, 
        n31703, n31702, n31701, n31700, n30282, n31699, n30281, 
        n30424, n30280, n31698, n31697, n30279, n31696, n31160, 
        n31161, n31695, n31694, n31162, n30423, n30422, n39589, 
        n31163, n30278, n30421, n30277, n31693, n30420, n45876, 
        n31692, n31691, n31690, n24_adj_4251, n22_adj_4252, n23_adj_4253, 
        n21_adj_4254, n4_adj_4255, n38076, n39504, n39505, n26_adj_4256, 
        n19_adj_4257, n16_adj_4258, n24_adj_4259, n28_adj_4260, n28_adj_4261, 
        n32_adj_4262, n30_adj_4263, n31_adj_4264, n30_adj_4265, n33679, 
        n29_adj_4266, n7476, n38194, n17_adj_4267, n29_adj_4268, n37_adj_4269, 
        n36_adj_4270, n42_adj_4271, n40_adj_4272, n41, n39_adj_4273, 
        n38174, n103, n37231, n40_adj_4274, n38_adj_4275, n39_adj_4276, 
        n37_adj_4277, n34_adj_4278, n42_adj_4279, n46_adj_4280, n33_adj_4281, 
        n33784, n8_adj_4282, n40825, n6_adj_4283, n27353, n12_adj_4284, 
        n14_adj_4285, n9_adj_4286, n33_adj_4287, n41_adj_4288, n38_adj_4289, 
        n43_adj_4290, n40_adj_4291, n46_adj_4292, n39_adj_4293, n47, 
        n19_adj_4294, n32958, n10_adj_4295, n12_adj_4296, n16_adj_4297, 
        n18_adj_4298, n18_adj_4299, n27289, n16_adj_4300, n17_adj_4301, 
        n44_adj_4302, n33_adj_4303, n40_adj_4304, n45_adj_4305, n42_adj_4306, 
        n48_adj_4307, n41_adj_4308, n49, n18_adj_4309, n20_adj_4310, 
        n15_adj_4311, n27379, n48_adj_4312, n46_adj_4313, n47_adj_4314, 
        n45_adj_4315, n44_adj_4316, n43_adj_4317, n54, n49_adj_4318, 
        n27449, n19_adj_4319, n42814, n25_adj_4320, n7_adj_4321, n20_adj_4322, 
        n13_adj_4323, n18_adj_4324, n22_adj_4325, n807;
    
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n31688), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_19 (.CI(n30418), .I0(timer[17]), .I1(n1[17]), 
            .CO(n30419));
    SB_LUT4 timer_1147_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n31157), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_21 (.CI(n31688), .I0(n2591), .I1(n2621), .CO(n31689));
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk32MHz), .E(n39942), .D(\neo_pixel_transmitter.done_N_570 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n31687), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_18_lut (.I0(one_wire_N_513[29]), .I1(timer[16]), 
            .I2(n1[16]), .I3(n30417), .O(n24)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1808_20 (.CI(n31687), .I0(n2592), .I1(n2621), .CO(n31688));
    SB_CARRY sub_14_add_2_18 (.CI(n30417), .I0(timer[16]), .I1(n1[16]), 
            .CO(n30418));
    SB_CARRY timer_1147_add_4_16 (.CI(n31157), .I0(GND_net), .I1(timer[14]), 
            .CO(n31158));
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n31686), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_19 (.CI(n31686), .I0(n2593), .I1(n2621), .CO(n31687));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n31685), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_18 (.CI(n31685), .I0(n2594), .I1(n2621), .CO(n31686));
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n31684), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_17 (.CI(n31684), .I0(n2595), .I1(n2621), .CO(n31685));
    SB_LUT4 timer_1147_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n31156), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1147_add_4_15 (.CI(n31156), .I0(GND_net), .I1(timer[13]), 
            .CO(n31157));
    SB_LUT4 add_21_19_lut (.I0(n19), .I1(bit_ctr[17]), .I2(GND_net), .I3(n30275), 
            .O(n42947)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n31683), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_16 (.CI(n31683), .I0(n2596), .I1(n2621), .CO(n31684));
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n31682), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1147_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n31155), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1147_add_4_14 (.CI(n31155), .I0(GND_net), .I1(timer[12]), 
            .CO(n31156));
    SB_LUT4 sub_14_add_2_17_lut (.I0(one_wire_N_513[20]), .I1(timer[15]), 
            .I2(n1[15]), .I3(n30416), .O(n6)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 timer_1147_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n31154), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_7_lut (.I0(n19), .I1(bit_ctr[5]), .I2(GND_net), .I3(n30263), 
            .O(n42956)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_14_add_2_17 (.CI(n30416), .I0(timer[15]), .I1(n1[15]), 
            .CO(n30417));
    SB_LUT4 sub_14_add_2_16_lut (.I0(one_wire_N_513[24]), .I1(timer[14]), 
            .I2(n1[14]), .I3(n30415), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1808_15 (.CI(n31682), .I0(n2597), .I1(n2621), .CO(n31683));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n31681), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_16 (.CI(n30415), .I0(timer[14]), .I1(n1[14]), 
            .CO(n30416));
    SB_CARRY mod_5_add_1808_14 (.CI(n31681), .I0(n2598), .I1(n2621), .CO(n31682));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n31680), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_13 (.CI(n31680), .I0(n2599), .I1(n2621), .CO(n31681));
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n31679), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_12 (.CI(n31679), .I0(n2600), .I1(n2621), .CO(n31680));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n31678), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_11 (.CI(n31678), .I0(n2601), .I1(n2621), .CO(n31679));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n31677), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_10 (.CI(n31677), .I0(n2602), .I1(n2621), .CO(n31678));
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n31676), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1147_add_4_13 (.CI(n31154), .I0(GND_net), .I1(timer[11]), 
            .CO(n31155));
    SB_CARRY mod_5_add_1808_9 (.CI(n31676), .I0(n2603), .I1(n2621), .CO(n31677));
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n31675), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_8 (.CI(n31675), .I0(n2604), .I1(n2621), .CO(n31676));
    SB_LUT4 sub_14_add_2_15_lut (.I0(one_wire_N_513[19]), .I1(timer[13]), 
            .I2(n1[13]), .I3(n30414), .O(n20)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n31674), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1147_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n31153), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_7 (.CI(n31674), .I0(n2605), .I1(n2621), .CO(n31675));
    SB_DFF bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(clk32MHz), .D(n35971));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(clk32MHz), .D(n35973));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(clk32MHz), .D(n35975));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(clk32MHz), .D(n35967));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(clk32MHz), .D(n35969));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(clk32MHz), .D(n35963));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(clk32MHz), .D(n35965));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(clk32MHz), .D(n35959));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(clk32MHz), .D(n35961));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(clk32MHz), .D(n35955));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(clk32MHz), .D(n35957));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(clk32MHz), .D(n35951));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(clk32MHz), .D(n35953));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(clk32MHz), .D(n35947));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(clk32MHz), .D(n35949));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(clk32MHz), .D(n35933));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(clk32MHz), .D(n35935));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(clk32MHz), .D(n35937));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(clk32MHz), .D(n35939));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(clk32MHz), .D(n35941));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(clk32MHz), .D(n35943));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(clk32MHz), .D(n35931));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(clk32MHz), .D(n35925));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(clk32MHz), .E(VCC_net), 
            .D(n35907));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(clk32MHz), .D(n35927));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(clk32MHz), .E(VCC_net), 
            .D(n35909));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(clk32MHz), .E(VCC_net), 
            .D(n35911));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(clk32MHz), .D(n35929));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY timer_1147_add_4_12 (.CI(n31153), .I0(GND_net), .I1(timer[10]), 
            .CO(n31154));
    SB_LUT4 timer_1147_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n31152), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1147_add_4_11 (.CI(n31152), .I0(GND_net), .I1(timer[9]), 
            .CO(n31153));
    SB_LUT4 timer_1147_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n31151), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1147_add_4_10 (.CI(n31151), .I0(GND_net), .I1(timer[8]), 
            .CO(n31152));
    SB_LUT4 timer_1147_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n31150), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i11_4_lut (.I0(n2302), .I1(n2292), .I2(n2293), .I3(n2301), 
            .O(n30));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22211_2_lut (.I0(bit_ctr[12]), .I1(n2309), .I2(GND_net), 
            .I3(GND_net), .O(n27219));
    defparam i22211_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15_4_lut (.I0(n2294), .I1(n30), .I2(n2306), .I3(n2304), 
            .O(n34));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut (.I0(n2291), .I1(n2303), .I2(n27219), .I3(n2305), 
            .O(n32));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY timer_1147_add_4_9 (.CI(n31150), .I0(GND_net), .I1(timer[7]), 
            .CO(n31151));
    SB_LUT4 i14_4_lut (.I0(n2298), .I1(n2295), .I2(n2296), .I3(n2300), 
            .O(n33));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n2308), .I1(n2297), .I2(n2307), .I3(n2299), 
            .O(n31));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut (.I0(n31), .I1(n33), .I2(n32), .I3(n34), .O(n2324));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 timer_1147_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n31149), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1147_add_4_8 (.CI(n31149), .I0(GND_net), .I1(timer[6]), 
            .CO(n31150));
    SB_LUT4 timer_1147_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n31148), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1147_add_4_7 (.CI(n31148), .I0(GND_net), .I1(timer[5]), 
            .CO(n31149));
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i38732_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45855));
    defparam i38732_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_14_add_2_15 (.CI(n30414), .I0(timer[13]), .I1(n1[13]), 
            .CO(n30415));
    SB_LUT4 timer_1147_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n31147), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n31673), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_3_lut (.I0(bit_ctr[11]), .I1(n2403), .I2(n2409), .I3(GND_net), 
            .O(n27));
    defparam i7_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut_adj_1480 (.I0(n2390), .I1(n2391), .I2(n2397), .I3(n2394), 
            .O(n33_adj_4196));
    defparam i13_4_lut_adj_1480.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1481 (.I0(n2392), .I1(n2405), .I2(n2400), .I3(n2398), 
            .O(n32_adj_4197));
    defparam i12_4_lut_adj_1481.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1482 (.I0(n2396), .I1(n2402), .I2(n2408), .I3(n2399), 
            .O(n31_adj_4198));
    defparam i11_4_lut_adj_1482.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1483 (.I0(n2393), .I1(n2406), .I2(n2395), .I3(n2407), 
            .O(n35));
    defparam i15_4_lut_adj_1483.LUT_INIT = 16'hfffe;
    SB_CARRY timer_1147_add_4_6 (.CI(n31147), .I0(GND_net), .I1(timer[4]), 
            .CO(n31148));
    SB_LUT4 i17_4_lut (.I0(n33_adj_4196), .I1(n27), .I2(n2404), .I3(n2401), 
            .O(n37));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n37), .I1(n35), .I2(n31_adj_4198), .I3(n32_adj_4197), 
            .O(n2423));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_1147_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n31146), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1147_add_4_5 (.CI(n31146), .I0(GND_net), .I1(timer[3]), 
            .CO(n31147));
    SB_LUT4 timer_1147_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n31145), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1147_add_4_4 (.CI(n31145), .I0(GND_net), .I1(timer[2]), 
            .CO(n31146));
    SB_LUT4 timer_1147_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n31144), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i38731_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45854));
    defparam i38731_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_1147_add_4_3 (.CI(n31144), .I0(GND_net), .I1(timer[1]), 
            .CO(n31145));
    SB_LUT4 timer_1147_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1147_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n31144));
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1808_6 (.CI(n31673), .I0(n2606), .I1(n2621), .CO(n31674));
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_add_2_14_lut (.I0(n18_adj_4200), .I1(timer[12]), .I2(n1[12]), 
            .I3(n30413), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n31672), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_14 (.CI(n30413), .I0(timer[12]), .I1(n1[12]), 
            .CO(n30414));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n30412), .O(\one_wire_N_513[11] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_14_add_2_13 (.CI(n30412), .I0(timer[11]), .I1(n1[11]), 
            .CO(n30413));
    SB_CARRY add_21_19 (.CI(n30275), .I0(bit_ctr[17]), .I1(GND_net), .CO(n30276));
    SB_CARRY mod_5_add_1808_5 (.CI(n31672), .I0(n2607), .I1(n2621), .CO(n31673));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n31671), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_4 (.CI(n31671), .I0(n2608), .I1(n2621), .CO(n31672));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n30411), .O(one_wire_N_513[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n45853), 
            .I3(n31670), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_3 (.CI(n31670), .I0(n2609), .I1(n45853), .CO(n31671));
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n45853), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n45853), 
            .CO(n31670));
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n31669), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_12 (.CI(n30411), .I0(timer[10]), .I1(n1[10]), 
            .CO(n30412));
    SB_LUT4 add_21_18_lut (.I0(n19), .I1(bit_ctr[16]), .I2(GND_net), .I3(n30274), 
            .O(n42943)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n31668), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_22 (.CI(n31668), .I0(n2490), .I1(n2522), .CO(n31669));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n31667), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n30410), .O(one_wire_N_513[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_21 (.CI(n31667), .I0(n2491), .I1(n2522), .CO(n31668));
    SB_LUT4 mod_5_add_1741_20_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n31666), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_11 (.CI(n30410), .I0(timer[9]), .I1(n1[9]), 
            .CO(n30411));
    SB_LUT4 sub_14_add_2_10_lut (.I0(one_wire_N_513[10]), .I1(timer[8]), 
            .I2(n1[8]), .I3(n30409), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i12_3_lut_4_lut_3_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(bit_ctr[29]), 
            .I3(GND_net), .O(n708));   // verilog/neopixel.v(22[26:36])
    defparam i12_3_lut_4_lut_3_lut.LUT_INIT = 16'h4242;
    SB_CARRY sub_14_add_2_10 (.CI(n30409), .I0(timer[8]), .I1(n1[8]), 
            .CO(n30410));
    SB_CARRY mod_5_add_1741_20 (.CI(n31666), .I0(n2492), .I1(n2522), .CO(n31667));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n31665), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_19 (.CI(n31665), .I0(n2493), .I1(n2522), .CO(n31666));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n31664), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_18 (.CI(n31664), .I0(n2494), .I1(n2522), .CO(n31665));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n31663), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_17 (.CI(n31663), .I0(n2495), .I1(n2522), .CO(n31664));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n31662), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_16 (.CI(n31662), .I0(n2496), .I1(n2522), .CO(n31663));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n31661), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_18 (.CI(n30274), .I0(bit_ctr[16]), .I1(GND_net), .CO(n30275));
    SB_CARRY mod_5_add_1741_15 (.CI(n31661), .I0(n2497), .I1(n2522), .CO(n31662));
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1741_14_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n31660), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_7 (.CI(n30263), .I0(bit_ctr[5]), .I1(GND_net), .CO(n30264));
    SB_LUT4 add_21_17_lut (.I0(n19), .I1(bit_ctr[15]), .I2(GND_net), .I3(n30273), 
            .O(n42966)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3718_2_lut_3_lut (.I0(n15780), .I1(bit_ctr[27]), .I2(n38037), 
            .I3(GND_net), .O(n60));   // verilog/neopixel.v(22[26:36])
    defparam i3718_2_lut_3_lut.LUT_INIT = 16'hf4f4;
    SB_CARRY mod_5_add_1741_14 (.CI(n31660), .I0(n2498), .I1(n2522), .CO(n31661));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n31659), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_13 (.CI(n31659), .I0(n2499), .I1(n2522), .CO(n31660));
    SB_LUT4 i22229_2_lut (.I0(bit_ctr[15]), .I1(n2009), .I2(GND_net), 
            .I3(GND_net), .O(n27237));
    defparam i22229_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38006_3_lut_4_lut (.I0(n15780), .I1(bit_ctr[27]), .I2(n838), 
            .I3(n38037), .O(n38039));   // verilog/neopixel.v(22[26:36])
    defparam i38006_3_lut_4_lut.LUT_INIT = 16'hf40b;
    SB_LUT4 i12_4_lut_adj_1484 (.I0(n2000), .I1(n1999), .I2(n2007), .I3(n2003), 
            .O(n28_adj_4203));
    defparam i12_4_lut_adj_1484.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1741_12_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n31658), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_12 (.CI(n31658), .I0(n2500), .I1(n2522), .CO(n31659));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n31657), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n30408), .O(\one_wire_N_513[7] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_9 (.CI(n30408), .I0(timer[7]), .I1(n1[7]), .CO(n30409));
    SB_CARRY mod_5_add_1741_11 (.CI(n31657), .I0(n2501), .I1(n2522), .CO(n31658));
    SB_LUT4 i10_4_lut (.I0(n1996), .I1(n1994), .I2(n2006), .I3(n27237), 
            .O(n26_adj_4204));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1485 (.I0(n1997), .I1(n2001), .I2(n1995), .I3(n2008), 
            .O(n27_adj_4205));
    defparam i11_4_lut_adj_1485.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1741_10_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n31656), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i9_4_lut (.I0(n2004), .I1(n2002), .I2(n2005), .I3(n1998), 
            .O(n25_adj_4206));
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1486 (.I0(n25_adj_4206), .I1(n27_adj_4205), .I2(n26_adj_4204), 
            .I3(n28_adj_4203), .O(n2027));
    defparam i15_4_lut_adj_1486.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1741_10 (.CI(n31656), .I0(n2502), .I1(n2522), .CO(n31657));
    SB_LUT4 mod_5_add_1741_9_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n31655), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_9 (.CI(n31655), .I0(n2503), .I1(n2522), .CO(n31656));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n31654), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_8_lut (.I0(one_wire_N_513[9]), .I1(timer[6]), .I2(n1[6]), 
            .I3(n30407), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_8 (.CI(n30407), .I0(timer[6]), .I1(n1[6]), .CO(n30408));
    SB_LUT4 add_21_6_lut (.I0(n19), .I1(bit_ctr[4]), .I2(GND_net), .I3(n30262), 
            .O(n42955)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_17 (.CI(n30273), .I0(bit_ctr[15]), .I1(GND_net), .CO(n30274));
    SB_CARRY mod_5_add_1741_8 (.CI(n31654), .I0(n2504), .I1(n2522), .CO(n31655));
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n30406), .O(\one_wire_N_513[5] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_7_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n31653), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1741_7 (.CI(n31653), .I0(n2505), .I1(n2522), .CO(n31654));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n31652), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_6 (.CI(n31652), .I0(n2506), .I1(n2522), .CO(n31653));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n31651), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_5 (.CI(n31651), .I0(n2507), .I1(n2522), .CO(n31652));
    SB_LUT4 mod_5_add_1741_4_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n31650), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_16_lut (.I0(n19), .I1(bit_ctr[14]), .I2(GND_net), .I3(n30272), 
            .O(n42965)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1741_4 (.CI(n31650), .I0(n2508), .I1(n2522), .CO(n31651));
    SB_LUT4 mod_5_add_1741_3_lut (.I0(n2509), .I1(n2509), .I2(n45854), 
            .I3(n31649), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY sub_14_add_2_7 (.CI(n30406), .I0(timer[5]), .I1(n1[5]), .CO(n30407));
    SB_CARRY mod_5_add_1741_3 (.CI(n31649), .I0(n2509), .I1(n45854), .CO(n31650));
    SB_LUT4 mod_5_add_1741_2_lut (.I0(bit_ctr[10]), .I1(bit_ctr[10]), .I2(n45854), 
            .I3(VCC_net), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n30405), .O(one_wire_N_513[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(n45854), 
            .CO(n31649));
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n31648), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n31647), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_21 (.CI(n31647), .I0(n2391), .I1(n2423), .CO(n31648));
    SB_LUT4 i38735_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45858));
    defparam i38735_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1674_20_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n31646), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_20 (.CI(n31646), .I0(n2392), .I1(n2423), .CO(n31647));
    SB_LUT4 mod_5_add_1674_19_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n31645), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_19 (.CI(n31645), .I0(n2393), .I1(n2423), .CO(n31646));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n31644), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_18 (.CI(n31644), .I0(n2394), .I1(n2423), .CO(n31645));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n31643), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_17 (.CI(n31643), .I0(n2395), .I1(n2423), .CO(n31644));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n31642), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_6 (.CI(n30405), .I0(timer[4]), .I1(n1[4]), .CO(n30406));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n30404), .O(one_wire_N_513[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_16 (.CI(n31642), .I0(n2396), .I1(n2423), .CO(n31643));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n31641), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_15 (.CI(n31641), .I0(n2397), .I1(n2423), .CO(n31642));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n31640), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_14 (.CI(n31640), .I0(n2398), .I1(n2423), .CO(n31641));
    SB_LUT4 mod_5_add_1674_13_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n31639), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_13 (.CI(n31639), .I0(n2399), .I1(n2423), .CO(n31640));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n31638), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_12 (.CI(n31638), .I0(n2400), .I1(n2423), .CO(n31639));
    SB_LUT4 mod_5_add_1674_11_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n31637), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_11 (.CI(n31637), .I0(n2401), .I1(n2423), .CO(n31638));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n31636), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_10 (.CI(n31636), .I0(n2402), .I1(n2423), .CO(n31637));
    SB_CARRY sub_14_add_2_5 (.CI(n30404), .I0(timer[3]), .I1(n1[3]), .CO(n30405));
    SB_LUT4 mod_5_add_1674_9_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n31635), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n30403), .O(one_wire_N_513[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_9 (.CI(n31635), .I0(n2403), .I1(n2423), .CO(n31636));
    SB_CARRY sub_14_add_2_4 (.CI(n30403), .I0(timer[2]), .I1(n1[2]), .CO(n30404));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n31634), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_8 (.CI(n31634), .I0(n2404), .I1(n2423), .CO(n31635));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n31633), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_7 (.CI(n31633), .I0(n2405), .I1(n2423), .CO(n31634));
    SB_LUT4 mod_5_add_1674_6_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n31632), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_6 (.CI(n31632), .I0(n2406), .I1(n2423), .CO(n31633));
    SB_LUT4 mod_5_add_1674_5_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n31631), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_5 (.CI(n31631), .I0(n2407), .I1(n2423), .CO(n31632));
    SB_LUT4 mod_5_add_1674_4_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n31630), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_4 (.CI(n31630), .I0(n2408), .I1(n2423), .CO(n31631));
    SB_LUT4 mod_5_add_1674_3_lut (.I0(n2409), .I1(n2409), .I2(n45855), 
            .I3(n31629), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_3 (.CI(n31629), .I0(n2409), .I1(n45855), .CO(n31630));
    SB_LUT4 sub_14_add_2_3_lut (.I0(n4), .I1(timer[1]), .I2(n1[1]), .I3(n30402), 
            .O(n32659)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1674_2_lut (.I0(bit_ctr[11]), .I1(bit_ctr[11]), .I2(n45855), 
            .I3(VCC_net), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(n45855), 
            .CO(n31629));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n31628), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n31627), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_20 (.CI(n31627), .I0(n2292), .I1(n2324), .CO(n31628));
    SB_LUT4 mod_5_add_1607_19_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n31626), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_19 (.CI(n31626), .I0(n2293), .I1(n2324), .CO(n31627));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n31625), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_18 (.CI(n31625), .I0(n2294), .I1(n2324), .CO(n31626));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n31624), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_17 (.CI(n31624), .I0(n2295), .I1(n2324), .CO(n31625));
    SB_LUT4 mod_5_add_1607_16_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n31623), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_3 (.CI(n30402), .I0(timer[1]), .I1(n1[1]), .CO(n30403));
    SB_CARRY mod_5_add_1607_16 (.CI(n31623), .I0(n2296), .I1(n2324), .CO(n31624));
    SB_LUT4 mod_5_add_1607_15_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n31622), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_15 (.CI(n31622), .I0(n2297), .I1(n2324), .CO(n31623));
    SB_LUT4 mod_5_add_1607_14_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n31621), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_14 (.CI(n31621), .I0(n2298), .I1(n2324), .CO(n31622));
    SB_LUT4 mod_5_add_1607_13_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n31620), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_16 (.CI(n30272), .I0(bit_ctr[14]), .I1(GND_net), .CO(n30273));
    SB_CARRY mod_5_add_1607_13 (.CI(n31620), .I0(n2299), .I1(n2324), .CO(n31621));
    SB_LUT4 mod_5_add_1607_12_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n31619), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_12 (.CI(n31619), .I0(n2300), .I1(n2324), .CO(n31620));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n31618), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_11 (.CI(n31618), .I0(n2301), .I1(n2324), .CO(n31619));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n31617), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_10 (.CI(n31617), .I0(n2302), .I1(n2324), .CO(n31618));
    SB_CARRY add_21_6 (.CI(n30262), .I0(bit_ctr[4]), .I1(GND_net), .CO(n30263));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n31616), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_2_lut (.I0(one_wire_N_513[2]), .I1(timer[0]), .I2(n1[0]), 
            .I3(VCC_net), .O(n4)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1607_9 (.CI(n31616), .I0(n2303), .I1(n2324), .CO(n31617));
    SB_LUT4 add_21_15_lut (.I0(n19), .I1(bit_ctr[13]), .I2(GND_net), .I3(n30271), 
            .O(n42964)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n30402));
    SB_LUT4 mod_5_add_1607_8_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n31615), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_8 (.CI(n31615), .I0(n2304), .I1(n2324), .CO(n31616));
    SB_LUT4 mod_5_add_1607_7_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n31614), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_7 (.CI(n31614), .I0(n2305), .I1(n2324), .CO(n31615));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n31613), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_6 (.CI(n31613), .I0(n2306), .I1(n2324), .CO(n31614));
    SB_LUT4 mod_5_add_1607_5_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n31612), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_5 (.CI(n31612), .I0(n2307), .I1(n2324), .CO(n31613));
    SB_LUT4 mod_5_add_1607_4_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n31611), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_4 (.CI(n31611), .I0(n2308), .I1(n2324), .CO(n31612));
    SB_LUT4 mod_5_add_1607_3_lut (.I0(n2309), .I1(n2309), .I2(n45856), 
            .I3(n31610), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_3 (.CI(n31610), .I0(n2309), .I1(n45856), .CO(n31611));
    SB_LUT4 mod_5_add_1607_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[12]), .I2(n45856), 
            .I3(VCC_net), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(n45856), 
            .CO(n31610));
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n31609), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_19_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n31608), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_19 (.CI(n31608), .I0(n2193), .I1(n2225), .CO(n31609));
    SB_LUT4 mod_5_add_1540_18_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n31607), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_18 (.CI(n31607), .I0(n2194), .I1(n2225), .CO(n31608));
    SB_LUT4 mod_5_add_1540_17_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n31606), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_17 (.CI(n31606), .I0(n2195), .I1(n2225), .CO(n31607));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n31605), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_16 (.CI(n31605), .I0(n2196), .I1(n2225), .CO(n31606));
    SB_LUT4 mod_5_add_1540_15_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n31604), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1540_15 (.CI(n31604), .I0(n2197), .I1(n2225), .CO(n31605));
    SB_LUT4 mod_5_add_1540_14_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n31603), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_14 (.CI(n31603), .I0(n2198), .I1(n2225), .CO(n31604));
    SB_LUT4 mod_5_add_1540_13_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n31602), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_13 (.CI(n31602), .I0(n2199), .I1(n2225), .CO(n31603));
    SB_LUT4 mod_5_add_1540_12_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n31601), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_12 (.CI(n31601), .I0(n2200), .I1(n2225), .CO(n31602));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n31600), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_2_lut (.I0(n2491), .I1(n2504), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_4208));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_1487 (.I0(n2496), .I1(n2505), .I2(n2500), .I3(n2499), 
            .O(n34_adj_4209));
    defparam i13_4_lut_adj_1487.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[10]), .I1(n2497), .I2(n2509), .I3(GND_net), 
            .O(n22_adj_4210));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i17_4_lut_adj_1488 (.I0(n2490), .I1(n34_adj_4209), .I2(n24_adj_4208), 
            .I3(n2494), .O(n38));
    defparam i17_4_lut_adj_1488.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_5_lut (.I0(n19), .I1(bit_ctr[3]), .I2(GND_net), .I3(n30261), 
            .O(n42954)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1540_11 (.CI(n31600), .I0(n2201), .I1(n2225), .CO(n31601));
    SB_LUT4 i15_4_lut_adj_1489 (.I0(n2501), .I1(n2502), .I2(n2506), .I3(n2492), 
            .O(n36));
    defparam i15_4_lut_adj_1489.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_10_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n31599), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_10 (.CI(n31599), .I0(n2202), .I1(n2225), .CO(n31600));
    SB_LUT4 mod_5_add_1540_9_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n31598), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_9 (.CI(n31598), .I0(n2203), .I1(n2225), .CO(n31599));
    SB_LUT4 i16_4_lut (.I0(n2495), .I1(n2498), .I2(n2493), .I3(n22_adj_4210), 
            .O(n37_adj_4211));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_8_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n31597), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i14_4_lut_adj_1490 (.I0(n2507), .I1(n2508), .I2(n2503), .I3(n2489), 
            .O(n35_adj_4212));
    defparam i14_4_lut_adj_1490.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1540_8 (.CI(n31597), .I0(n2204), .I1(n2225), .CO(n31598));
    SB_LUT4 i20_4_lut (.I0(n35_adj_4212), .I1(n37_adj_4211), .I2(n36), 
            .I3(n38), .O(n2522));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut (.I0(n27335), .I1(n17206), .I2(n38094), .I3(\state[1] ), 
            .O(n38456));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 mod_5_add_1540_7_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n31596), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_7 (.CI(n31596), .I0(n2205), .I1(n2225), .CO(n31597));
    SB_CARRY add_21_15 (.CI(n30271), .I0(bit_ctr[13]), .I1(GND_net), .CO(n30272));
    SB_LUT4 mod_5_add_1540_6_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n31595), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i38730_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45853));
    defparam i38730_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1540_6 (.CI(n31595), .I0(n2206), .I1(n2225), .CO(n31596));
    SB_LUT4 mod_5_add_1540_5_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n31594), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_5 (.CI(n31594), .I0(n2207), .I1(n2225), .CO(n31595));
    SB_LUT4 add_21_14_lut (.I0(n19), .I1(bit_ctr[12]), .I2(GND_net), .I3(n30270), 
            .O(n42963)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1540_4_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n31593), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_4 (.CI(n31593), .I0(n2208), .I1(n2225), .CO(n31594));
    SB_LUT4 mod_5_add_1540_3_lut (.I0(n2209), .I1(n2209), .I2(n45857), 
            .I3(n31592), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1540_3 (.CI(n31592), .I0(n2209), .I1(n45857), .CO(n31593));
    SB_LUT4 mod_5_add_1540_2_lut (.I0(bit_ctr[13]), .I1(bit_ctr[13]), .I2(n45857), 
            .I3(VCC_net), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(n45857), 
            .CO(n31592));
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n31591), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_18_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n31590), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i36355_3_lut_4_lut (.I0(n27335), .I1(n17206), .I2(start), 
            .I3(n38094), .O(n42968));
    defparam i36355_3_lut_4_lut.LUT_INIT = 16'hf0fe;
    SB_LUT4 i224_2_lut_3_lut (.I0(n27335), .I1(n17206), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n1108));
    defparam i224_2_lut_3_lut.LUT_INIT = 16'hf1f1;
    SB_CARRY mod_5_add_1473_18 (.CI(n31590), .I0(n2094), .I1(n2126), .CO(n31591));
    SB_CARRY add_21_14 (.CI(n30270), .I0(bit_ctr[12]), .I1(GND_net), .CO(n30271));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n31589), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_17 (.CI(n31589), .I0(n2095), .I1(n2126), .CO(n31590));
    SB_LUT4 mod_5_add_1473_16_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n31588), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_16 (.CI(n31588), .I0(n2096), .I1(n2126), .CO(n31589));
    SB_LUT4 mod_5_add_1473_15_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n31587), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_15 (.CI(n31587), .I0(n2097), .I1(n2126), .CO(n31588));
    SB_LUT4 mod_5_add_1473_14_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n31586), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_14 (.CI(n31586), .I0(n2098), .I1(n2126), .CO(n31587));
    SB_LUT4 mod_5_add_1473_13_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n31585), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_13 (.CI(n31585), .I0(n2099), .I1(n2126), .CO(n31586));
    SB_LUT4 mod_5_add_1473_12_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n31584), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_12 (.CI(n31584), .I0(n2100), .I1(n2126), .CO(n31585));
    SB_LUT4 mod_5_add_1473_11_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n31583), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_13_lut (.I0(n19), .I1(bit_ctr[11]), .I2(GND_net), .I3(n30269), 
            .O(n42962)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1473_11 (.CI(n31583), .I0(n2101), .I1(n2126), .CO(n31584));
    SB_LUT4 mod_5_add_1473_10_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n31582), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_10 (.CI(n31582), .I0(n2102), .I1(n2126), .CO(n31583));
    SB_LUT4 mod_5_add_1473_9_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n31581), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_DFF bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(clk32MHz), .D(n35923));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1473_9 (.CI(n31581), .I0(n2103), .I1(n2126), .CO(n31582));
    SB_LUT4 mod_5_add_1473_8_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n31580), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_8 (.CI(n31580), .I0(n2104), .I1(n2126), .CO(n31581));
    SB_LUT4 mod_5_add_1473_7_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n31579), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut_adj_1491 (.I0(bit_ctr[17]), .I1(bit_ctr[31]), .I2(bit_ctr[28]), 
            .I3(bit_ctr[12]), .O(n27_adj_4213));
    defparam i10_4_lut_adj_1491.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1473_7 (.CI(n31579), .I0(n2105), .I1(n2126), .CO(n31580));
    SB_CARRY add_21_13 (.CI(n30269), .I0(bit_ctr[11]), .I1(GND_net), .CO(n30270));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n31578), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_5 (.CI(n30261), .I0(bit_ctr[3]), .I1(GND_net), .CO(n30262));
    SB_LUT4 add_21_4_lut (.I0(n19), .I1(bit_ctr[2]), .I2(GND_net), .I3(n30260), 
            .O(n42953)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1473_6 (.CI(n31578), .I0(n2106), .I1(n2126), .CO(n31579));
    SB_LUT4 mod_5_add_1473_5_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n31577), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_5 (.CI(n31577), .I0(n2107), .I1(n2126), .CO(n31578));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n31576), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_12_lut (.I0(n19), .I1(bit_ctr[10]), .I2(GND_net), .I3(n30268), 
            .O(n42961)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1473_4 (.CI(n31576), .I0(n2108), .I1(n2126), .CO(n31577));
    SB_LUT4 mod_5_add_1473_3_lut (.I0(n2109), .I1(n2109), .I2(n45858), 
            .I3(n31575), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_3 (.CI(n31575), .I0(n2109), .I1(n45858), .CO(n31576));
    SB_LUT4 mod_5_add_1473_2_lut (.I0(bit_ctr[14]), .I1(bit_ctr[14]), .I2(n45858), 
            .I3(VCC_net), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(n45858), 
            .CO(n31575));
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n31574), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_12 (.CI(n30268), .I0(bit_ctr[10]), .I1(GND_net), .CO(n30269));
    SB_LUT4 mod_5_add_1406_17_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n31573), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_17 (.CI(n31573), .I0(n1995), .I1(n2027), .CO(n31574));
    SB_LUT4 mod_5_add_1406_16_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n31572), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_16 (.CI(n31572), .I0(n1996), .I1(n2027), .CO(n31573));
    SB_LUT4 mod_5_add_1406_15_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n31571), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_15 (.CI(n31571), .I0(n1997), .I1(n2027), .CO(n31572));
    SB_LUT4 mod_5_add_1406_14_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n31570), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_14 (.CI(n31570), .I0(n1998), .I1(n2027), .CO(n31571));
    SB_LUT4 mod_5_add_1406_13_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n31569), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_13 (.CI(n31569), .I0(n1999), .I1(n2027), .CO(n31570));
    SB_LUT4 mod_5_add_1406_12_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n31568), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_12 (.CI(n31568), .I0(n2000), .I1(n2027), .CO(n31569));
    SB_DFF timer_1147__i0 (.Q(timer[0]), .C(clk32MHz), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 mod_5_add_1406_11_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n31567), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i2007_3_lut (.I0(n17196), .I1(\state_3__N_362[1] ), .I2(\state[1] ), 
            .I3(GND_net), .O(n4724));
    defparam i2007_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i22156_2_lut (.I0(bit_ctr[3]), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(GND_net), .O(n27164));
    defparam i22156_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12_4_lut_adj_1492 (.I0(bit_ctr[5]), .I1(bit_ctr[16]), .I2(bit_ctr[14]), 
            .I3(bit_ctr[7]), .O(n29_adj_4214));
    defparam i12_4_lut_adj_1492.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1493 (.I0(bit_ctr[29]), .I1(bit_ctr[23]), .I2(bit_ctr[21]), 
            .I3(bit_ctr[20]), .O(n28_adj_4215));
    defparam i11_4_lut_adj_1493.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut (.I0(one_wire_N_513[3]), .I1(one_wire_N_513[4]), .I2(one_wire_N_513[2]), 
            .I3(GND_net), .O(n32476));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i22355_2_lut (.I0(n32476), .I1(n17064), .I2(GND_net), .I3(GND_net), 
            .O(n27365));
    defparam i22355_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut (.I0(n27172), .I1(one_wire_N_513[4]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4216));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1494 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n17195));   // verilog/neopixel.v(52[18] 72[12])
    defparam i1_2_lut_adj_1494.LUT_INIT = 16'hbbbb;
    SB_LUT4 i6_4_lut (.I0(\one_wire_N_513[5] ), .I1(\one_wire_N_513[11] ), 
            .I2(\one_wire_N_513[7] ), .I3(n17206), .O(n14));   // verilog/neopixel.v(104[14:39])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1495 (.I0(n8), .I1(n14), .I2(n10), .I3(GND_net), 
            .O(n17064));   // verilog/neopixel.v(104[14:39])
    defparam i7_3_lut_adj_1495.LUT_INIT = 16'hfefe;
    SB_LUT4 i31012_2_lut (.I0(\state[1] ), .I1(n17196), .I2(GND_net), 
            .I3(GND_net), .O(n38070));
    defparam i31012_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_1406_11 (.CI(n31567), .I0(n2001), .I1(n2027), .CO(n31568));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n31566), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_10 (.CI(n31566), .I0(n2002), .I1(n2027), .CO(n31567));
    SB_LUT4 mod_5_add_1406_9_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n31565), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i1_3_lut_adj_1496 (.I0(bit_ctr[14]), .I1(n2096), .I2(n2109), 
            .I3(GND_net), .O(n18_adj_4217));
    defparam i1_3_lut_adj_1496.LUT_INIT = 16'hecec;
    SB_CARRY mod_5_add_1406_9 (.CI(n31565), .I0(n2003), .I1(n2027), .CO(n31566));
    SB_LUT4 mod_5_add_1406_8_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n31564), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_8 (.CI(n31564), .I0(n2004), .I1(n2027), .CO(n31565));
    SB_LUT4 i13_4_lut_adj_1497 (.I0(n2105), .I1(n2107), .I2(n2094), .I3(n18_adj_4217), 
            .O(n30_adj_4218));
    defparam i13_4_lut_adj_1497.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1406_7_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n31563), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i11_4_lut_adj_1498 (.I0(n2106), .I1(n2097), .I2(n2102), .I3(n2093), 
            .O(n28_adj_4219));
    defparam i11_4_lut_adj_1498.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1499 (.I0(n2095), .I1(n2100), .I2(n2103), .I3(n2104), 
            .O(n29_adj_4220));
    defparam i12_4_lut_adj_1499.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1406_7 (.CI(n31563), .I0(n2005), .I1(n2027), .CO(n31564));
    SB_LUT4 mod_5_add_1406_6_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n31562), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_6 (.CI(n31562), .I0(n2006), .I1(n2027), .CO(n31563));
    SB_LUT4 i10_4_lut_adj_1500 (.I0(n2099), .I1(n2108), .I2(n2101), .I3(n2098), 
            .O(n27_adj_4221));
    defparam i10_4_lut_adj_1500.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1406_5_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n31561), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i16_4_lut_adj_1501 (.I0(n27_adj_4221), .I1(n29_adj_4220), .I2(n28_adj_4219), 
            .I3(n30_adj_4218), .O(n2126));
    defparam i16_4_lut_adj_1501.LUT_INIT = 16'hfffe;
    SB_LUT4 i38734_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45857));
    defparam i38734_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1406_5 (.CI(n31561), .I0(n2007), .I1(n2027), .CO(n31562));
    SB_LUT4 mod_5_add_1406_4_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n31560), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_4 (.CI(n31560), .I0(n2008), .I1(n2027), .CO(n31561));
    SB_LUT4 mod_5_add_1406_3_lut (.I0(n2009), .I1(n2009), .I2(n45859), 
            .I3(n31559), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1406_3 (.CI(n31559), .I0(n2009), .I1(n45859), .CO(n31560));
    SB_DFFE bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(clk32MHz), .E(VCC_net), 
            .D(n35913));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(clk32MHz), .D(n35917));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1406_2_lut (.I0(bit_ctr[15]), .I1(bit_ctr[15]), .I2(n45859), 
            .I3(VCC_net), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(n45859), 
            .CO(n31559));
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n31558), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_DFF bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(clk32MHz), .D(n35915));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk32MHz), .D(n18886));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1339_16_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n31557), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_16 (.CI(n31557), .I0(n1896), .I1(n1928), .CO(n31558));
    SB_LUT4 mod_5_add_1339_15_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n31556), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_15 (.CI(n31556), .I0(n1897), .I1(n1928), .CO(n31557));
    SB_LUT4 mod_5_add_1339_14_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n31555), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_14 (.CI(n31555), .I0(n1898), .I1(n1928), .CO(n31556));
    SB_LUT4 mod_5_add_1339_13_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n31554), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_13 (.CI(n31554), .I0(n1899), .I1(n1928), .CO(n31555));
    SB_LUT4 mod_5_add_1339_12_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n31553), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_12 (.CI(n31553), .I0(n1900), .I1(n1928), .CO(n31554));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n31552), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_11 (.CI(n31552), .I0(n1901), .I1(n1928), .CO(n31553));
    SB_LUT4 mod_5_add_1339_10_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n31551), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_10 (.CI(n31551), .I0(n1902), .I1(n1928), .CO(n31552));
    SB_LUT4 mod_5_add_1339_9_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n31550), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_9 (.CI(n31550), .I0(n1903), .I1(n1928), .CO(n31551));
    SB_LUT4 mod_5_add_1339_8_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n31549), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_8 (.CI(n31549), .I0(n1904), .I1(n1928), .CO(n31550));
    SB_LUT4 mod_5_add_1339_7_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n31548), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_7 (.CI(n31548), .I0(n1905), .I1(n1928), .CO(n31549));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n31547), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk32MHz), .D(n18885));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk32MHz), .D(n18884));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk32MHz), .D(n18883));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk32MHz), .D(n18882));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk32MHz), .D(n18881));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk32MHz), .D(n18880));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk32MHz), .D(n18879));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk32MHz), .D(n18878));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk32MHz), .D(n18877));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk32MHz), .D(n18876));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk32MHz), .D(n18875));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk32MHz), .D(n18874));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk32MHz), .D(n18873));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk32MHz), .D(n18872));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk32MHz), .D(n18871));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk32MHz), .D(n18870));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk32MHz), .D(n18869));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk32MHz), .D(n18868));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk32MHz), .D(n18867));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk32MHz), .D(n18866));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1339_6 (.CI(n31547), .I0(n1906), .I1(n1928), .CO(n31548));
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk32MHz), .D(n18865));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk32MHz), .D(n18864));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk32MHz), .D(n18863));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1339_5_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n31546), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_5 (.CI(n31546), .I0(n1907), .I1(n1928), .CO(n31547));
    SB_LUT4 mod_5_add_1339_4_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n31545), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_4 (.CI(n31545), .I0(n1908), .I1(n1928), .CO(n31546));
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk32MHz), .D(n18862));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk32MHz), .D(n18861));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk32MHz), .D(n18860));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk32MHz), .D(n18859));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk32MHz), .D(n18858));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk32MHz), .D(n18857));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk32MHz), .D(n18856));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk32MHz), .E(VCC_net), .D(n18855));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1339_3_lut (.I0(n1909), .I1(n1909), .I2(n45860), 
            .I3(n31544), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1339_3 (.CI(n31544), .I0(n1909), .I1(n45860), .CO(n31545));
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1502 (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n37332));
    defparam i1_2_lut_adj_1502.LUT_INIT = 16'h2222;
    SB_LUT4 i11_2_lut (.I0(n21_adj_4222), .I1(n22_adj_4223), .I2(GND_net), 
            .I3(GND_net), .O(n28_adj_4224));   // verilog/neopixel.v(104[14:39])
    defparam i11_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1503 (.I0(n23_adj_4225), .I1(n25_adj_4226), .I2(n24), 
            .I3(n26), .O(n32_adj_4227));   // verilog/neopixel.v(104[14:39])
    defparam i15_4_lut_adj_1503.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1504 (.I0(n19_adj_4228), .I1(n32_adj_4227), .I2(n28_adj_4224), 
            .I3(n20), .O(n17206));   // verilog/neopixel.v(104[14:39])
    defparam i16_4_lut_adj_1504.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1505 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4229));
    defparam i1_2_lut_adj_1505.LUT_INIT = 16'heeee;
    SB_LUT4 i31026_2_lut (.I0(one_wire_N_513[3]), .I1(one_wire_N_513[2]), 
            .I2(GND_net), .I3(GND_net), .O(n38086));
    defparam i31026_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22164_2_lut (.I0(n32659), .I1(one_wire_N_513[3]), .I2(GND_net), 
            .I3(GND_net), .O(n27172));
    defparam i22164_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(one_wire_N_513[4]), .I1(n37374), .I2(n27172), 
            .I3(n38086), .O(n116));
    defparam i1_4_lut.LUT_INIT = 16'h45cd;
    SB_LUT4 i38715_3_lut (.I0(n38192), .I1(n116), .I2(n17206), .I3(GND_net), 
            .O(n39942));
    defparam i38715_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_3_lut (.I0(n2600), .I1(bit_ctr[9]), .I2(n2609), .I3(GND_net), 
            .O(n26_adj_4230));
    defparam i4_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i14_4_lut_adj_1506 (.I0(n2601), .I1(n2604), .I2(n2593), .I3(n2596), 
            .O(n36_adj_4231));
    defparam i14_4_lut_adj_1506.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1507 (.I0(n2595), .I1(n2605), .I2(n2608), .I3(n2603), 
            .O(n34_adj_4232));
    defparam i12_4_lut_adj_1507.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1508 (.I0(n2590), .I1(n36_adj_4231), .I2(n26_adj_4230), 
            .I3(n2602), .O(n40));
    defparam i18_4_lut_adj_1508.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1509 (.I0(n2592), .I1(n2606), .I2(n2589), .I3(n2598), 
            .O(n38_adj_4233));
    defparam i16_4_lut_adj_1509.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2599), .I1(n34_adj_4232), .I2(n2588), .I3(GND_net), 
            .O(n39));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1510 (.I0(n2591), .I1(n2594), .I2(n2597), .I3(n2607), 
            .O(n37_adj_4234));
    defparam i15_4_lut_adj_1510.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(n37_adj_4234), .I1(n39), .I2(n38_adj_4233), 
            .I3(n40), .O(n2621));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1339_2_lut (.I0(bit_ctr[16]), .I1(bit_ctr[16]), .I2(n45860), 
            .I3(VCC_net), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(n45860), 
            .CO(n31544));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n31543), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n31542), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_15 (.CI(n31542), .I0(n1797), .I1(n1829), .CO(n31543));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n31541), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_14 (.CI(n31541), .I0(n1798), .I1(n1829), .CO(n31542));
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n31540), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_13 (.CI(n31540), .I0(n1799), .I1(n1829), .CO(n31541));
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n31539), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_12 (.CI(n31539), .I0(n1800), .I1(n1829), .CO(n31540));
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n31538), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_4 (.CI(n30260), .I0(bit_ctr[2]), .I1(GND_net), .CO(n30261));
    SB_CARRY mod_5_add_1272_11 (.CI(n31538), .I0(n1801), .I1(n1829), .CO(n31539));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n31537), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_10 (.CI(n31537), .I0(n1802), .I1(n1829), .CO(n31538));
    SB_LUT4 add_21_11_lut (.I0(n19), .I1(bit_ctr[9]), .I2(GND_net), .I3(n30267), 
            .O(n42960)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n31536), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_9 (.CI(n31536), .I0(n1803), .I1(n1829), .CO(n31537));
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n31535), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_8 (.CI(n31535), .I0(n1804), .I1(n1829), .CO(n31536));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n31534), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n31816), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_7 (.CI(n31534), .I0(n1805), .I1(n1829), .CO(n31535));
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n31533), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n31815), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_6 (.CI(n31533), .I0(n1806), .I1(n1829), .CO(n31534));
    SB_CARRY mod_5_add_2143_28 (.CI(n31815), .I0(n3084), .I1(n3116), .CO(n31816));
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n31532), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n31814), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_5 (.CI(n31532), .I0(n1807), .I1(n1829), .CO(n31533));
    SB_CARRY mod_5_add_2143_27 (.CI(n31814), .I0(n3085), .I1(n3116), .CO(n31815));
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n31531), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n31813), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_4 (.CI(n31531), .I0(n1808), .I1(n1829), .CO(n31532));
    SB_CARRY mod_5_add_2143_26 (.CI(n31813), .I0(n3086), .I1(n3116), .CO(n31814));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n45861), 
            .I3(n31530), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n31812), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_3 (.CI(n31530), .I0(n1809), .I1(n45861), .CO(n31531));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n45861), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_25 (.CI(n31812), .I0(n3087), .I1(n3116), .CO(n31813));
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n45861), 
            .CO(n31530));
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n31811), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n31529), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_24 (.CI(n31811), .I0(n3088), .I1(n3116), .CO(n31812));
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n31528), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n31810), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_23 (.CI(n31810), .I0(n3089), .I1(n3116), .CO(n31811));
    SB_CARRY mod_5_add_1205_14 (.CI(n31528), .I0(n1698), .I1(n1730), .CO(n31529));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n31527), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n31809), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_13 (.CI(n31527), .I0(n1699), .I1(n1730), .CO(n31528));
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n31526), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_22 (.CI(n31809), .I0(n3090), .I1(n3116), .CO(n31810));
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n31808), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_12 (.CI(n31526), .I0(n1700), .I1(n1730), .CO(n31527));
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n31525), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_21 (.CI(n31808), .I0(n3091), .I1(n3116), .CO(n31809));
    SB_CARRY mod_5_add_1205_11 (.CI(n31525), .I0(n1701), .I1(n1730), .CO(n31526));
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n31807), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n31524), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_20 (.CI(n31807), .I0(n3092), .I1(n3116), .CO(n31808));
    SB_CARRY mod_5_add_1205_10 (.CI(n31524), .I0(n1702), .I1(n1730), .CO(n31525));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n31806), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_19 (.CI(n31806), .I0(n3093), .I1(n3116), .CO(n31807));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n31523), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n31805), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_9 (.CI(n31523), .I0(n1703), .I1(n1730), .CO(n31524));
    SB_CARRY mod_5_add_2143_18 (.CI(n31805), .I0(n3094), .I1(n3116), .CO(n31806));
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n31522), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_8 (.CI(n31522), .I0(n1704), .I1(n1730), .CO(n31523));
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n31804), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_17 (.CI(n31804), .I0(n3095), .I1(n3116), .CO(n31805));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n31521), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_7 (.CI(n31521), .I0(n1705), .I1(n1730), .CO(n31522));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n31520), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n31803), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_6 (.CI(n31520), .I0(n1706), .I1(n1730), .CO(n31521));
    SB_CARRY mod_5_add_2143_16 (.CI(n31803), .I0(n3096), .I1(n3116), .CO(n31804));
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n31802), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n31519), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_15 (.CI(n31802), .I0(n3097), .I1(n3116), .CO(n31803));
    SB_CARRY mod_5_add_1205_5 (.CI(n31519), .I0(n1707), .I1(n1730), .CO(n31520));
    SB_LUT4 i9_4_lut_adj_1511 (.I0(n1707), .I1(n1702), .I2(n1697), .I3(n1703), 
            .O(n22_adj_4235));
    defparam i9_4_lut_adj_1511.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1512 (.I0(n1704), .I1(n1701), .I2(n1708), .I3(GND_net), 
            .O(n20_adj_4236));
    defparam i7_3_lut_adj_1512.LUT_INIT = 16'hfefe;
    SB_LUT4 i8_4_lut (.I0(n1698), .I1(n1700), .I2(n1705), .I3(n1706), 
            .O(n21_adj_4237));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_3_lut (.I0(n1699), .I1(bit_ctr[18]), .I2(n1709), .I3(GND_net), 
            .O(n19_adj_4238));
    defparam i6_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i12_4_lut_adj_1513 (.I0(n19_adj_4238), .I1(n21_adj_4237), .I2(n20_adj_4236), 
            .I3(n22_adj_4235), .O(n1730));
    defparam i12_4_lut_adj_1513.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n31801), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n31518), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_4 (.CI(n31518), .I0(n1708), .I1(n1730), .CO(n31519));
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n45864), 
            .I3(n31517), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_3 (.CI(n31517), .I0(n1709), .I1(n45864), .CO(n31518));
    SB_LUT4 add_21_3_lut (.I0(n19), .I1(bit_ctr[1]), .I2(GND_net), .I3(n30259), 
            .O(n42952)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_11 (.CI(n30267), .I0(bit_ctr[9]), .I1(GND_net), .CO(n30268));
    SB_CARRY mod_5_add_2143_14 (.CI(n31801), .I0(n3098), .I1(n3116), .CO(n31802));
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n45864), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n31800), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n45864), 
            .CO(n31517));
    SB_CARRY mod_5_add_2143_13 (.CI(n31800), .I0(n3099), .I1(n3116), .CO(n31801));
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n31516), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n31799), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n31515), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_12 (.CI(n31799), .I0(n3100), .I1(n3116), .CO(n31800));
    SB_CARRY mod_5_add_1138_13 (.CI(n31515), .I0(n1599), .I1(n1631), .CO(n31516));
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n31514), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n31798), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_12 (.CI(n31514), .I0(n1600), .I1(n1631), .CO(n31515));
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n31513), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_11 (.CI(n31798), .I0(n3101), .I1(n3116), .CO(n31799));
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n31797), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_11 (.CI(n31513), .I0(n1601), .I1(n1631), .CO(n31514));
    SB_CARRY mod_5_add_2143_10 (.CI(n31797), .I0(n3102), .I1(n3116), .CO(n31798));
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n31512), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n31796), .O(n3202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_10 (.CI(n31512), .I0(n1602), .I1(n1631), .CO(n31513));
    SB_CARRY mod_5_add_2143_9 (.CI(n31796), .I0(n3103), .I1(n3116), .CO(n31797));
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n31511), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n31795), .O(n3203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_9 (.CI(n31511), .I0(n1603), .I1(n1631), .CO(n31512));
    SB_CARRY mod_5_add_2143_8 (.CI(n31795), .I0(n3104), .I1(n3116), .CO(n31796));
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n31510), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n31794), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_8 (.CI(n31510), .I0(n1604), .I1(n1631), .CO(n31511));
    SB_CARRY mod_5_add_2143_7 (.CI(n31794), .I0(n3105), .I1(n3116), .CO(n31795));
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n31509), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_7 (.CI(n31509), .I0(n1605), .I1(n1631), .CO(n31510));
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(clk32MHz), .E(n18416), .D(state_3__N_362[0]), 
            .S(n18584));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n31508), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_3 (.CI(n30259), .I0(bit_ctr[1]), .I1(GND_net), .CO(n30260));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n31793), .O(n3205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_6 (.CI(n31508), .I0(n1606), .I1(n1631), .CO(n31509));
    SB_CARRY mod_5_add_2143_6 (.CI(n31793), .I0(n3106), .I1(n3116), .CO(n31794));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n31507), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_5 (.CI(n31507), .I0(n1607), .I1(n1631), .CO(n31508));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n31792), .O(n3206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_5 (.CI(n31792), .I0(n3107), .I1(n3116), .CO(n31793));
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n31506), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_4 (.CI(n31506), .I0(n1608), .I1(n1631), .CO(n31507));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n31791), .O(n3207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_10_lut (.I0(n19), .I1(bit_ctr[8]), .I2(GND_net), .I3(n30266), 
            .O(n42959)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_2143_4 (.CI(n31791), .I0(n3108), .I1(n3116), .CO(n31792));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n45866), 
            .I3(n31505), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n45863), 
            .I3(n31790), .O(n3208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_3 (.CI(n31505), .I0(n1609), .I1(n45866), .CO(n31506));
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n45866), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n45866), 
            .CO(n31505));
    SB_CARRY mod_5_add_2143_3 (.CI(n31790), .I0(n3109), .I1(n45863), .CO(n31791));
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n31504), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n45863), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n45863), 
            .CO(n31790));
    SB_LUT4 mod_5_add_1071_12_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n31503), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n31789), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_12 (.CI(n31503), .I0(n1500), .I1(n1532), .CO(n31504));
    SB_LUT4 add_21_33_lut (.I0(n19), .I1(bit_ctr[31]), .I2(GND_net), .I3(n30289), 
            .O(n42951)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n31788), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_11_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n31502), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_27 (.CI(n31788), .I0(n2985), .I1(n3017), .CO(n31789));
    SB_CARRY mod_5_add_1071_11 (.CI(n31502), .I0(n1501), .I1(n1532), .CO(n31503));
    SB_LUT4 mod_5_add_1071_10_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n31501), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n31787), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_26 (.CI(n31787), .I0(n2986), .I1(n3017), .CO(n31788));
    SB_CARRY mod_5_add_1071_10 (.CI(n31501), .I0(n1502), .I1(n1532), .CO(n31502));
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n31786), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_25 (.CI(n31786), .I0(n2987), .I1(n3017), .CO(n31787));
    SB_LUT4 mod_5_add_1071_9_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n31500), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n31785), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_9 (.CI(n31500), .I0(n1503), .I1(n1532), .CO(n31501));
    SB_CARRY mod_5_add_2076_24 (.CI(n31785), .I0(n2988), .I1(n3017), .CO(n31786));
    SB_LUT4 mod_5_add_1071_8_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n31499), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n31784), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_8 (.CI(n31499), .I0(n1504), .I1(n1532), .CO(n31500));
    SB_LUT4 mod_5_add_1071_7_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n31498), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_23 (.CI(n31784), .I0(n2989), .I1(n3017), .CO(n31785));
    SB_CARRY mod_5_add_1071_7 (.CI(n31498), .I0(n1505), .I1(n1532), .CO(n31499));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n31783), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_6_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n31497), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_22 (.CI(n31783), .I0(n2990), .I1(n3017), .CO(n31784));
    SB_CARRY mod_5_add_1071_6 (.CI(n31497), .I0(n1506), .I1(n1532), .CO(n31498));
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n31782), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_21 (.CI(n31782), .I0(n2991), .I1(n3017), .CO(n31783));
    SB_LUT4 mod_5_add_1071_5_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n31496), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n31781), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_5 (.CI(n31496), .I0(n1507), .I1(n1532), .CO(n31497));
    SB_CARRY mod_5_add_2076_20 (.CI(n31781), .I0(n2992), .I1(n3017), .CO(n31782));
    SB_LUT4 mod_5_add_1071_4_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n31495), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n31780), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_19 (.CI(n31780), .I0(n2993), .I1(n3017), .CO(n31781));
    SB_CARRY mod_5_add_1071_4 (.CI(n31495), .I0(n1508), .I1(n1532), .CO(n31496));
    SB_LUT4 mod_5_add_1071_3_lut (.I0(n1509), .I1(n1509), .I2(n45867), 
            .I3(n31494), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n31779), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_18 (.CI(n31779), .I0(n2994), .I1(n3017), .CO(n31780));
    SB_CARRY mod_5_add_1071_3 (.CI(n31494), .I0(n1509), .I1(n45867), .CO(n31495));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(bit_ctr[20]), .I1(bit_ctr[20]), .I2(n45867), 
            .I3(VCC_net), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(n45867), 
            .CO(n31494));
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1400), .I1(n1400), .I2(n1433), 
            .I3(n31493), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n31778), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_11_lut (.I0(n1401), .I1(n1401), .I2(n1433), 
            .I3(n31492), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_DFF timer_1147__i1 (.Q(timer[1]), .C(clk32MHz), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i2 (.Q(timer[2]), .C(clk32MHz), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY mod_5_add_2076_17 (.CI(n31778), .I0(n2995), .I1(n3017), .CO(n31779));
    SB_CARRY mod_5_add_1004_11 (.CI(n31492), .I0(n1401), .I1(n1433), .CO(n31493));
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n31777), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_16 (.CI(n31777), .I0(n2996), .I1(n3017), .CO(n31778));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(n1402), .I1(n1402), .I2(n1433), 
            .I3(n31491), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_10 (.CI(n31491), .I0(n1402), .I1(n1433), .CO(n31492));
    SB_LUT4 add_21_32_lut (.I0(n19), .I1(bit_ctr[30]), .I2(GND_net), .I3(n30288), 
            .O(n42950)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1004_9_lut (.I0(n1403), .I1(n1403), .I2(n1433), 
            .I3(n31490), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n31776), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_DFF timer_1147__i3 (.Q(timer[3]), .C(clk32MHz), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i4 (.Q(timer[4]), .C(clk32MHz), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i5 (.Q(timer[5]), .C(clk32MHz), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i6 (.Q(timer[6]), .C(clk32MHz), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i7 (.Q(timer[7]), .C(clk32MHz), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i8 (.Q(timer[8]), .C(clk32MHz), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i9 (.Q(timer[9]), .C(clk32MHz), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i10 (.Q(timer[10]), .C(clk32MHz), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i11 (.Q(timer[11]), .C(clk32MHz), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i12 (.Q(timer[12]), .C(clk32MHz), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i13 (.Q(timer[13]), .C(clk32MHz), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i14 (.Q(timer[14]), .C(clk32MHz), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i15 (.Q(timer[15]), .C(clk32MHz), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i16 (.Q(timer[16]), .C(clk32MHz), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i17 (.Q(timer[17]), .C(clk32MHz), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i18 (.Q(timer[18]), .C(clk32MHz), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i19 (.Q(timer[19]), .C(clk32MHz), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i20 (.Q(timer[20]), .C(clk32MHz), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i21 (.Q(timer[21]), .C(clk32MHz), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i22 (.Q(timer[22]), .C(clk32MHz), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i23 (.Q(timer[23]), .C(clk32MHz), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i24 (.Q(timer[24]), .C(clk32MHz), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i25 (.Q(timer[25]), .C(clk32MHz), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i26 (.Q(timer[26]), .C(clk32MHz), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i27 (.Q(timer[27]), .C(clk32MHz), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i28 (.Q(timer[28]), .C(clk32MHz), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i29 (.Q(timer[29]), .C(clk32MHz), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i30 (.Q(timer[30]), .C(clk32MHz), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1147__i31 (.Q(timer[31]), .C(clk32MHz), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_DFF start_103 (.Q(start), .C(clk32MHz), .D(n35977));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_2076_15 (.CI(n31776), .I0(n2997), .I1(n3017), .CO(n31777));
    SB_CARRY mod_5_add_1004_9 (.CI(n31490), .I0(n1403), .I1(n1433), .CO(n31491));
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n31775), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_8_lut (.I0(n1404), .I1(n1404), .I2(n1433), 
            .I3(n31489), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_8 (.CI(n31489), .I0(n1404), .I1(n1433), .CO(n31490));
    SB_LUT4 mod_5_add_1004_7_lut (.I0(n1405), .I1(n1405), .I2(n1433), 
            .I3(n31488), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_14 (.CI(n31775), .I0(n2998), .I1(n3017), .CO(n31776));
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n31774), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_13 (.CI(n31774), .I0(n2999), .I1(n3017), .CO(n31775));
    SB_CARRY mod_5_add_1004_7 (.CI(n31488), .I0(n1405), .I1(n1433), .CO(n31489));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n31773), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_12 (.CI(n31773), .I0(n3000), .I1(n3017), .CO(n31774));
    SB_LUT4 mod_5_add_1004_6_lut (.I0(n1406), .I1(n1406), .I2(n1433), 
            .I3(n31487), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_6 (.CI(n31487), .I0(n1406), .I1(n1433), .CO(n31488));
    SB_LUT4 i38738_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45861));
    defparam i38738_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n31772), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_11 (.CI(n31772), .I0(n3001), .I1(n3017), .CO(n31773));
    SB_LUT4 mod_5_add_1004_5_lut (.I0(n1407), .I1(n1407), .I2(n1433), 
            .I3(n31486), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_5 (.CI(n31486), .I0(n1407), .I1(n1433), .CO(n31487));
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n31771), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_4_lut (.I0(n1408), .I1(n1408), .I2(n1433), 
            .I3(n31485), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_32 (.CI(n30288), .I0(bit_ctr[30]), .I1(GND_net), .CO(n30289));
    SB_CARRY mod_5_add_2076_10 (.CI(n31771), .I0(n3002), .I1(n3017), .CO(n31772));
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n31770), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_4 (.CI(n31485), .I0(n1408), .I1(n1433), .CO(n31486));
    SB_CARRY mod_5_add_2076_9 (.CI(n31770), .I0(n3003), .I1(n3017), .CO(n31771));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(n1409), .I1(n1409), .I2(n45869), 
            .I3(n31484), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n31769), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_3 (.CI(n31484), .I0(n1409), .I1(n45869), .CO(n31485));
    SB_CARRY mod_5_add_2076_8 (.CI(n31769), .I0(n3004), .I1(n3017), .CO(n31770));
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n31768), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_2_lut (.I0(bit_ctr[21]), .I1(bit_ctr[21]), .I2(n45869), 
            .I3(VCC_net), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_7 (.CI(n31768), .I0(n3005), .I1(n3017), .CO(n31769));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n31767), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(n45869), 
            .CO(n31484));
    SB_CARRY mod_5_add_2076_6 (.CI(n31767), .I0(n3006), .I1(n3017), .CO(n31768));
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1301), .I1(n1301), .I2(n1334), 
            .I3(n31483), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_10_lut (.I0(n1302), .I1(n1302), .I2(n1334), 
            .I3(n31482), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_10 (.CI(n31482), .I0(n1302), .I1(n1334), .CO(n31483));
    SB_LUT4 mod_5_add_937_9_lut (.I0(n1303), .I1(n1303), .I2(n1334), .I3(n31481), 
            .O(n1402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_9 (.CI(n31481), .I0(n1303), .I1(n1334), .CO(n31482));
    SB_LUT4 mod_5_add_937_8_lut (.I0(n1304), .I1(n1304), .I2(n1334), .I3(n31480), 
            .O(n1403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n31766), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_8 (.CI(n31480), .I0(n1304), .I1(n1334), .CO(n31481));
    SB_LUT4 mod_5_add_937_7_lut (.I0(n1305), .I1(n1305), .I2(n1334), .I3(n31479), 
            .O(n1404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_5 (.CI(n31766), .I0(n3007), .I1(n3017), .CO(n31767));
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n31765), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_7 (.CI(n31479), .I0(n1305), .I1(n1334), .CO(n31480));
    SB_CARRY mod_5_add_2076_4 (.CI(n31765), .I0(n3008), .I1(n3017), .CO(n31766));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n3009), .I1(n3009), .I2(n45868), 
            .I3(n31764), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_937_6_lut (.I0(n1306), .I1(n1306), .I2(n1334), .I3(n31478), 
            .O(n1405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_6 (.CI(n31478), .I0(n1306), .I1(n1334), .CO(n31479));
    SB_CARRY mod_5_add_2076_3 (.CI(n31764), .I0(n3009), .I1(n45868), .CO(n31765));
    SB_LUT4 mod_5_add_937_5_lut (.I0(n1307), .I1(n1307), .I2(n1334), .I3(n31477), 
            .O(n1406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_5 (.CI(n31477), .I0(n1307), .I1(n1334), .CO(n31478));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n45868), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n45868), 
            .CO(n31764));
    SB_LUT4 mod_5_add_937_4_lut (.I0(n1308), .I1(n1308), .I2(n1334), .I3(n31476), 
            .O(n1407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n31763), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_4 (.CI(n31476), .I0(n1308), .I1(n1334), .CO(n31477));
    SB_LUT4 mod_5_add_2009_26_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n31762), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_26 (.CI(n31762), .I0(n2886), .I1(n2918), .CO(n31763));
    SB_LUT4 mod_5_add_2009_25_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n31761), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_25 (.CI(n31761), .I0(n2887), .I1(n2918), .CO(n31762));
    SB_LUT4 mod_5_add_937_3_lut (.I0(n1309), .I1(n1309), .I2(n45870), 
            .I3(n31475), .O(n1408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2009_24_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n31760), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_3 (.CI(n31475), .I0(n1309), .I1(n45870), .CO(n31476));
    SB_LUT4 mod_5_add_937_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[22]), .I2(n45870), 
            .I3(VCC_net), .O(n1409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(n45870), 
            .CO(n31475));
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n31474), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n31473), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n31473), .I0(n1203), .I1(n1235), .CO(n31474));
    SB_CARRY mod_5_add_2009_24 (.CI(n31760), .I0(n2888), .I1(n2918), .CO(n31761));
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n31472), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_23_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n31759), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_23 (.CI(n31759), .I0(n2889), .I1(n2918), .CO(n31760));
    SB_CARRY mod_5_add_870_8 (.CI(n31472), .I0(n1204), .I1(n1235), .CO(n31473));
    SB_LUT4 mod_5_add_2009_22_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n31758), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n31471), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_31_lut (.I0(n19), .I1(bit_ctr[29]), .I2(GND_net), .I3(n30287), 
            .O(n42946)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_31 (.CI(n30287), .I0(bit_ctr[29]), .I1(GND_net), .CO(n30288));
    SB_CARRY mod_5_add_2009_22 (.CI(n31758), .I0(n2890), .I1(n2918), .CO(n31759));
    SB_CARRY mod_5_add_870_7 (.CI(n31471), .I0(n1205), .I1(n1235), .CO(n31472));
    SB_LUT4 mod_5_add_2009_21_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n31757), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n31470), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_6 (.CI(n31470), .I0(n1206), .I1(n1235), .CO(n31471));
    SB_CARRY mod_5_add_2009_21 (.CI(n31757), .I0(n2891), .I1(n2918), .CO(n31758));
    SB_LUT4 mod_5_add_2009_20_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n31756), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n31469), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_5 (.CI(n31469), .I0(n1207), .I1(n1235), .CO(n31470));
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n31468), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_20 (.CI(n31756), .I0(n2892), .I1(n2918), .CO(n31757));
    SB_CARRY mod_5_add_870_4 (.CI(n31468), .I0(n1208), .I1(n1235), .CO(n31469));
    SB_LUT4 mod_5_add_2009_19_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n31755), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n45872), 
            .I3(n31467), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_19 (.CI(n31755), .I0(n2893), .I1(n2918), .CO(n31756));
    SB_CARRY mod_5_add_870_3 (.CI(n31467), .I0(n1209), .I1(n45872), .CO(n31468));
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n45872), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n45872), 
            .CO(n31467));
    SB_LUT4 mod_5_add_2009_18_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n31754), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n31466), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_18 (.CI(n31754), .I0(n2894), .I1(n2918), .CO(n31755));
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n31465), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_17_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n31753), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_8 (.CI(n31465), .I0(n1104), .I1(n1136), .CO(n31466));
    SB_CARRY mod_5_add_2009_17 (.CI(n31753), .I0(n2895), .I1(n2918), .CO(n31754));
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105_adj_4239), .I1(n1105_adj_4239), 
            .I2(n1136), .I3(n31464), .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_30_lut (.I0(n19), .I1(bit_ctr[28]), .I2(GND_net), .I3(n30286), 
            .O(n42945)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2009_16_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n31752), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_7 (.CI(n31464), .I0(n1105_adj_4239), .I1(n1136), 
            .CO(n31465));
    SB_CARRY mod_5_add_2009_16 (.CI(n31752), .I0(n2896), .I1(n2918), .CO(n31753));
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n31463), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_15_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n31751), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_15 (.CI(n31751), .I0(n2897), .I1(n2918), .CO(n31752));
    SB_CARRY mod_5_add_803_6 (.CI(n31463), .I0(n1106), .I1(n1136), .CO(n31464));
    SB_LUT4 mod_5_add_2009_14_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n31750), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n31462), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_5 (.CI(n31462), .I0(n1107), .I1(n1136), .CO(n31463));
    SB_CARRY mod_5_add_2009_14 (.CI(n31750), .I0(n2898), .I1(n2918), .CO(n31751));
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108_adj_4240), .I1(n1108_adj_4240), 
            .I2(n1136), .I3(n31461), .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_13_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n31749), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_13 (.CI(n31749), .I0(n2899), .I1(n2918), .CO(n31750));
    SB_CARRY mod_5_add_803_4 (.CI(n31461), .I0(n1108_adj_4240), .I1(n1136), 
            .CO(n31462));
    SB_CARRY add_21_30 (.CI(n30286), .I0(bit_ctr[28]), .I1(GND_net), .CO(n30287));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n31748), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_12 (.CI(n31748), .I0(n2900), .I1(n2918), .CO(n31749));
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n45873), 
            .I3(n31460), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_3 (.CI(n31460), .I0(n1109), .I1(n45873), .CO(n31461));
    SB_LUT4 mod_5_add_2009_11_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n31747), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n45873), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_11 (.CI(n31747), .I0(n2901), .I1(n2918), .CO(n31748));
    SB_LUT4 mod_5_add_2009_10_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n31746), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n45873), 
            .CO(n31460));
    SB_LUT4 mod_5_add_736_8_lut (.I0(n4_adj_4241), .I1(n4_adj_4241), .I2(n1037), 
            .I3(n31459), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_10 (.CI(n31746), .I0(n2902), .I1(n2918), .CO(n31747));
    SB_LUT4 mod_5_add_736_7_lut (.I0(n1005), .I1(n1005), .I2(n1037), .I3(n31458), 
            .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_9_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n31745), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_7 (.CI(n31458), .I0(n1005), .I1(n1037), .CO(n31459));
    SB_CARRY mod_5_add_2009_9 (.CI(n31745), .I0(n2903), .I1(n2918), .CO(n31746));
    SB_LUT4 mod_5_add_736_6_lut (.I0(n1006), .I1(n1006), .I2(n1037), .I3(n31457), 
            .O(n1105_adj_4239)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_8_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n31744), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_6 (.CI(n31457), .I0(n1006), .I1(n1037), .CO(n31458));
    SB_CARRY mod_5_add_2009_8 (.CI(n31744), .I0(n2904), .I1(n2918), .CO(n31745));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n31743), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_5_lut (.I0(n1007), .I1(n1007), .I2(n1037), .I3(n31456), 
            .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_5 (.CI(n31456), .I0(n1007), .I1(n1037), .CO(n31457));
    SB_CARRY mod_5_add_2009_7 (.CI(n31743), .I0(n2905), .I1(n2918), .CO(n31744));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n31742), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n31455), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_4 (.CI(n31455), .I0(n1008), .I1(n1037), .CO(n31456));
    SB_CARRY mod_5_add_2009_6 (.CI(n31742), .I0(n2906), .I1(n2918), .CO(n31743));
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n45874), 
            .I3(n31454), .O(n1108_adj_4240)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2009_5_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n31741), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_3 (.CI(n31454), .I0(n1009), .I1(n45874), .CO(n31455));
    SB_CARRY mod_5_add_2009_5 (.CI(n31741), .I0(n2907), .I1(n2918), .CO(n31742));
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n45874), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n45874), 
            .CO(n31454));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n31740), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(n905), .I2(VCC_net), 
            .I3(n31453), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_4 (.CI(n31740), .I0(n2908), .I1(n2918), .CO(n31741));
    SB_LUT4 mod_5_add_2009_3_lut (.I0(n2909), .I1(n2909), .I2(n45871), 
            .I3(n31739), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n31452), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_6 (.CI(n31452), .I0(n906), .I1(VCC_net), .CO(n31453));
    SB_CARRY mod_5_add_2009_3 (.CI(n31739), .I0(n2909), .I1(n45871), .CO(n31740));
    SB_LUT4 mod_5_add_2009_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[6]), .I2(n45871), 
            .I3(VCC_net), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n38039), .I2(VCC_net), 
            .I3(n31451), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_5 (.CI(n31451), .I0(n38039), .I1(VCC_net), 
            .CO(n31452));
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(n45871), 
            .CO(n31739));
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n18523), .I2(VCC_net), 
            .I3(n31450), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_4 (.CI(n31450), .I0(n18523), .I1(VCC_net), 
            .CO(n31451));
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n31738), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n31737), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n15788), .I2(GND_net), 
            .I3(n31449), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_3 (.CI(n31449), .I0(n15788), .I1(GND_net), 
            .CO(n31450));
    SB_CARRY mod_5_add_1942_25 (.CI(n31737), .I0(n2787), .I1(n2819), .CO(n31738));
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n31736), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n31449));
    SB_CARRY mod_5_add_1942_24 (.CI(n31736), .I0(n2788), .I1(n2819), .CO(n31737));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n31735), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_23 (.CI(n31735), .I0(n2789), .I1(n2819), .CO(n31736));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n31734), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_22 (.CI(n31734), .I0(n2790), .I1(n2819), .CO(n31735));
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n31733), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_21 (.CI(n31733), .I0(n2791), .I1(n2819), .CO(n31734));
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n31732), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_20 (.CI(n31732), .I0(n2792), .I1(n2819), .CO(n31733));
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n31731), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_19 (.CI(n31731), .I0(n2793), .I1(n2819), .CO(n31732));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n31730), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_18 (.CI(n31730), .I0(n2794), .I1(n2819), .CO(n31731));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n31729), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_DFFESR one_wire_108 (.Q(PIN_8_c), .C(clk32MHz), .E(n18367), .D(\neo_pixel_transmitter.done_N_576 ), 
            .R(n38456));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1942_17 (.CI(n31729), .I0(n2795), .I1(n2819), .CO(n31730));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n31728), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_16 (.CI(n31728), .I0(n2796), .I1(n2819), .CO(n31729));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n31727), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1147_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n31174), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1147_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n31173), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_15 (.CI(n31727), .I0(n2797), .I1(n2819), .CO(n31728));
    SB_CARRY timer_1147_add_4_32 (.CI(n31173), .I0(GND_net), .I1(timer[30]), 
            .CO(n31174));
    SB_LUT4 timer_1147_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n31172), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_10 (.CI(n30266), .I0(bit_ctr[8]), .I1(GND_net), .CO(n30267));
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n31726), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_14 (.CI(n31726), .I0(n2798), .I1(n2819), .CO(n31727));
    SB_CARRY timer_1147_add_4_31 (.CI(n31172), .I0(GND_net), .I1(timer[29]), 
            .CO(n31173));
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n31725), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_13 (.CI(n31725), .I0(n2799), .I1(n2819), .CO(n31726));
    SB_LUT4 timer_1147_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n31171), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n31724), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1147_add_4_30 (.CI(n31171), .I0(GND_net), .I1(timer[28]), 
            .CO(n31172));
    SB_LUT4 timer_1147_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n31170), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_12 (.CI(n31724), .I0(n2800), .I1(n2819), .CO(n31725));
    SB_CARRY timer_1147_add_4_29 (.CI(n31170), .I0(GND_net), .I1(timer[27]), 
            .CO(n31171));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n31723), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1147_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n31169), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_11 (.CI(n31723), .I0(n2801), .I1(n2819), .CO(n31724));
    SB_CARRY timer_1147_add_4_28 (.CI(n31169), .I0(GND_net), .I1(timer[26]), 
            .CO(n31170));
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n31722), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_10 (.CI(n31722), .I0(n2802), .I1(n2819), .CO(n31723));
    SB_LUT4 timer_1147_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n31168), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n31721), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1147_add_4_27 (.CI(n31168), .I0(GND_net), .I1(timer[25]), 
            .CO(n31169));
    SB_CARRY mod_5_add_1942_9 (.CI(n31721), .I0(n2803), .I1(n2819), .CO(n31722));
    SB_LUT4 timer_1147_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n31167), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1147_add_4_26 (.CI(n31167), .I0(GND_net), .I1(timer[24]), 
            .CO(n31168));
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n31720), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1147_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n31166), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_29_lut (.I0(n11), .I1(bit_ctr[27]), .I2(GND_net), .I3(n30285), 
            .O(n42939)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1942_8 (.CI(n31720), .I0(n2804), .I1(n2819), .CO(n31721));
    SB_CARRY timer_1147_add_4_25 (.CI(n31166), .I0(GND_net), .I1(timer[23]), 
            .CO(n31167));
    SB_LUT4 timer_1147_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n31165), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n31719), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1147_add_4_24 (.CI(n31165), .I0(GND_net), .I1(timer[22]), 
            .CO(n31166));
    SB_CARRY mod_5_add_1942_7 (.CI(n31719), .I0(n2805), .I1(n2819), .CO(n31720));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n31718), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_6 (.CI(n31718), .I0(n2806), .I1(n2819), .CO(n31719));
    SB_LUT4 timer_1147_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n31164), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1147_add_4_17 (.CI(n31158), .I0(GND_net), .I1(timer[15]), 
            .CO(n31159));
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n31717), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_5 (.CI(n31717), .I0(n2807), .I1(n2819), .CO(n31718));
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n31716), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_4 (.CI(n31716), .I0(n2808), .I1(n2819), .CO(n31717));
    SB_LUT4 sub_14_add_2_33_lut (.I0(one_wire_N_513[22]), .I1(timer[31]), 
            .I2(n1[31]), .I3(n30432), .O(n19_adj_4228)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_14_add_2_32_lut (.I0(one_wire_N_513[25]), .I1(timer[30]), 
            .I2(n1[30]), .I3(n30431), .O(n21_adj_4222)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_29 (.CI(n30285), .I0(bit_ctr[27]), .I1(GND_net), .CO(n30286));
    SB_CARRY sub_14_add_2_32 (.CI(n30431), .I0(timer[30]), .I1(n1[30]), 
            .CO(n30432));
    SB_LUT4 add_21_2_lut (.I0(n19), .I1(bit_ctr[0]), .I2(GND_net), .I3(VCC_net), 
            .O(n42940)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_14_add_2_31_lut (.I0(GND_net), .I1(timer[29]), .I2(n1[29]), 
            .I3(n30430), .O(one_wire_N_513[29])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n45875), 
            .I3(n31715), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_3 (.CI(n31715), .I0(n2809), .I1(n45875), .CO(n31716));
    SB_LUT4 add_21_9_lut (.I0(n19), .I1(bit_ctr[7]), .I2(GND_net), .I3(n30265), 
            .O(n42958)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_28_lut (.I0(n11), .I1(bit_ctr[26]), .I2(GND_net), .I3(n30284), 
            .O(n42936)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n45875), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY sub_14_add_2_31 (.CI(n30430), .I0(timer[29]), .I1(n1[29]), 
            .CO(n30431));
    SB_LUT4 sub_14_add_2_30_lut (.I0(one_wire_N_513[26]), .I1(timer[28]), 
            .I2(n1[28]), .I3(n30429), .O(n22_adj_4223)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n45875), 
            .CO(n31715));
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n31714), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_24_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n31713), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_24 (.CI(n31713), .I0(n2688), .I1(n2720), .CO(n31714));
    SB_LUT4 mod_5_add_1875_23_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n31712), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_30 (.CI(n30429), .I0(timer[28]), .I1(n1[28]), 
            .CO(n30430));
    SB_CARRY mod_5_add_1875_23 (.CI(n31712), .I0(n2689), .I1(n2720), .CO(n31713));
    SB_LUT4 sub_14_add_2_29_lut (.I0(one_wire_N_513[18]), .I1(timer[27]), 
            .I2(n1[27]), .I3(n30428), .O(n18_adj_4200)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1875_22_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n31711), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_29 (.CI(n30428), .I0(timer[27]), .I1(n1[27]), 
            .CO(n30429));
    SB_LUT4 i15_4_lut_adj_1514 (.I0(n3107), .I1(n3097), .I2(n3105), .I3(n3090), 
            .O(n42));
    defparam i15_4_lut_adj_1514.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1875_22 (.CI(n31711), .I0(n2690), .I1(n2720), .CO(n31712));
    SB_LUT4 mod_5_add_1875_21_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n31710), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_28_lut (.I0(GND_net), .I1(timer[26]), .I2(n1[26]), 
            .I3(n30427), .O(one_wire_N_513[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19_4_lut_adj_1515 (.I0(n3083), .I1(n3095), .I2(n3101), .I3(n3103), 
            .O(n46));
    defparam i19_4_lut_adj_1515.LUT_INIT = 16'hfffe;
    SB_CARRY add_21_28 (.CI(n30284), .I0(bit_ctr[26]), .I1(GND_net), .CO(n30285));
    SB_LUT4 i17_4_lut_adj_1516 (.I0(n3092), .I1(n3102), .I2(n3098), .I3(n3086), 
            .O(n44));
    defparam i17_4_lut_adj_1516.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_27_lut (.I0(n11), .I1(bit_ctr[25]), .I2(GND_net), .I3(n30283), 
            .O(n42935)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i18_4_lut_adj_1517 (.I0(n3093), .I1(n3108), .I2(n3088), .I3(n3100), 
            .O(n45));
    defparam i18_4_lut_adj_1517.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1518 (.I0(n3089), .I1(n3096), .I2(n3094), .I3(n3091), 
            .O(n43));
    defparam i16_4_lut_adj_1518.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1875_21 (.CI(n31710), .I0(n2691), .I1(n2720), .CO(n31711));
    SB_CARRY sub_14_add_2_28 (.CI(n30427), .I0(timer[26]), .I1(n1[26]), 
            .CO(n30428));
    SB_CARRY add_21_9 (.CI(n30265), .I0(bit_ctr[7]), .I1(GND_net), .CO(n30266));
    SB_LUT4 sub_14_add_2_27_lut (.I0(GND_net), .I1(timer[25]), .I2(n1[25]), 
            .I3(n30426), .O(one_wire_N_513[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1875_20_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n31709), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_27 (.CI(n30283), .I0(bit_ctr[25]), .I1(GND_net), .CO(n30284));
    SB_CARRY mod_5_add_1875_20 (.CI(n31709), .I0(n2692), .I1(n2720), .CO(n31710));
    SB_CARRY sub_14_add_2_27 (.CI(n30426), .I0(timer[25]), .I1(n1[25]), 
            .CO(n30427));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n31708), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_19 (.CI(n31708), .I0(n2693), .I1(n2720), .CO(n31709));
    SB_LUT4 mod_5_add_1875_18_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n31707), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk32MHz), .D(n18663));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i13_2_lut (.I0(n3087), .I1(n3084), .I2(GND_net), .I3(GND_net), 
            .O(n40_adj_4246));
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_1875_18 (.CI(n31707), .I0(n2694), .I1(n2720), .CO(n31708));
    SB_LUT4 i21_4_lut_adj_1519 (.I0(n3106), .I1(n42), .I2(n3085), .I3(n3099), 
            .O(n48));
    defparam i21_4_lut_adj_1519.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n43), .I1(n45), .I2(n44), .I3(n46), .O(n52));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1875_17_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n31706), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_17 (.CI(n31706), .I0(n2695), .I1(n2720), .CO(n31707));
    SB_LUT4 i12_3_lut (.I0(n3104), .I1(bit_ctr[4]), .I2(n3109), .I3(GND_net), 
            .O(n39_adj_4247));
    defparam i12_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 mod_5_add_1875_16_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n31705), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_16 (.CI(n31705), .I0(n2696), .I1(n2720), .CO(n31706));
    SB_LUT4 i26_4_lut (.I0(n39_adj_4247), .I1(n52), .I2(n48), .I3(n40_adj_4246), 
            .O(n3116));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1875_15_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n31704), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_26_lut (.I0(GND_net), .I1(timer[24]), .I2(n1[24]), 
            .I3(n30425), .O(one_wire_N_513[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n30259));
    SB_CARRY mod_5_add_1875_15 (.CI(n31704), .I0(n2697), .I1(n2720), .CO(n31705));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n31703), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_26 (.CI(n30425), .I0(timer[24]), .I1(n1[24]), 
            .CO(n30426));
    SB_CARRY mod_5_add_1875_14 (.CI(n31703), .I0(n2698), .I1(n2720), .CO(n31704));
    SB_LUT4 mod_5_add_1875_13_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n31702), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_13 (.CI(n31702), .I0(n2699), .I1(n2720), .CO(n31703));
    SB_LUT4 mod_5_add_1875_12_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n31701), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_12 (.CI(n31701), .I0(n2700), .I1(n2720), .CO(n31702));
    SB_LUT4 mod_5_add_1875_11_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n31700), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_26_lut (.I0(n11), .I1(bit_ctr[24]), .I2(GND_net), .I3(n30282), 
            .O(n42934)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1875_11 (.CI(n31700), .I0(n2701), .I1(n2720), .CO(n31701));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n31699), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_8_lut (.I0(n19), .I1(bit_ctr[6]), .I2(GND_net), .I3(n30264), 
            .O(n42957)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_26 (.CI(n30282), .I0(bit_ctr[24]), .I1(GND_net), .CO(n30283));
    SB_LUT4 add_21_25_lut (.I0(n11), .I1(bit_ctr[23]), .I2(GND_net), .I3(n30281), 
            .O(n42933)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_25 (.CI(n30281), .I0(bit_ctr[23]), .I1(GND_net), .CO(n30282));
    SB_LUT4 sub_14_add_2_25_lut (.I0(one_wire_N_513[17]), .I1(timer[23]), 
            .I2(n1[23]), .I3(n30424), .O(n25_adj_4226)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1875_10 (.CI(n31699), .I0(n2702), .I1(n2720), .CO(n31700));
    SB_LUT4 add_21_24_lut (.I0(n19), .I1(bit_ctr[22]), .I2(GND_net), .I3(n30280), 
            .O(n42944)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1875_9_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n31698), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_9 (.CI(n31698), .I0(n2703), .I1(n2720), .CO(n31699));
    SB_CARRY add_21_24 (.CI(n30280), .I0(bit_ctr[22]), .I1(GND_net), .CO(n30281));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n31697), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_8 (.CI(n31697), .I0(n2704), .I1(n2720), .CO(n31698));
    SB_LUT4 timer_1147_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n31158), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_25 (.CI(n30424), .I0(timer[23]), .I1(n1[23]), 
            .CO(n30425));
    SB_LUT4 add_21_23_lut (.I0(n19), .I1(bit_ctr[21]), .I2(GND_net), .I3(n30279), 
            .O(n42942)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1875_7_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n31696), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1147_add_4_18 (.CI(n31159), .I0(GND_net), .I1(timer[16]), 
            .CO(n31160));
    SB_CARRY add_21_23 (.CI(n30279), .I0(bit_ctr[21]), .I1(GND_net), .CO(n30280));
    SB_CARRY mod_5_add_1875_7 (.CI(n31696), .I0(n2705), .I1(n2720), .CO(n31697));
    SB_LUT4 timer_1147_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n31159), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1147_add_4_19 (.CI(n31160), .I0(GND_net), .I1(timer[17]), 
            .CO(n31161));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n31695), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_6 (.CI(n31695), .I0(n2706), .I1(n2720), .CO(n31696));
    SB_LUT4 timer_1147_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n31160), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1875_5_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n31694), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1147_add_4_20 (.CI(n31161), .I0(GND_net), .I1(timer[18]), 
            .CO(n31162));
    SB_LUT4 sub_14_add_2_24_lut (.I0(GND_net), .I1(timer[22]), .I2(n1[22]), 
            .I3(n30423), .O(one_wire_N_513[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_24 (.CI(n30423), .I0(timer[22]), .I1(n1[22]), 
            .CO(n30424));
    SB_LUT4 timer_1147_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n31161), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_23_lut (.I0(n39589), .I1(timer[21]), .I2(n1[21]), 
            .I3(n30422), .O(n23_adj_4225)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY timer_1147_add_4_21 (.CI(n31162), .I0(GND_net), .I1(timer[19]), 
            .CO(n31163));
    SB_CARRY sub_14_add_2_23 (.CI(n30422), .I0(timer[21]), .I1(n1[21]), 
            .CO(n30423));
    SB_LUT4 add_21_22_lut (.I0(n19), .I1(bit_ctr[20]), .I2(GND_net), .I3(n30278), 
            .O(n42941)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_14_add_2_22_lut (.I0(GND_net), .I1(timer[20]), .I2(n1[20]), 
            .I3(n30421), .O(one_wire_N_513[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_22 (.CI(n30278), .I0(bit_ctr[20]), .I1(GND_net), .CO(n30279));
    SB_CARRY sub_14_add_2_22 (.CI(n30421), .I0(timer[20]), .I1(n1[20]), 
            .CO(n30422));
    SB_CARRY mod_5_add_1875_5 (.CI(n31694), .I0(n2707), .I1(n2720), .CO(n31695));
    SB_LUT4 timer_1147_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n31162), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_21_lut (.I0(n19), .I1(bit_ctr[19]), .I2(GND_net), .I3(n30277), 
            .O(n42949)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1875_4_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n31693), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1147_add_4_22 (.CI(n31163), .I0(GND_net), .I1(timer[20]), 
            .CO(n31164));
    SB_LUT4 sub_14_add_2_21_lut (.I0(GND_net), .I1(timer[19]), .I2(n1[19]), 
            .I3(n30420), .O(one_wire_N_513[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_4 (.CI(n31693), .I0(n2708), .I1(n2720), .CO(n31694));
    SB_LUT4 timer_1147_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n31163), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1147_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1147_add_4_23 (.CI(n31164), .I0(GND_net), .I1(timer[21]), 
            .CO(n31165));
    SB_CARRY sub_14_add_2_21 (.CI(n30420), .I0(timer[19]), .I1(n1[19]), 
            .CO(n30421));
    SB_CARRY add_21_8 (.CI(n30264), .I0(bit_ctr[6]), .I1(GND_net), .CO(n30265));
    SB_LUT4 sub_14_add_2_20_lut (.I0(GND_net), .I1(timer[18]), .I2(n1[18]), 
            .I3(n30419), .O(one_wire_N_513[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1875_3_lut (.I0(n2709), .I1(n2709), .I2(n45876), 
            .I3(n31692), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY sub_14_add_2_20 (.CI(n30419), .I0(timer[18]), .I1(n1[18]), 
            .CO(n30420));
    SB_LUT4 sub_14_add_2_19_lut (.I0(GND_net), .I1(timer[17]), .I2(n1[17]), 
            .I3(n30418), .O(one_wire_N_513[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_3 (.CI(n31692), .I0(n2709), .I1(n45876), .CO(n31693));
    SB_LUT4 mod_5_add_1875_2_lut (.I0(bit_ctr[8]), .I1(bit_ctr[8]), .I2(n45876), 
            .I3(VCC_net), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_21_21 (.CI(n30277), .I0(bit_ctr[19]), .I1(GND_net), .CO(n30278));
    SB_LUT4 add_21_20_lut (.I0(n19), .I1(bit_ctr[18]), .I2(GND_net), .I3(n30276), 
            .O(n42948)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(n45876), 
            .CO(n31692));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n31691), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n31690), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_20 (.CI(n30276), .I0(bit_ctr[18]), .I1(GND_net), .CO(n30277));
    SB_CARRY mod_5_add_1808_23 (.CI(n31690), .I0(n2589), .I1(n2621), .CO(n31691));
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n31689), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_22 (.CI(n31689), .I0(n2590), .I1(n2621), .CO(n31690));
    SB_LUT4 i14_4_lut_adj_1520 (.I0(n1105), .I1(n4724), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n4754));
    defparam i14_4_lut_adj_1520.LUT_INIT = 16'hcfca;
    SB_LUT4 i10_4_lut_adj_1521 (.I0(n1806), .I1(n1803), .I2(n1805), .I3(n1798), 
            .O(n24_adj_4251));
    defparam i10_4_lut_adj_1521.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1522 (.I0(n1808), .I1(n1804), .I2(n1802), .I3(n1801), 
            .O(n22_adj_4252));
    defparam i8_4_lut_adj_1522.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1523 (.I0(n1800), .I1(n1799), .I2(n1797), .I3(n1807), 
            .O(n23_adj_4253));
    defparam i9_4_lut_adj_1523.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1524 (.I0(n1796), .I1(bit_ctr[17]), .I2(n1809), 
            .I3(GND_net), .O(n21_adj_4254));
    defparam i7_3_lut_adj_1524.LUT_INIT = 16'heaea;
    SB_LUT4 i13_4_lut_adj_1525 (.I0(n21_adj_4254), .I1(n23_adj_4253), .I2(n22_adj_4252), 
            .I3(n24_adj_4251), .O(n1829));
    defparam i13_4_lut_adj_1525.LUT_INIT = 16'hfffe;
    SB_LUT4 i38737_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45860));
    defparam i38737_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22325_3_lut (.I0(one_wire_N_513[9]), .I1(\one_wire_N_513[11] ), 
            .I2(one_wire_N_513[10]), .I3(GND_net), .O(n27335));
    defparam i22325_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1526 (.I0(\state[0] ), .I1(n4_adj_4255), .I2(n1108), 
            .I3(\state[1] ), .O(n18416));
    defparam i1_4_lut_adj_1526.LUT_INIT = 16'hafcc;
    SB_LUT4 i15_4_lut_adj_1527 (.I0(n4_adj_4255), .I1(\state[0] ), .I2(\state[1] ), 
            .I3(n1108), .O(n18584));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15_4_lut_adj_1527.LUT_INIT = 16'h0a3a;
    SB_LUT4 i31109_4_lut (.I0(n17064), .I1(n32476), .I2(n4_adj_4216), 
            .I3(\state[0] ), .O(n27453));
    defparam i31109_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i3_4_lut (.I0(n5_adj_4229), .I1(\state[1] ), .I2(n17064), 
            .I3(n38076), .O(n39504));
    defparam i3_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i2_4_lut (.I0(\state[1] ), .I1(n39504), .I2(start), .I3(n39505), 
            .O(n39307));
    defparam i2_4_lut.LUT_INIT = 16'h8c00;
    SB_LUT4 i11_4_lut_adj_1528 (.I0(n1895), .I1(n1902), .I2(n1899), .I3(n1897), 
            .O(n26_adj_4256));
    defparam i11_4_lut_adj_1528.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1529 (.I0(n1907), .I1(bit_ctr[16]), .I2(n1909), 
            .I3(GND_net), .O(n19_adj_4257));
    defparam i4_3_lut_adj_1529.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut_adj_1530 (.I0(n1908), .I1(n1900), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4258));
    defparam i1_2_lut_adj_1530.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1531 (.I0(n1904), .I1(n1901), .I2(n1906), .I3(n1898), 
            .O(n24_adj_4259));
    defparam i9_4_lut_adj_1531.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1532 (.I0(n19_adj_4257), .I1(n26_adj_4256), .I2(n1905), 
            .I3(n1903), .O(n28_adj_4260));
    defparam i13_4_lut_adj_1532.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1533 (.I0(n1896), .I1(n28_adj_4260), .I2(n24_adj_4259), 
            .I3(n16_adj_4258), .O(n1928));
    defparam i14_4_lut_adj_1533.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1534 (.I0(n2193), .I1(n2194), .I2(n2206), .I3(n2204), 
            .O(n28_adj_4261));
    defparam i10_4_lut_adj_1534.LUT_INIT = 16'hfffe;
    SB_LUT4 i38736_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45859));
    defparam i38736_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut_adj_1535 (.I0(n2203), .I1(n28_adj_4261), .I2(bit_ctr[13]), 
            .I3(n2209), .O(n32_adj_4262));
    defparam i14_4_lut_adj_1535.LUT_INIT = 16'hfeee;
    SB_LUT4 i12_4_lut_adj_1536 (.I0(n2208), .I1(n2201), .I2(n2192), .I3(n2196), 
            .O(n30_adj_4263));
    defparam i12_4_lut_adj_1536.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1537 (.I0(n2195), .I1(n2207), .I2(n2205), .I3(n2199), 
            .O(n31_adj_4264));
    defparam i13_4_lut_adj_1537.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1538 (.I0(n27_adj_4213), .I1(n29_adj_4214), .I2(n28_adj_4215), 
            .I3(n30_adj_4265), .O(n33679));
    defparam i16_4_lut_adj_1538.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1539 (.I0(n2202), .I1(n2197), .I2(n2198), .I3(n2200), 
            .O(n29_adj_4266));
    defparam i11_4_lut_adj_1539.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1540 (.I0(n29_adj_4266), .I1(n31_adj_4264), .I2(n30_adj_4263), 
            .I3(n32_adj_4262), .O(n2225));
    defparam i17_4_lut_adj_1540.LUT_INIT = 16'hfffe;
    SB_LUT4 i38733_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45856));
    defparam i38733_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3433_2_lut_4_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(bit_ctr[29]), 
            .I3(bit_ctr[28]), .O(n7476));   // verilog/neopixel.v(22[26:36])
    defparam i3433_2_lut_4_lut.LUT_INIT = 16'h9400;
    SB_LUT4 i31133_2_lut_3_lut (.I0(n38192), .I1(one_wire_N_513[4]), .I2(n38086), 
            .I3(GND_net), .O(n38194));
    defparam i31133_2_lut_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut_3_lut (.I0(bit_ctr[3]), .I1(bit_ctr[4]), .I2(n33679), 
            .I3(GND_net), .O(\state_3__N_362[1] ));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hf8f8;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i38753_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45876));
    defparam i38753_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6_3_lut_adj_1541 (.I0(bit_ctr[26]), .I1(bit_ctr[13]), .I2(bit_ctr[11]), 
            .I3(GND_net), .O(n17_adj_4267));
    defparam i6_3_lut_adj_1541.LUT_INIT = 16'hfefe;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i3_2_lut_adj_1542 (.I0(n5), .I1(n6), .I2(GND_net), .I3(GND_net), 
            .O(n39589));   // verilog/neopixel.v(104[14:39])
    defparam i3_2_lut_adj_1542.LUT_INIT = 16'heeee;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut_adj_1543 (.I0(n27453), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[1] ), .O(n39505));
    defparam i2_3_lut_4_lut_adj_1543.LUT_INIT = 16'hffdf;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23_3_lut_4_lut (.I0(n27172), .I1(one_wire_N_513[4]), .I2(n32476), 
            .I3(\state[0] ), .O(n38076));
    defparam i23_3_lut_4_lut.LUT_INIT = 16'hf0ee;
    SB_LUT4 i1_2_lut_3_lut_adj_1544 (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(n27453), .I3(GND_net), .O(n4_adj_4255));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_2_lut_3_lut_adj_1544.LUT_INIT = 16'h4040;
    SB_LUT4 i6_3_lut_adj_1545 (.I0(n2689), .I1(bit_ctr[8]), .I2(n2709), 
            .I3(GND_net), .O(n29_adj_4268));
    defparam i6_3_lut_adj_1545.LUT_INIT = 16'heaea;
    SB_LUT4 i14_4_lut_adj_1546 (.I0(n2700), .I1(n2701), .I2(n2702), .I3(n2688), 
            .O(n37_adj_4269));
    defparam i14_4_lut_adj_1546.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1547 (.I0(n2687), .I1(n2703), .I2(n2697), .I3(n2699), 
            .O(n36_adj_4270));
    defparam i13_4_lut_adj_1547.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1548 (.I0(n37_adj_4269), .I1(n29_adj_4268), .I2(n2692), 
            .I3(n2691), .O(n42_adj_4271));
    defparam i19_4_lut_adj_1548.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1549 (.I0(n2695), .I1(n2690), .I2(n2707), .I3(n2693), 
            .O(n40_adj_4272));
    defparam i17_4_lut_adj_1549.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1550 (.I0(n2706), .I1(n36_adj_4270), .I2(n2694), 
            .I3(n2704), .O(n41));
    defparam i18_4_lut_adj_1550.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1551 (.I0(n2708), .I1(n2705), .I2(n2696), .I3(n2698), 
            .O(n39_adj_4273));
    defparam i16_4_lut_adj_1551.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n39_adj_4273), .I1(n41), .I2(n40_adj_4272), 
            .I3(n42_adj_4271), .O(n2720));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i38752_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45875));
    defparam i38752_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i31113_2_lut (.I0(one_wire_N_513[4]), .I1(n38086), .I2(GND_net), 
            .I3(GND_net), .O(n38174));
    defparam i31113_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i130_4_lut (.I0(n27335), .I1(n38194), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[1] ), .O(n103));
    defparam i130_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i1_4_lut_adj_1552 (.I0(n38192), .I1(n38174), .I2(n4_adj_4216), 
            .I3(n37332), .O(n37231));
    defparam i1_4_lut_adj_1552.LUT_INIT = 16'h1505;
    SB_LUT4 i1_4_lut_adj_1553 (.I0(n17206), .I1(\state[0] ), .I2(n37231), 
            .I3(n103), .O(n18367));
    defparam i1_4_lut_adj_1553.LUT_INIT = 16'h5150;
    SB_LUT4 i86_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_576 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i86_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i16_4_lut_adj_1554 (.I0(n2798), .I1(n2804), .I2(n2791), .I3(n2795), 
            .O(n40_adj_4274));
    defparam i16_4_lut_adj_1554.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1555 (.I0(n2796), .I1(n2793), .I2(n2788), .I3(n2808), 
            .O(n38_adj_4275));
    defparam i14_4_lut_adj_1555.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1556 (.I0(n2789), .I1(n2800), .I2(n2803), .I3(n2805), 
            .O(n39_adj_4276));
    defparam i15_4_lut_adj_1556.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1557 (.I0(n2792), .I1(n2787), .I2(n2801), .I3(n2799), 
            .O(n37_adj_4277));
    defparam i13_4_lut_adj_1557.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_2_lut (.I0(n2786), .I1(n2797), .I2(GND_net), .I3(GND_net), 
            .O(n34_adj_4278));
    defparam i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i18_4_lut_adj_1558 (.I0(n2794), .I1(n2806), .I2(n2807), .I3(n2790), 
            .O(n42_adj_4279));
    defparam i18_4_lut_adj_1558.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1559 (.I0(n37_adj_4277), .I1(n39_adj_4276), .I2(n38_adj_4275), 
            .I3(n40_adj_4274), .O(n46_adj_4280));
    defparam i22_4_lut_adj_1559.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_3_lut (.I0(bit_ctr[7]), .I1(n2802), .I2(n2809), .I3(GND_net), 
            .O(n33_adj_4281));
    defparam i9_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i23_4_lut (.I0(n33_adj_4281), .I1(n46_adj_4280), .I2(n42_adj_4279), 
            .I3(n34_adj_4278), .O(n2819));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i38748_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45871));
    defparam i38748_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i38751_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45874));
    defparam i38751_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i38721_2_lut (.I0(n33784), .I1(n971[28]), .I2(GND_net), .I3(GND_net), 
            .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i38721_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i38719_2_lut (.I0(n33784), .I1(n971[29]), .I2(GND_net), .I3(GND_net), 
            .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam i38719_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_i672_3_lut (.I0(n906), .I1(n971[30]), .I2(n33784), .I3(GND_net), 
            .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i605_3_lut_4_lut (.I0(n708), .I1(n7476), .I2(n60), .I3(n838), 
            .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_3_lut_4_lut.LUT_INIT = 16'h8887;
    SB_LUT4 mod_5_i604_4_lut_4_lut (.I0(n708), .I1(n7476), .I2(n838), 
            .I3(n60), .O(n905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i604_4_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i36445_3_lut (.I0(n15780), .I1(bit_ctr[27]), .I2(n838), .I3(GND_net), 
            .O(n18523));
    defparam i36445_3_lut.LUT_INIT = 16'h5959;
    SB_LUT4 i3_4_lut_adj_1560 (.I0(bit_ctr[26]), .I1(n906), .I2(n15788), 
            .I3(n18523), .O(n8_adj_4282));   // verilog/neopixel.v(22[26:36])
    defparam i3_4_lut_adj_1560.LUT_INIT = 16'h0013;
    SB_LUT4 i4_3_lut_adj_1561 (.I0(n38039), .I1(n8_adj_4282), .I2(n905), 
            .I3(GND_net), .O(n33784));   // verilog/neopixel.v(22[26:36])
    defparam i4_3_lut_adj_1561.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_adj_1562 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n15788));
    defparam i1_2_lut_adj_1562.LUT_INIT = 16'h9999;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n33784), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i675_3_lut (.I0(n15788), .I1(n971[27]), .I2(n33784), 
            .I3(GND_net), .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33759_3_lut (.I0(n971[28]), .I1(n971[31]), .I2(n971[29]), 
            .I3(GND_net), .O(n40825));
    defparam i33759_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_adj_1563 (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), 
            .I3(GND_net), .O(n6_adj_4283));
    defparam i2_3_lut_adj_1563.LUT_INIT = 16'heaea;
    SB_LUT4 i3_4_lut_adj_1564 (.I0(n33784), .I1(n6_adj_4283), .I2(n1005), 
            .I3(n40825), .O(n1037));
    defparam i3_4_lut_adj_1564.LUT_INIT = 16'hfdfc;
    SB_LUT4 i38717_2_lut (.I0(n33784), .I1(n971[31]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_4241));   // verilog/neopixel.v(22[26:36])
    defparam i38717_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i38750_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45873));
    defparam i38750_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22343_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n27353));
    defparam i22343_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(n1105_adj_4239), .I1(n1103), .I2(n27353), .I3(n1108_adj_4240), 
            .O(n12_adj_4284));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1565 (.I0(n1107), .I1(n12_adj_4284), .I2(n1106), 
            .I3(n1104), .O(n1136));
    defparam i6_4_lut_adj_1565.LUT_INIT = 16'hfffe;
    SB_LUT4 i38749_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45872));
    defparam i38749_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6_4_lut_adj_1566 (.I0(n1205), .I1(n1206), .I2(n1204), .I3(n1207), 
            .O(n14_adj_4285));
    defparam i6_4_lut_adj_1566.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1567 (.I0(bit_ctr[23]), .I1(n1203), .I2(n1209), 
            .I3(GND_net), .O(n9_adj_4286));
    defparam i1_3_lut_adj_1567.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut (.I0(n9_adj_4286), .I1(n14_adj_4285), .I2(n1202), 
            .I3(n1208), .O(n1235));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i38747_1_lut (.I0(n1334), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45870));
    defparam i38747_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_3_lut (.I0(bit_ctr[6]), .I1(n2907), .I2(n2909), .I3(GND_net), 
            .O(n33_adj_4287));
    defparam i8_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i16_4_lut_adj_1568 (.I0(n2900), .I1(n2891), .I2(n2897), .I3(n2888), 
            .O(n41_adj_4288));
    defparam i16_4_lut_adj_1568.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n2906), .I1(n2887), .I2(n2892), .I3(GND_net), 
            .O(n38_adj_4289));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut_adj_1569 (.I0(n2896), .I1(n2885), .I2(n2905), .I3(n2902), 
            .O(n43_adj_4290));
    defparam i18_4_lut_adj_1569.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1570 (.I0(n2899), .I1(n2890), .I2(n2898), .I3(n2908), 
            .O(n40_adj_4291));
    defparam i15_4_lut_adj_1570.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1571 (.I0(n41_adj_4288), .I1(n33_adj_4287), .I2(n2889), 
            .I3(n2901), .O(n46_adj_4292));
    defparam i21_4_lut_adj_1571.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1572 (.I0(n2886), .I1(n2894), .I2(n2895), .I3(n2903), 
            .O(n39_adj_4293));
    defparam i14_4_lut_adj_1572.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1573 (.I0(n43_adj_4290), .I1(n2904), .I2(n38_adj_4289), 
            .I3(n2893), .O(n47));
    defparam i22_4_lut_adj_1573.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n47), .I1(n39_adj_4293), .I2(n46_adj_4292), 
            .I3(n40_adj_4291), .O(n2918));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i38745_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45868));
    defparam i38745_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_4_lut_adj_1574 (.I0(bit_ctr[9]), .I1(bit_ctr[8]), .I2(bit_ctr[18]), 
            .I3(bit_ctr[10]), .O(n19_adj_4294));
    defparam i8_4_lut_adj_1574.LUT_INIT = 16'hfffe;
    SB_LUT4 i36451_3_lut_4_lut_4_lut (.I0(n708), .I1(n7476), .I2(n32958), 
            .I3(bit_ctr[28]), .O(n38037));   // verilog/neopixel.v(22[26:36])
    defparam i36451_3_lut_4_lut_4_lut.LUT_INIT = 16'h1ef0;
    SB_LUT4 i1_2_lut_adj_1575 (.I0(n1304), .I1(n1305), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_4295));
    defparam i1_2_lut_adj_1575.LUT_INIT = 16'heeee;
    SB_LUT4 i3_3_lut (.I0(bit_ctr[22]), .I1(n1303), .I2(n1309), .I3(GND_net), 
            .O(n12_adj_4296));
    defparam i3_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1576 (.I0(n1306), .I1(n1308), .I2(n1302), .I3(n10_adj_4295), 
            .O(n16_adj_4297));
    defparam i7_4_lut_adj_1576.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1577 (.I0(n1307), .I1(n16_adj_4297), .I2(n12_adj_4296), 
            .I3(n1301), .O(n1334));
    defparam i8_4_lut_adj_1577.LUT_INIT = 16'hfffe;
    SB_LUT4 i38746_1_lut (.I0(n1433), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45869));
    defparam i38746_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1578 (.I0(n19_adj_4294), .I1(bit_ctr[22]), .I2(n17_adj_4267), 
            .I3(n18_adj_4298), .O(n18_adj_4299));
    defparam i1_4_lut_adj_1578.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1579 (.I0(bit_ctr[25]), .I1(bit_ctr[24]), .I2(bit_ctr[30]), 
            .I3(n18_adj_4299), .O(n30_adj_4265));
    defparam i13_4_lut_adj_1579.LUT_INIT = 16'hfffe;
    SB_LUT4 i22281_2_lut (.I0(bit_ctr[21]), .I1(n1409), .I2(GND_net), 
            .I3(GND_net), .O(n27289));
    defparam i22281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_1580 (.I0(n1405), .I1(n27289), .I2(n1403), .I3(n1406), 
            .O(n16_adj_4300));
    defparam i6_4_lut_adj_1580.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1581 (.I0(n1402), .I1(n1404), .I2(n1400), .I3(n1407), 
            .O(n17_adj_4301));
    defparam i7_4_lut_adj_1581.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1582 (.I0(n17_adj_4301), .I1(n1408), .I2(n16_adj_4300), 
            .I3(n1401), .O(n1433));
    defparam i9_4_lut_adj_1582.LUT_INIT = 16'hfffe;
    SB_LUT4 i38744_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45867));
    defparam i38744_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i18_4_lut_adj_1583 (.I0(n2990), .I1(n2986), .I2(n2996), .I3(n2995), 
            .O(n44_adj_4302));
    defparam i18_4_lut_adj_1583.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1584 (.I0(bit_ctr[5]), .I1(n2992), .I2(n3009), 
            .I3(GND_net), .O(n33_adj_4303));
    defparam i7_3_lut_adj_1584.LUT_INIT = 16'hecec;
    SB_LUT4 i14_4_lut_adj_1585 (.I0(n3008), .I1(n2994), .I2(n2987), .I3(n2988), 
            .O(n40_adj_4304));
    defparam i14_4_lut_adj_1585.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1586 (.I0(n2984), .I1(n2997), .I2(n3001), .I3(n2993), 
            .O(n45_adj_4305));
    defparam i19_4_lut_adj_1586.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1587 (.I0(n2999), .I1(n3006), .I2(n3007), .I3(n3004), 
            .O(n42_adj_4306));
    defparam i16_4_lut_adj_1587.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1588 (.I0(n33_adj_4303), .I1(n44_adj_4302), .I2(n2985), 
            .I3(n2989), .O(n48_adj_4307));
    defparam i22_4_lut_adj_1588.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1589 (.I0(n3003), .I1(n2998), .I2(n2991), .I3(n3000), 
            .O(n41_adj_4308));
    defparam i15_4_lut_adj_1589.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut_adj_1590 (.I0(n45_adj_4305), .I1(n3002), .I2(n40_adj_4304), 
            .I3(n3005), .O(n49));
    defparam i23_4_lut_adj_1590.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut_adj_1591 (.I0(n49), .I1(n41_adj_4308), .I2(n48_adj_4307), 
            .I3(n42_adj_4306), .O(n3017));
    defparam i25_4_lut_adj_1591.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1592 (.I0(n1500), .I1(n1499), .I2(n1505), .I3(n1501), 
            .O(n18_adj_4309));
    defparam i7_4_lut_adj_1592.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1593 (.I0(n1502), .I1(n18_adj_4309), .I2(n1508), 
            .I3(n1503), .O(n20_adj_4310));
    defparam i9_4_lut_adj_1593.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1594 (.I0(n1506), .I1(bit_ctr[20]), .I2(n1509), 
            .I3(GND_net), .O(n15_adj_4311));
    defparam i4_3_lut_adj_1594.LUT_INIT = 16'heaea;
    SB_LUT4 i10_4_lut_adj_1595 (.I0(n15_adj_4311), .I1(n20_adj_4310), .I2(n1504), 
            .I3(n1507), .O(n1532));
    defparam i10_4_lut_adj_1595.LUT_INIT = 16'hfffe;
    SB_LUT4 i38740_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45863));
    defparam i38740_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i38743_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45866));
    defparam i38743_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22369_2_lut (.I0(bit_ctr[3]), .I1(n3209), .I2(GND_net), .I3(GND_net), 
            .O(n27379));
    defparam i22369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20_4_lut_adj_1596 (.I0(n3196), .I1(n3208), .I2(n3199), .I3(n3188), 
            .O(n48_adj_4312));
    defparam i20_4_lut_adj_1596.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1597 (.I0(n3195), .I1(n3202), .I2(n3187), .I3(n3194), 
            .O(n46_adj_4313));
    defparam i18_4_lut_adj_1597.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1598 (.I0(n3200), .I1(n3185), .I2(n3182), .I3(n3192), 
            .O(n47_adj_4314));
    defparam i19_4_lut_adj_1598.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1599 (.I0(n3201), .I1(n3197), .I2(n3190), .I3(n3183), 
            .O(n45_adj_4315));
    defparam i17_4_lut_adj_1599.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1600 (.I0(n3184), .I1(n3205), .I2(n3206), .I3(n3186), 
            .O(n44_adj_4316));
    defparam i16_4_lut_adj_1600.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1601 (.I0(n3198), .I1(n3193), .I2(n3189), .I3(n27379), 
            .O(n43_adj_4317));
    defparam i15_4_lut_adj_1601.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1602 (.I0(n45_adj_4315), .I1(n47_adj_4314), .I2(n46_adj_4313), 
            .I3(n48_adj_4312), .O(n54));
    defparam i26_4_lut_adj_1602.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1603 (.I0(n3191), .I1(n3207), .I2(n3204), .I3(n3203), 
            .O(n49_adj_4318));
    defparam i21_4_lut_adj_1603.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n49_adj_4318), .I1(n54), .I2(n43_adj_4317), 
            .I3(n44_adj_4316), .O(n27449));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 color_bit_I_0_i19_3_lut (.I0(\color[20] ), .I1(\color[21] ), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n19_adj_4319));   // verilog/neopixel.v(22[26:36])
    defparam color_bit_I_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35953_2_lut (.I0(\color[17] ), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(GND_net), .O(n42814));
    defparam i35953_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i48_3_lut (.I0(n27449), .I1(bit_ctr[3]), .I2(n3209), .I3(GND_net), 
            .O(n25_adj_4320));
    defparam i48_3_lut.LUT_INIT = 16'h1818;
    SB_LUT4 i2_4_lut_adj_1604 (.I0(n42814), .I1(bit_ctr[1]), .I2(n19_adj_4319), 
            .I3(bit_ctr[2]), .O(n7_adj_4321));
    defparam i2_4_lut_adj_1604.LUT_INIT = 16'h3022;
    SB_LUT4 i4_4_lut (.I0(n7_adj_4321), .I1(n25_adj_4320), .I2(n27164), 
            .I3(n33679), .O(state_3__N_362[0]));
    defparam i4_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 mux_654_Mux_0_i3_3_lut_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_570 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_654_Mux_0_i3_3_lut_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 i8_4_lut_adj_1605 (.I0(n1608), .I1(n1606), .I2(n1604), .I3(n1603), 
            .O(n20_adj_4322));
    defparam i8_4_lut_adj_1605.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1606 (.I0(bit_ctr[19]), .I1(n1602), .I2(n1609), 
            .I3(GND_net), .O(n13_adj_4323));
    defparam i1_3_lut_adj_1606.LUT_INIT = 16'hecec;
    SB_LUT4 i6_2_lut (.I0(n1598), .I1(n1600), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4324));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1607 (.I0(n13_adj_4323), .I1(n20_adj_4322), .I2(n1605), 
            .I3(n1599), .O(n22_adj_4325));
    defparam i10_4_lut_adj_1607.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1608 (.I0(n1601), .I1(n22_adj_4325), .I2(n18_adj_4324), 
            .I3(n1607), .O(n1631));
    defparam i11_4_lut_adj_1608.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_2_lut (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n37374));
    defparam i1_3_lut_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i38741_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45864));
    defparam i38741_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_4_lut (.I0(n32476), .I1(n17064), .I2(start), .I3(\neo_pixel_transmitter.done ), 
            .O(n1105));   // verilog/neopixel.v(79[18] 99[12])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hf1ff;
    SB_LUT4 i1_3_lut_4_lut (.I0(n17064), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(n4_adj_4216), .O(n17196));   // verilog/neopixel.v(52[18] 72[12])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hcfdf;
    SB_LUT4 i3_4_lut_4_lut (.I0(n38037), .I1(n15780), .I2(n807), .I3(bit_ctr[27]), 
            .O(n838));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 i7_4_lut_adj_1609 (.I0(bit_ctr[19]), .I1(bit_ctr[15]), .I2(bit_ctr[27]), 
            .I3(bit_ctr[6]), .O(n18_adj_4298));
    defparam i7_4_lut_adj_1609.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i538_3_lut_4_lut_3_lut (.I0(n708), .I1(n7476), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i538_3_lut_4_lut_3_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n708), .I1(n7476), .I2(bit_ctr[28]), 
            .I3(GND_net), .O(n15780));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 i1_3_lut_4_lut_3_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(bit_ctr[29]), 
            .I3(GND_net), .O(n32958));   // verilog/neopixel.v(22[26:36])
    defparam i1_3_lut_4_lut_3_lut.LUT_INIT = 16'h9494;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis lattice_noprune=1, syn_instantiated=1, LSE_LINE_FILE_ID=49, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=35, LSE_RLINE=38, syn_preserve=0 */ ;   // verilog/TinyFPGA_B.v(35[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module coms
//

module coms (rx_data, PWMLimit, clk32MHz, GND_net, n19434, setpoint, 
            n19435, n19436, n19437, n19438, n19439, n19440, n19427, 
            n19428, n19429, n19430, n19431, control_mode, VCC_net, 
            n19448, n19449, n19446, n19447, n19444, n19445, n19441, 
            n19442, n19443, n19432, n19433, n46050, n19145, \data_out_frame[20] , 
            n19144, n19143, n19142, n19141, n19140, n19139, n19138, 
            n19137, \data_out_frame[19] , n19136, n19135, n19134, 
            n19133, n19132, n19131, n19130, n19129, \data_out_frame[18] , 
            n19128, n19127, n19126, n17199, \data_out_frame[5] , \data_out_frame[7] , 
            \FRAME_MATCHER.state[3] , \FRAME_MATCHER.state[0] , n63, n17268, 
            n2857, n38098, n17200, n17202, n19125, n19124, n19123, 
            n19122, \data_out_frame[8] , \data_out_frame[11] , n19121, 
            \data_out_frame[17] , n19120, n19119, n19118, n19117, 
            n19116, n19115, n19114, n19113, \data_out_frame[16] , 
            n4661, n19112, n19111, n19110, n4659, \data_out_frame[12] , 
            n19109, n19108, n19107, n19106, n19105, \data_out_frame[15] , 
            n19104, n18435, n6119, ID0, n19103, n19102, rx_data_ready, 
            ID2, \data_out_frame[14] , n19101, n19272, \data_in_frame[15] , 
            n19271, n19270, n19100, n19099, n19098, n19097, \data_out_frame[13] , 
            \data_out_frame[6] , n19096, n19095, \data_out_frame[4][0] , 
            n19094, \data_out_frame[4][2] , \data_out_frame[10] , \data_out_frame[9] , 
            n19093, n19092, n19091, n19090, n19089, n19088, n19087, 
            n19086, n19085, n19084, n19083, n19082, n19081, n19080, 
            n19079, n19078, n19077, n19076, n19075, n19074, n19073, 
            n19072, n19071, n19070, n19069, n19068, n19067, n19066, 
            n19065, n19269, n19064, n19268, n19063, n19062, n19061, 
            n19060, n19059, n19058, n19057, n19056, n19055, n19054, 
            n19053, n19052, n19051, n19050, n19049, n19048, n19047, 
            n19046, n19045, n19044, n19043, n19267, n19042, n19041, 
            n19040, n19039, n19038, n19266, n19037, n19036, n19035, 
            n19034, n19033, n19032, n19265, n19031, n19030, n19029, 
            n19028, n19027, ID1, n14536, n4660, n19026, n19025, 
            n19024, n19023, n19022, n4673, n19021, n19020, n4672, 
            n4671, n4670, n4669, n4668, n19019, n19018, n19017, 
            n19014, n19013, \data_out_frame[0][4] , n19012, \data_out_frame[0][3] , 
            n19011, \data_in[3] , n19010, n19009, n19008, n19007, 
            n19006, n19005, n19004, n19003, \data_in[2] , n19002, 
            n19001, n19000, n18999, n18998, n18997, n18996, n18995, 
            \data_in[1] , n18994, n18993, n18992, n18991, n18990, 
            n18989, n18988, n18987, \data_in[0] , n18986, n18985, 
            n18984, n18983, n18982, n18981, \Ki[7] , \Ki[6] , \Ki[5] , 
            \Ki[4] , \Ki[3] , \Ki[2] , \Ki[1] , \Kp[7] , \Kp[6] , 
            \Kp[5] , \Kp[4] , \Kp[3] , \Kp[2] , \Kp[1] , gearBoxRatio, 
            IntegralLimit, \Kp[0] , \Ki[0] , \data_in_frame[7] , n37368, 
            n17264, n37348, n18829, n19208, n3761, n740, n19207, 
            n19206, n19205, n19204, n2664, n36597, n19203, n18798, 
            LED_c, n20639, n5, n46559, n5_adj_3, n19202, n19201, 
            n37376, n40, n4666, n4665, n4676, n4675, n4674, n4678, 
            n4677, n4680, n4679, n4682, n4681, n39863, n4667, 
            n4664, n4663, n4662, n18758, n18755, n18752, n18749, 
            n19426, r_SM_Main, n18746, n18767, n18764, n18761, n18744, 
            n18747, \r_SM_Main_2__N_3320[1] , n18750, n18753, n18756, 
            n18759, n18762, n18765, n18896, n18898, n18816, n18815, 
            tx_active, n18814, tx_o, n45935, tx_enable, n18402, 
            n12501, n18897, n36985, \r_Clock_Count[2] , n36987, \r_Clock_Count[3] , 
            n36989, \r_Clock_Count[4] , n36919, \r_Clock_Count[5] , 
            n36743, \r_Clock_Count[6] , n36695, \r_Clock_Count[7] , 
            n36983, \r_Clock_Count[1] , n18780, r_Bit_Index, n18777, 
            n19419, n27445, \r_SM_Main[1]_adj_4 , n95, n16, \r_SM_Main[2]_adj_5 , 
            r_Rx_Data, PIN_13_N_105, n37215, n37220, n37217, n37216, 
            n37218, n37219, n37214, n18943, n18806, n18793, n18786, 
            n18785, n18784, n18783, n18782, n18781, n42920, n20874, 
            n42919, n17255, n4, n26349, n4_adj_6, n4_adj_7, n17250, 
            n4926, n18467, n20896, n18602) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [7:0]rx_data;
    output [23:0]PWMLimit;
    input clk32MHz;
    input GND_net;
    input n19434;
    output [23:0]setpoint;
    input n19435;
    input n19436;
    input n19437;
    input n19438;
    input n19439;
    input n19440;
    input n19427;
    input n19428;
    input n19429;
    input n19430;
    input n19431;
    output [7:0]control_mode;
    input VCC_net;
    input n19448;
    input n19449;
    input n19446;
    input n19447;
    input n19444;
    input n19445;
    input n19441;
    input n19442;
    input n19443;
    input n19432;
    input n19433;
    input n46050;
    input n19145;
    output [7:0]\data_out_frame[20] ;
    input n19144;
    input n19143;
    input n19142;
    input n19141;
    input n19140;
    input n19139;
    input n19138;
    input n19137;
    output [7:0]\data_out_frame[19] ;
    input n19136;
    input n19135;
    input n19134;
    input n19133;
    input n19132;
    input n19131;
    input n19130;
    input n19129;
    output [7:0]\data_out_frame[18] ;
    input n19128;
    input n19127;
    input n19126;
    output n17199;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[7] ;
    output \FRAME_MATCHER.state[3] ;
    output \FRAME_MATCHER.state[0] ;
    output n63;
    output n17268;
    output n2857;
    output n38098;
    output n17200;
    output n17202;
    input n19125;
    input n19124;
    input n19123;
    input n19122;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[11] ;
    input n19121;
    output [7:0]\data_out_frame[17] ;
    input n19120;
    input n19119;
    input n19118;
    input n19117;
    input n19116;
    input n19115;
    input n19114;
    input n19113;
    output [7:0]\data_out_frame[16] ;
    output n4661;
    input n19112;
    input n19111;
    input n19110;
    output n4659;
    output [7:0]\data_out_frame[12] ;
    input n19109;
    input n19108;
    input n19107;
    input n19106;
    input n19105;
    output [7:0]\data_out_frame[15] ;
    input n19104;
    output n18435;
    output n6119;
    input ID0;
    input n19103;
    input n19102;
    output rx_data_ready;
    input ID2;
    output [7:0]\data_out_frame[14] ;
    input n19101;
    input n19272;
    output [7:0]\data_in_frame[15] ;
    input n19271;
    input n19270;
    input n19100;
    input n19099;
    input n19098;
    input n19097;
    output [7:0]\data_out_frame[13] ;
    output [7:0]\data_out_frame[6] ;
    input n19096;
    input n19095;
    output \data_out_frame[4][0] ;
    input n19094;
    output \data_out_frame[4][2] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[9] ;
    input n19093;
    input n19092;
    input n19091;
    input n19090;
    input n19089;
    input n19088;
    input n19087;
    input n19086;
    input n19085;
    input n19084;
    input n19083;
    input n19082;
    input n19081;
    input n19080;
    input n19079;
    input n19078;
    input n19077;
    input n19076;
    input n19075;
    input n19074;
    input n19073;
    input n19072;
    input n19071;
    input n19070;
    input n19069;
    input n19068;
    input n19067;
    input n19066;
    input n19065;
    input n19269;
    input n19064;
    input n19268;
    input n19063;
    input n19062;
    input n19061;
    input n19060;
    input n19059;
    input n19058;
    input n19057;
    input n19056;
    input n19055;
    input n19054;
    input n19053;
    input n19052;
    input n19051;
    input n19050;
    input n19049;
    input n19048;
    input n19047;
    input n19046;
    input n19045;
    input n19044;
    input n19043;
    input n19267;
    input n19042;
    input n19041;
    input n19040;
    input n19039;
    input n19038;
    input n19266;
    input n19037;
    input n19036;
    input n19035;
    input n19034;
    input n19033;
    input n19032;
    input n19265;
    input n19031;
    input n19030;
    input n19029;
    input n19028;
    input n19027;
    input ID1;
    output n14536;
    output n4660;
    input n19026;
    input n19025;
    input n19024;
    input n19023;
    input n19022;
    output n4673;
    input n19021;
    input n19020;
    output n4672;
    output n4671;
    output n4670;
    output n4669;
    output n4668;
    input n19019;
    input n19018;
    input n19017;
    input n19014;
    input n19013;
    output \data_out_frame[0][4] ;
    input n19012;
    output \data_out_frame[0][3] ;
    input n19011;
    output [7:0]\data_in[3] ;
    input n19010;
    input n19009;
    input n19008;
    input n19007;
    input n19006;
    input n19005;
    input n19004;
    input n19003;
    output [7:0]\data_in[2] ;
    input n19002;
    input n19001;
    input n19000;
    input n18999;
    input n18998;
    input n18997;
    input n18996;
    input n18995;
    output [7:0]\data_in[1] ;
    input n18994;
    input n18993;
    input n18992;
    input n18991;
    input n18990;
    input n18989;
    input n18988;
    input n18987;
    output [7:0]\data_in[0] ;
    input n18986;
    input n18985;
    input n18984;
    input n18983;
    input n18982;
    input n18981;
    output \Ki[7] ;
    output \Ki[6] ;
    output \Ki[5] ;
    output \Ki[4] ;
    output \Ki[3] ;
    output \Ki[2] ;
    output \Ki[1] ;
    output \Kp[7] ;
    output \Kp[6] ;
    output \Kp[5] ;
    output \Kp[4] ;
    output \Kp[3] ;
    output \Kp[2] ;
    output \Kp[1] ;
    output [23:0]gearBoxRatio;
    output [23:0]IntegralLimit;
    output \Kp[0] ;
    output \Ki[0] ;
    output [7:0]\data_in_frame[7] ;
    output n37368;
    output n17264;
    output n37348;
    input n18829;
    input n19208;
    output n3761;
    output n740;
    input n19207;
    input n19206;
    input n19205;
    input n19204;
    output n2664;
    input n36597;
    input n19203;
    input n18798;
    output LED_c;
    output n20639;
    output n5;
    output n46559;
    output n5_adj_3;
    input n19202;
    input n19201;
    output n37376;
    output n40;
    output n4666;
    output n4665;
    output n4676;
    output n4675;
    output n4674;
    output n4678;
    output n4677;
    output n4680;
    output n4679;
    output n4682;
    output n4681;
    output n39863;
    output n4667;
    output n4664;
    output n4663;
    output n4662;
    input n18758;
    input n18755;
    input n18752;
    input n18749;
    input n19426;
    output [2:0]r_SM_Main;
    input n18746;
    input n18767;
    input n18764;
    input n18761;
    output n18744;
    output n18747;
    output \r_SM_Main_2__N_3320[1] ;
    output n18750;
    output n18753;
    output n18756;
    output n18759;
    output n18762;
    output n18765;
    output n18896;
    input n18898;
    input n18816;
    input n18815;
    output tx_active;
    input n18814;
    output tx_o;
    output n45935;
    output tx_enable;
    output n18402;
    output n12501;
    output n18897;
    input n36985;
    output \r_Clock_Count[2] ;
    input n36987;
    output \r_Clock_Count[3] ;
    input n36989;
    output \r_Clock_Count[4] ;
    input n36919;
    output \r_Clock_Count[5] ;
    input n36743;
    output \r_Clock_Count[6] ;
    input n36695;
    output \r_Clock_Count[7] ;
    input n36983;
    output \r_Clock_Count[1] ;
    input n18780;
    output [2:0]r_Bit_Index;
    input n18777;
    input n19419;
    input n27445;
    output \r_SM_Main[1]_adj_4 ;
    output n95;
    input n16;
    output \r_SM_Main[2]_adj_5 ;
    output r_Rx_Data;
    input PIN_13_N_105;
    output n37215;
    output n37220;
    output n37217;
    output n37216;
    output n37218;
    output n37219;
    output n37214;
    input n18943;
    input n18806;
    input n18793;
    input n18786;
    input n18785;
    input n18784;
    input n18783;
    input n18782;
    input n18781;
    output n42920;
    output n20874;
    output n42919;
    output n17255;
    output n4;
    output n26349;
    output n4_adj_6;
    output n4_adj_7;
    output n17250;
    output n4926;
    output n18467;
    output n20896;
    output n18602;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire LED_c /* synthesis SET_AS_NETWORK=LED_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(4[10:13])
    
    wire n8, n37361;
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(94[12:25])
    
    wire n19163, n19351, n19174;
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(94[12:25])
    
    wire n19294;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(94[12:25])
    
    wire n19293, n19292, n19291, n19290, n19289, n19350, n19349, 
        n19288;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(94[12:25])
    
    wire n19287, n19286, n19285, n19284, n19283, n19282, n19173, 
        n2;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(113[11:12])
    
    wire n30318, n1972, n30319, n19172, n2_adj_3902, n3, n19281, 
        n2_adj_3903, n30317, n19280;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(94[12:25])
    
    wire n19279, n19171, n19170, n2_adj_3904, n30316, n2_adj_3905, 
        n30315, n19169, n19168, n19167, n19278, n19277, n19276, 
        n19275, n19274, n19198;
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(94[12:25])
    
    wire n19197, n19348, n19196, n19347, n19195, n19194;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(94[12:25])
    
    wire n6, n19193, n19346, n19166, n19345, n19192;
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(94[12:25])
    
    wire n19344, n19343, n19342, n19341, n19340, n19339, n19338, 
        n19337, n19336, n19335, n19334, n19333, n19332, n19331, 
        n19330, n19329, n19328, n19327, n19326, n19456;
    wire [7:0]\data_out_frame[0] ;   // verilog/coms.v(95[12:26])
    
    wire n19325;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(100[12:33])
    
    wire n19324, n19453, n20482, n19321, n19320, n19319, n19318, 
        n19354, n19317, n19316, n19315, n19314, n19313, n19312;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(94[12:25])
    
    wire n19311, n19310, n19191, n19309, n19190;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(110[11:16])
    
    wire n19308, n19307, n19306, n19305, n19304;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(94[12:25])
    
    wire n19303, n19302, n19301, n19300, n19299, n19298, n19297, 
        n19296, n19295, n19165, n19164, n19162, n19161, n19160;
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(94[12:25])
    
    wire n19159, n19158, n19157, n19156, n19155, n19154, n19153, 
        n19152;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(94[12:25])
    
    wire n19151, n19150, n19149, n19148, n19147, n19236;
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(94[12:25])
    
    wire n19235, n19234, n19233, n19146, n19232;
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(94[12:25])
    
    wire n19231, n19230, n19241;
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(94[12:25])
    
    wire n37401, n18140, n17542, n38588, n19189, n19229, n19188, 
        n19187, n19228, n19227, n19226, n19225, n19186, n19185, 
        n19184;
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(94[12:25])
    
    wire n19183, n19182, n19181, n8_adj_3906, n37953, n10, n19180, 
        n19179, n19178, n19177, n19176, n30320, n8_adj_3907, n37342;
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(94[12:25])
    
    wire n19209, n17266, n14748, n14721, n9, n19210, n37588, n37520, 
        n17988, n19211, n19212, n200, n322, n326, n6_adj_3908, 
        n19213, n17170;
    wire [31:0]\FRAME_MATCHER.state_31__N_2492 ;
    
    wire n17025, n36609, n324, n301, n36589, n31, Kp_23__N_1745, 
        tx_transmit_N_3215;
    wire [0:0]n3086;
    
    wire n63_c, n63_adj_3909, n20661, n19214;
    wire [31:0]n93;
    
    wire n5_c, n4658, n6_adj_3911, n19215;
    wire [31:0]\FRAME_MATCHER.state_31__N_2460 ;
    
    wire n46228, n19216, n40932, n40931;
    wire [7:0]tx_data;   // verilog/coms.v(103[13:20])
    
    wire n37839, n17979, n19224;
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(94[12:25])
    
    wire n19223, n40929, n40928, n40926, n40925, n40923, n40922, 
        n19222, n8_adj_3912;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(94[12:25])
    
    wire n19257, n19258, n19259, n19260, n19261, n19262, n19263, 
        n19264, n37440, n37786, n37735, n33079, n33882, n17664, 
        n38713, n18200, n37604, n37549, n2_adj_3913, n30314, n37738, 
        n37723, n38953, n2_adj_3914, n30313, n33902, n32998, n17671, 
        n6_adj_3915, n37801, n37640, n33047, n37666, n37467, n12, 
        \FRAME_MATCHER.rx_data_ready_prev , n33016, n37482, n37869, 
        n37872, n10_adj_3916, n38644, n18850, n2_adj_3917, n30312, 
        n37514, n37386, n12_adj_3918, n18381, n10308;
    wire [7:0]n2236;
    
    wire n33049, n6_adj_3919, n38639, n33941, n37720, n37721, n37744, 
        n10_adj_3920, n37673, n4_c, n39012, n37479, n19221, n19273, 
        n37508, n37701, n32950, n10_adj_3921, n37814, n32979, n1595, 
        n14, n39220, n1185, n33822, n17325, n37530, n17782, n12_adj_3922, 
        n17626, n37890, n37647, n37962, n10_adj_3923, n33067, n16_c, 
        n37380, n37911, n1642, n17, n38802, n32717, n37717, n17969, 
        n37707, n17746, n17183, n36679, n33880, n17778, n33893, 
        n10_adj_3924, n37407, n6_adj_3925, n16772, n19352, n6_adj_3926, 
        n37613, n37807, n32719, n19238, n6_adj_3927, n37539, n17963, 
        n37504, n37578, n33875, n19237, n2_adj_3928, n30311, n2_adj_3929, 
        n30310, n33845, n42985, n40910;
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(95[12:26])
    
    wire n19, n19220, n37863, n37492, n39208;
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(95[12:26])
    
    wire n40934, n40911, n37601, n18143, n17916, n17638, n18147, 
        n10_adj_3930, n37422, n40909, n46031, n45881, n44499, n39027, 
        n33815, n37561, n37884, n10_adj_3931, n37413, n45941, n40935, 
        n37634, n40912, n44728, n37486, n37763, n10_adj_3932, n8_adj_3933, 
        n37354, n37552, n18209, n54, n37473, n37395, n52, n53, 
        n51, n37935, n48, n37804, n37419, n50, n37652, n18079, 
        n49, n60, n37501, n1559, n55, n16906, n32972, n37704, 
        n39565, n37575, n18, n37404, n20, n15, n37687, n18119, 
        n17404, n37517, n33035, n38540, n2_adj_3934, n30309, n17860, 
        n17422, n12_adj_3935, n17365, n10_adj_3936;
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(94[12:25])
    
    wire n19249, n37572, n17817, n37655, n37875, n17844, n37992, 
        n6_adj_3937, n25, n37643, n38695, n37866, n19_adj_3938, 
        n30, n19250, n17764, n37923, n28, n37792, n29, n37941, 
        n27, n37766, n12_adj_3939, n16787, n19251, n37416, n16915, 
        n19252, n19253, n6_adj_3940, n2_adj_3941, n30308, n37757, 
        n10_adj_3942, n19254, n1119, n6_adj_3943, n6_adj_3944, n19255, 
        n4_adj_3945, n37741, n38435, n37658, n19256, n52_adj_3946, 
        n8_adj_3947, n37965, n50_adj_3948, n17330, n51_adj_3949, n49_adj_3950, 
        n37977, n46, n2_adj_3951, n30307, n48_adj_3952, n32716, 
        n47, n58, n37665, n53_adj_3953, n2_adj_3954, n30306, n39387, 
        n37798, n16_adj_3955, n17_adj_3956, n16817, n38620, n10_adj_3957, 
        n33008, n10_adj_3958, n2_adj_3959, n30305, n38514, n2_adj_3960, 
        n30304, n19219;
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(95[12:26])
    
    wire n19016, n37830, n37555, n17833, n39798, n17418, n19218, 
        n17725, n17742, n6_adj_3961, n18031, n14_adj_3962, n37810, 
        n33891, n37944, n15_adj_3963, n37827, n37496, n39794, n16_adj_3964, 
        n17_adj_3965, n18073, Kp_23__N_893, n11, n37817, n37899, 
        n15612, n17687, n2_adj_3966, n30303, n17648, n6_adj_3967, 
        n37591, n1287, n37920, n15_adj_3968, n18219, n14_adj_3969, 
        n12_adj_3970, n2_adj_3971, n30302, n164, n18292, n42885, 
        n30339, n30338, n32986, n17821, n37750, n37914, n18082, 
        n37677, n10_adj_3972, n6_adj_3973, n42882, n30337, n37842, 
        n18_adj_3974, n16_adj_3975, n20_adj_3976, n6_adj_3977, n38809, 
        n14_adj_3978, n10_adj_3979, n6121, n18436, n42884, n30336, 
        n18980, n18979, n18978, n18977, n18976, n18975, n18974, 
        n18973, n18972, n18971, n18970, n18969, n18968, n18967, 
        n18966, n18965, n18964, n18963, n18962, n18961, n18960, 
        n18959, n18958, n18957, n18956, n18955, n18954, n18953, 
        n18952, n18951, n18950, n18949, n18948, n18947, n18946, 
        n4_adj_3980, n18945, n18944, n19199, n18937, n18936, Kp_23__N_718, 
        n63_adj_3981, n18664, n19353, n18935, n18934, n18933, n18795, 
        n18796, n37545, n37610, n38719, n18932, n18931, n18930, 
        n18929, n18797, n18800, n42881, n30335, n18801, n18915, 
        n18928, n18927, n18926, n17482, n18925, n18916, n18924, 
        n18923, n18922, n18917, n18921, n18920, n18919, n18918, 
        n18914, n18913, n36219, n36213, n18910, n37860, n19200, 
        n42974, n30334, n27114, n10_adj_3982, n17031, n17045, n33852, 
        n37476, n18122, n17874, Kp_23__N_1353, Kp_23__N_1372, n37881, 
        n18155, n37795, n17500, n37893, n37848, n37950, n37436, 
        n14_adj_3983, n10_adj_3984, n37594, n17445, n37769, n37980, 
        n37845, n37947, n20_adj_3985, n37430, n19_adj_3986, n17696, 
        n17492, n21, n17222, n18_adj_3987, n20_adj_3988, n5_adj_3989, 
        n37929, Kp_23__N_1083, n37783, n37536, n37905, n17449, n37780, 
        n6_adj_3990, n37690, n37729, n37908, n10_adj_3991, n18006, 
        n37747, n14_adj_3992, n10_adj_3993, n37878, n17425, n15_adj_3994, 
        n14_adj_3995, n37597, n37661, n37956, n10_adj_3996, n37463, 
        Kp_23__N_858, n37526, n3_adj_3997, n26, n24, n25_adj_3998, 
        n37631, n23, n37710, n33070, n37983, n33854, n33864, n7, 
        n37989, n14_adj_3999, n10_adj_4000, n39322, n37616, n48_adj_4001, 
        n33886, n54_adj_4002, n37773, n37693, n52_adj_4003, n37470, 
        n53_adj_4004, n37887, n51_adj_4005, n37714, n37533, n50_adj_4006, 
        Kp_23__N_760, n49_adj_4007, n60_adj_4008, n5_adj_4009, n37959, 
        n37433, n55_adj_4010, n39467, n37917, n42, n31_adj_4011, 
        Kp_23__N_1406, n28_adj_4012, n37968, n26_adj_4013, n37974, 
        n37443, n27_adj_4014, n25_adj_4015, n26_adj_4016, n39193, 
        n37820, n28_adj_4017, n40_c, n37726, n46_adj_4018, n44, 
        n45, n37760, n43, n37669, n37383, n15_adj_4019, n6_adj_4020, 
        n37926, n17827, n37902, n33843, n18228, n12_adj_4021, n18091, 
        n17379, n37622, n10_adj_4022, n37511, n17863, n37564, n37567, 
        n37851, n37776, n12_adj_4023, n17559, n17055, n8_adj_4024, 
        n12_adj_4025, n38781, n37939, n17_adj_4026, n16_adj_4027, 
        n39117, n22, n40829, n17167, n16_adj_4028, n3_adj_4029, 
        n3_adj_4030, n17_adj_4031, n3_adj_4032, n3_adj_4033, n3_adj_4034, 
        n3_adj_4035, n3_adj_4036, n3_adj_4037, n3_adj_4038, n3_adj_4039, 
        n3_adj_4040, n3_adj_4041, n3_adj_4042, n3_adj_4043, n3_adj_4044, 
        n3_adj_4045, n3_adj_4046, n2_adj_4047, n3_adj_4048, n2_adj_4049, 
        n3_adj_4050, n2_adj_4051, n3_adj_4052, n2_adj_4053, n3_adj_4054, 
        n2_adj_4055, n3_adj_4056, n2_adj_4057, n3_adj_4058, n2_adj_4059, 
        n3_adj_4060, n2_adj_4061, n3_adj_4062, n2_adj_4063, n3_adj_4064, 
        n2_adj_4065, n3_adj_4066, n2_adj_4067, n3_adj_4068, n2_adj_4069, 
        n3_adj_4070, n2_adj_4071, n3_adj_4072, n2_adj_4073, n3_adj_4074, 
        n38745, n46028, n38922, n38629, n38857, n37802, n37826, 
        n37825, n37551, n17597, n39432, n36585, n36783, n36787, 
        n36599, n36791, n36601, n36795, n36659, n36799, n36657, 
        n36803, n36655, n36811, n36651, n36815, n36649, n36819, 
        n36647, n36823, n36645, n36827, n36643, n7_adj_4075, n8_adj_4076, 
        n36831, n36603, n7_adj_4077, n8_adj_4078, n7_adj_4079, n8_adj_4080, 
        n36751, n36579, n7_adj_4081, n36683, n36807, n36653, n36763, 
        n36641, n7_adj_4082, n8_adj_4083, n7_adj_4084, n36639, n36767, 
        n36693, n36771, n36637, n7_adj_4085, n8_adj_4086, n36775, 
        n36635, n7_adj_4087, n8_adj_4088, n36779, n8_adj_4089, n7_adj_4090, 
        n19217, n46022, n46025, n12_adj_4091, n46016, n46019, n37754, 
        n46010, n46013, n37392, n46004, n46007, n37896, n45998, 
        n46001, n37698, n18_adj_4092, n45992, n45995, n16_adj_4093, 
        n45986, n45989, n42973, n30333, n17247, n16_adj_4094, n17_adj_4095, 
        n30321, n8_adj_4096, Kp_23__N_820, n20_adj_4097, n45980, n43083;
    wire [2:0]r_SM_Main_2__N_3323;
    
    wire n38178, n19240, n17900, n7_adj_4098, n28_adj_4099, n39620, 
        n7_adj_4100, n8_adj_4101, n39166, n17208, n26492, n40790, 
        n26_adj_4102, n30_adj_4103, n17_adj_4104, Kp_23__N_1433, n31_adj_4105, 
        n27441, n20_adj_4106, n6_adj_4107, n33677, n30_adj_4108, n34, 
        n32, n33, n4_adj_4109, n31_adj_4110, n17265, n26317, n38092, 
        n17201, n30332, n17636, n26_adj_4111, n37607, n37489, n8_adj_4112, 
        n42_adj_4113, n40_adj_4114, n41, n17263, n39, n38, n37, 
        n48_adj_4115, n43_adj_4116, n40827, n30331, n18799, n45983, 
        n9_adj_4117, n30330, n38165, n22_adj_4118, n27_adj_4119, n25_adj_4120, 
        n19175, n37209, n10_adj_4121, n14_adj_4122, n10_adj_4123, 
        n40809, n21_adj_4124, n37398, n20_adj_4125, n37378, n30329, 
        n30328, n24_adj_4126, n33828, n30327, n30326, n30325, n30324, 
        n19248, n19247, n19246, n30323, n40965, n40963, n40918, 
        n40956, n40954, n40915, n19245, n19239, n30322, n47_adj_4129, 
        n37854, n17853, n37619, n19244, n19243, n19242, n6_adj_4130, 
        n45974, n45977, n37986, n37971, n14_adj_4131, n45968, n45971, 
        n10_adj_4132, n37523, n45962, n44437, n45956, n40996, n45950, 
        n45953, n10_adj_4133, n16_adj_4134, n45944, n45947, n18295, 
        n15_adj_4135, n45938, n45926, n40946, n40945, n45929, n12503, 
        Kp_23__N_839, n33430, n12_adj_4136, n6_adj_4137, n37699, n18001, 
        n16726, n17928, n37732, n10_adj_4138, n17840, n33850, n37628, 
        n12_adj_4139, n37932, n37410, Kp_23__N_1562, n38088, n10_adj_4140, 
        n37789, n12_adj_4141, n18023, n32943, n4_adj_4142, n10_adj_4143, 
        n6_adj_4144, n37450, n16859, n32982, n37857, n10_adj_4146, 
        n16_adj_4147, n17_adj_4148, n42810, n19_adj_4149, n16_adj_4150, 
        n17_adj_4151, n42811, n19_adj_4152, n18_adj_4153, n16_adj_4154, 
        n17_adj_4155, n42818, n19_adj_4156, n16_adj_4157, n17_adj_4158, 
        n42987, n19_adj_4159, n16_adj_4160, n17_adj_4161, n42819, 
        n19_adj_4162, n5_adj_4163, n22_adj_4164, n14340, n33295, n33087, 
        n16_adj_4165, n8_adj_4166, n26281, n45920, n8_adj_4167, n20_adj_4168, 
        n40802, n45923, n27475, n6_adj_4169, n20642, n40815, n40813, 
        n13, Kp_23__N_1746, n45914, n39564, n26_adj_4170, n17_adj_4171, 
        n28_adj_4172, n29_adj_4173, n45917, n10_adj_4174, n45908, 
        n45911, n45902, n45905, n14_adj_4175, n44_adj_4176, n43081;
    wire [0:0]n3139;
    
    wire n45896, n45899, n13_adj_4177, n43367, n5_adj_4178, n40930, 
        n43362, n5_adj_4179, n40927, n43357, n5_adj_4180, n40924, 
        n42914, n6_adj_4181, n5_adj_4182, n40921, n42930, n40964, 
        n19_adj_4183, n40940, n45893, n44489, n45890, n40941, n44734, 
        n42938, n40955, n19_adj_4184, n40937, n45887, n44491, n40938, 
        n44732, n45884, n45878;
    
    SB_LUT4 i14131_3_lut_4_lut (.I0(n8), .I1(n37361), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n19163));
    defparam i14131_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n19351));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n19174));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n19294));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n19293));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n19292));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n19291));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n19290));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n19289));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n19350));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n19349));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n19288));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n19287));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n19286));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n19285));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n19284));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n19283));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n19282));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n19173));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_19_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n30318), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_19 (.CI(n30318), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n30319));
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n19172));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2_adj_3902), .S(n3));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n19281));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_18_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n30317), .O(n2_adj_3903)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_18_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n19280));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n19279));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n19171));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_18 (.CI(n30317), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n30318));
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n19170));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_17_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n30316), .O(n2_adj_3904)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_17 (.CI(n30316), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n30317));
    SB_LUT4 add_44_16_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n30315), .O(n2_adj_3905)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_16_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n19169));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n19168));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n19167));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n19278));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n19277));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n19276));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n19275));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n19274));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n19198));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n19197));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n19348));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n19196));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n19347));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n19195));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n19194));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut (.I0(\data_in_frame[21] [6]), .I1(\data_in_frame[17] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n19193));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n19346));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n19166));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n19345));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n19192));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n19344));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n19343));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n19342));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n19341));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n19340));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n19339));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n19338));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n19337));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n19336));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .D(n19434));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .D(n19435));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .D(n19436));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .D(n19437));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .D(n19438));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .D(n19439));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .D(n19440));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n19335));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .D(n19427));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .D(n19428));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .D(n19429));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .D(n19430));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .D(n19431));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n19334));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n19333));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n19332));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n19331));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n19330));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n19329));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n19328));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n19327));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n19326));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i1 (.Q(\data_out_frame[0] [0]), .C(clk32MHz), 
            .E(VCC_net), .D(n19456));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(clk32MHz), 
           .D(n19325));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk32MHz), 
           .D(n19324));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE byte_transmit_counter_i0_i0 (.Q(byte_transmit_counter[0]), .C(clk32MHz), 
            .E(VCC_net), .D(n19453));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(clk32MHz), 
           .D(n20482));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .D(n19448));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .D(n19449));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n19321));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .D(n19446));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .D(n19447));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n19320));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .D(n19444));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .D(n19445));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .D(n19441));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .D(n19442));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .D(n19443));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .D(n19432));   // verilog/coms.v(126[12] 289[6])
    SB_DFF setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .D(n19433));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n19319));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n19318));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n19354));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n19317));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n19316));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n19315));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n19314));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n19313));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n19312));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n19311));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n19310));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n19191));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n19309));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n19190));   // verilog/coms.v(126[12] 289[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk32MHz), 
           .D(n46050));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n19308));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n19307));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n19306));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n19305));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n19304));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n19303));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n19302));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n19301));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n19300));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n19299));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n19298));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n19297));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n19296));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n19295));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n19165));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n19164));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n19163));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n19162));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n19161));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n19160));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n19159));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n19158));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n19157));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n19156));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n19155));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n19154));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n19153));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n19152));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n19151));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n19150));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n19149));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n19148));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n19147));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n19236));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n19235));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n19234));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n19233));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n19146));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n19232));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n19231));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n19230));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n19145));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n19144));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n19143));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n19142));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n19141));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n19140));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n19139));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n19138));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n19241));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n19137));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n19136));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut (.I0(n37401), .I1(n18140), .I2(n17542), .I3(n6), 
            .O(n38588));   // verilog/coms.v(69[16:27])
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n19135));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n19189));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n19229));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n19188));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n19134));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n19133));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n19132));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n19187));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n19131));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n19130));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n19228));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i14132_3_lut_4_lut (.I0(n8), .I1(n37361), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n19164));
    defparam i14132_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n19227));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n19226));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n19225));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n19186));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n19129));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n19185));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n19128));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n19184));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i14133_3_lut_4_lut (.I0(n8), .I1(n37361), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n19165));
    defparam i14133_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n19183));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n19182));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n19181));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n19127));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_871 (.I0(\data_in_frame[18] [2]), .I1(n8_adj_3906), 
            .I2(\data_in_frame[20] [3]), .I3(n37953), .O(n10));
    defparam i4_4_lut_adj_871.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n19180));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n19179));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n19178));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n19177));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n19176));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i14134_3_lut_4_lut (.I0(n8), .I1(n37361), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n19166));
    defparam i14134_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14135_3_lut_4_lut (.I0(n8), .I1(n37361), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n19167));
    defparam i14135_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14136_3_lut_4_lut (.I0(n8), .I1(n37361), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n19168));
    defparam i14136_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n19126));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_20 (.CI(n30319), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n30320));
    SB_LUT4 i14177_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37342), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n19209));
    defparam i14177_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut (.I0(n17266), .I1(n14748), .I2(n14721), .I3(n17199), 
            .O(n9));
    defparam i1_4_lut.LUT_INIT = 16'h50dc;
    SB_LUT4 i14178_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37342), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n19210));
    defparam i14178_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_out_frame[5] [2]), .I1(n37588), .I2(n37520), 
            .I3(\data_out_frame[7] [4]), .O(n17988));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14179_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37342), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n19211));
    defparam i14179_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14180_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37342), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n19212));
    defparam i14180_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_872 (.I0(\FRAME_MATCHER.state[3] ), .I1(n200), 
            .I2(n322), .I3(n326), .O(n6_adj_3908));   // verilog/coms.v(113[11:12])
    defparam i1_4_lut_adj_872.LUT_INIT = 16'haaa8;
    SB_LUT4 i14181_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37342), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n19213));
    defparam i14181_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_873 (.I0(n17170), .I1(n6_adj_3908), .I2(\FRAME_MATCHER.state_31__N_2492 [3]), 
            .I3(n17025), .O(n36609));   // verilog/coms.v(113[11:12])
    defparam i1_4_lut_adj_873.LUT_INIT = 16'hccdc;
    SB_LUT4 i1_3_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(n324), .I2(n301), 
            .I3(GND_net), .O(n36589));
    defparam i1_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 mux_666_i1_3_lut_4_lut (.I0(n31), .I1(Kp_23__N_1745), .I2(\FRAME_MATCHER.state[0] ), 
            .I3(tx_transmit_N_3215), .O(n3086[0]));   // verilog/coms.v(230[9] 232[65])
    defparam mux_666_i1_3_lut_4_lut.LUT_INIT = 16'hf404;
    SB_LUT4 i1_2_lut_adj_874 (.I0(n63_c), .I1(n63_adj_3909), .I2(GND_net), 
            .I3(GND_net), .O(n20661));   // verilog/coms.v(139[7:80])
    defparam i1_2_lut_adj_874.LUT_INIT = 16'h8888;
    SB_LUT4 i14182_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37342), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n19214));
    defparam i14182_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_357_Select_1_i5_4_lut (.I0(n63), .I1(n17268), .I2(n2857), 
            .I3(n93[1]), .O(n5_c));
    defparam select_357_Select_1_i5_4_lut.LUT_INIT = 16'h3331;
    SB_LUT4 i1_2_lut_3_lut (.I0(n31), .I1(Kp_23__N_1745), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n4658));   // verilog/coms.v(230[9] 232[65])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i2_4_lut (.I0(n93[1]), .I1(n5_c), .I2(n38098), .I3(n63), 
            .O(n6_adj_3911));
    defparam i2_4_lut.LUT_INIT = 16'hcecf;
    SB_LUT4 i14183_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37342), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n19215));
    defparam i14183_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut (.I0(n17200), .I1(n6_adj_3911), .I2(\FRAME_MATCHER.state_31__N_2460 [1]), 
            .I3(n17202), .O(n46228));
    defparam i3_4_lut.LUT_INIT = 16'hddfd;
    SB_LUT4 i14184_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37342), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n19216));
    defparam i14184_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n19125));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n40932), .I3(n40931), .O(tx_data[7]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n19124));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n19123));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n19122));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[8] [7]), .I3(\data_out_frame[11] [3]), .O(n37839));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n19121));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_adj_875 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[5] [0]), .I3(GND_net), .O(n17979));
    defparam i1_2_lut_3_lut_adj_875.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n19120));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n19119));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n19118));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n19117));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n19116));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n19115));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n19114));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n19224));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n19113));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 mux_1033_i3_3_lut (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n4658), .I3(GND_net), .O(n4661));
    defparam mux_1033_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n19112));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n19223));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n40929), .I3(n40928), .O(tx_data[6]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n19111));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n40926), .I3(n40925), .O(tx_data[5]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n19110));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut (.I0(byte_transmit_counter[4]), 
            .I1(byte_transmit_counter[3]), .I2(n40923), .I3(n40922), .O(tx_data[3]));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n19222));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i14225_3_lut_4_lut (.I0(n8_adj_3912), .I1(n37342), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n19257));
    defparam i14225_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14226_3_lut_4_lut (.I0(n8_adj_3912), .I1(n37342), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n19258));
    defparam i14226_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14227_3_lut_4_lut (.I0(n8_adj_3912), .I1(n37342), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n19259));
    defparam i14227_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14228_3_lut_4_lut (.I0(n8_adj_3912), .I1(n37342), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n19260));
    defparam i14228_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14229_3_lut_4_lut (.I0(n8_adj_3912), .I1(n37342), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n19261));
    defparam i14229_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1033_i1_3_lut (.I0(\data_in_frame[16] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n4658), .I3(GND_net), .O(n4659));
    defparam mux_1033_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14230_3_lut_4_lut (.I0(n8_adj_3912), .I1(n37342), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n19262));
    defparam i14230_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14231_3_lut_4_lut (.I0(n8_adj_3912), .I1(n37342), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n19263));
    defparam i14231_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14232_3_lut_4_lut (.I0(n8_adj_3912), .I1(n37342), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n19264));
    defparam i14232_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_876 (.I0(n37440), .I1(n37786), .I2(\data_out_frame[12] [2]), 
            .I3(GND_net), .O(n37735));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_3_lut_adj_876.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_877 (.I0(n33079), .I1(n33882), .I2(n17664), .I3(\data_out_frame[20] [5]), 
            .O(n38713));
    defparam i3_4_lut_adj_877.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_878 (.I0(n18200), .I1(\data_out_frame[20] [2]), 
            .I2(n37604), .I3(GND_net), .O(n37549));   // verilog/coms.v(71[16:42])
    defparam i1_3_lut_adj_878.LUT_INIT = 16'h9696;
    SB_CARRY add_44_16 (.CI(n30315), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n30316));
    SB_LUT4 add_44_15_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n30314), .O(n2_adj_3913)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_15 (.CI(n30314), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n30315));
    SB_LUT4 i3_4_lut_adj_879 (.I0(\data_in_frame[19] [7]), .I1(n37738), 
            .I2(n37723), .I3(\data_in_frame[20] [1]), .O(n38953));
    defparam i3_4_lut_adj_879.LUT_INIT = 16'h6996;
    SB_LUT4 add_44_14_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n30313), .O(n2_adj_3914)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_14_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n19109));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_880 (.I0(n33902), .I1(n33882), .I2(GND_net), 
            .I3(GND_net), .O(n32998));
    defparam i1_2_lut_adj_880.LUT_INIT = 16'h6666;
    SB_CARRY add_44_14 (.CI(n30313), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n30314));
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n19108));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n19107));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n19106));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n19105));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n19104));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_881 (.I0(n17671), .I1(n32998), .I2(n18200), .I3(n6_adj_3915), 
            .O(n37801));
    defparam i4_4_lut_adj_881.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_882 (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[19] [6]), 
            .I2(n37640), .I3(n33047), .O(n37666));
    defparam i3_4_lut_adj_882.LUT_INIT = 16'h6996;
    SB_LUT4 i14424_4_lut_4_lut (.I0(n18435), .I1(n6119), .I2(ID0), .I3(\data_out_frame[0] [0]), 
            .O(n19456));
    defparam i14424_4_lut_4_lut.LUT_INIT = 16'h7520;
    SB_LUT4 i5_4_lut (.I0(\data_out_frame[20] [4]), .I1(n37467), .I2(\data_out_frame[20] [3]), 
            .I3(\data_out_frame[20] [5]), .O(n12));   // verilog/coms.v(71[16:42])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n19103));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n19102));   // verilog/coms.v(126[12] 289[6])
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3228  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut (.I0(\data_out_frame[20] [1]), .I1(n12), .I2(n33016), 
            .I3(\data_out_frame[20] [2]), .O(n37482));   // verilog/coms.v(71[16:42])
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_883 (.I0(n37869), .I1(\data_out_frame[20] [0]), 
            .I2(n33902), .I3(n37872), .O(n10_adj_3916));
    defparam i4_4_lut_adj_883.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(n37482), .I1(n10_adj_3916), .I2(\data_out_frame[19] [5]), 
            .I3(GND_net), .O(n38644));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i13818_4_lut_4_lut (.I0(n18435), .I1(n6119), .I2(ID2), .I3(\data_out_frame[0] [2]), 
            .O(n18850));
    defparam i13818_4_lut_4_lut.LUT_INIT = 16'hfda8;
    SB_LUT4 add_44_13_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n30312), .O(n2_adj_3917)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15524_3_lut_4_lut (.I0(\data_in_frame[2] [0]), .I1(n37514), 
            .I2(\data_in_frame[1] [0]), .I3(n37386), .O(n12_adj_3918));   // verilog/coms.v(83[17:70])
    defparam i15524_3_lut_4_lut.LUT_INIT = 16'h0990;
    SB_LUT4 i1_4_lut_4_lut (.I0(n18381), .I1(n10308), .I2(n2236[0]), .I3(byte_transmit_counter[0]), 
            .O(n19453));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hd580;
    SB_LUT4 i4_4_lut_adj_884 (.I0(\data_out_frame[19] [3]), .I1(\data_out_frame[19] [4]), 
            .I2(n33049), .I3(n6_adj_3919), .O(n38639));
    defparam i4_4_lut_adj_884.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_885 (.I0(n33941), .I1(n37720), .I2(GND_net), 
            .I3(GND_net), .O(n37721));
    defparam i1_2_lut_adj_885.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_886 (.I0(n37735), .I1(\data_out_frame[18] [6]), 
            .I2(\data_out_frame[14] [5]), .I3(n37744), .O(n10_adj_3920));
    defparam i4_4_lut_adj_886.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_887 (.I0(n37673), .I1(n4_c), .I2(n10_adj_3920), 
            .I3(\data_out_frame[18] [7]), .O(n39012));
    defparam i2_4_lut_adj_887.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut (.I0(n33902), .I1(n37479), .I2(\data_out_frame[19] [0]), 
            .I3(GND_net), .O(n33016));
    defparam i2_3_lut.LUT_INIT = 16'h6969;
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n19101));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n19221));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n19273));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n19272));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n19271));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n19270));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n19100));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n19099));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_4_lut_adj_888 (.I0(n37508), .I1(\data_out_frame[12] [5]), 
            .I2(n37701), .I3(n32950), .O(n10_adj_3921));
    defparam i2_4_lut_adj_888.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_889 (.I0(n37814), .I1(\data_out_frame[14] [7]), 
            .I2(n32979), .I3(n1595), .O(n14));
    defparam i6_4_lut_adj_889.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(n39220), .I1(n14), .I2(n10_adj_3921), .I3(n1185), 
            .O(n33822));
    defparam i7_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i5_4_lut_adj_890 (.I0(\data_out_frame[15] [0]), .I1(n17325), 
            .I2(n37530), .I3(n17782), .O(n12_adj_3922));   // verilog/coms.v(74[16:43])
    defparam i5_4_lut_adj_890.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_891 (.I0(n17626), .I1(n12_adj_3922), .I2(\data_out_frame[17] [2]), 
            .I3(\data_out_frame[12] [6]), .O(n33049));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_891.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_892 (.I0(n37890), .I1(n37647), .I2(\data_out_frame[16] [7]), 
            .I3(n37962), .O(n10_adj_3923));
    defparam i4_4_lut_adj_892.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_4_lut_adj_893 (.I0(n18381), .I1(n10308), .I2(n2236[6]), 
            .I3(byte_transmit_counter[6]), .O(n19324));
    defparam i1_4_lut_4_lut_adj_893.LUT_INIT = 16'hd580;
    SB_LUT4 i6_4_lut_adj_894 (.I0(n33067), .I1(n37962), .I2(n37744), .I3(\data_out_frame[17] [0]), 
            .O(n16_c));
    defparam i6_4_lut_adj_894.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_895 (.I0(n33822), .I1(n37380), .I2(n37911), .I3(n1642), 
            .O(n17));
    defparam i7_4_lut_adj_895.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(n38802), .I2(n16_c), .I3(n37735), 
            .O(n32717));
    defparam i9_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_896 (.I0(\data_out_frame[19] [3]), .I1(\data_out_frame[19] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n37720));
    defparam i1_2_lut_adj_896.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_897 (.I0(\data_out_frame[19] [5]), .I1(\data_out_frame[19] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n37717));
    defparam i1_2_lut_adj_897.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_898 (.I0(n17969), .I1(n37707), .I2(GND_net), 
            .I3(GND_net), .O(n17746));
    defparam i1_2_lut_adj_898.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut (.I0(n324), .I1(n17183), .I2(n9), .I3(\FRAME_MATCHER.state [4]), 
            .O(n36679));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hba00;
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n19098));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n19097));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_899 (.I0(n33880), .I1(n17778), .I2(n33893), .I3(\data_in_frame[18] [2]), 
            .O(n10_adj_3924));
    defparam i4_4_lut_adj_899.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_900 (.I0(\data_out_frame[13] [4]), .I1(n32979), 
            .I2(n37407), .I3(n6_adj_3925), .O(n16772));
    defparam i4_4_lut_adj_900.LUT_INIT = 16'h6996;
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n19352));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_901 (.I0(\data_out_frame[18] [1]), .I1(\data_out_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3926));
    defparam i1_2_lut_adj_901.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_902 (.I0(n16772), .I1(n17969), .I2(n37613), .I3(n6_adj_3926), 
            .O(n37604));
    defparam i4_4_lut_adj_902.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_903 (.I0(n16772), .I1(n37807), .I2(\data_out_frame[18] [2]), 
            .I3(GND_net), .O(n17671));
    defparam i2_3_lut_adj_903.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_904 (.I0(n17671), .I1(n37604), .I2(GND_net), 
            .I3(GND_net), .O(n32719));
    defparam i1_2_lut_adj_904.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n19238));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_905 (.I0(\data_out_frame[17] [6]), .I1(n37508), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3927));
    defparam i1_2_lut_adj_905.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_906 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[13] [3]), .I3(n6_adj_3927), .O(n37707));
    defparam i4_4_lut_adj_906.LUT_INIT = 16'h6996;
    SB_CARRY add_44_13 (.CI(n30312), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n30313));
    SB_LUT4 i2_3_lut_adj_907 (.I0(n37539), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[15] [6]), .I3(GND_net), .O(n37613));
    defparam i2_3_lut_adj_907.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_908 (.I0(n17963), .I1(n37504), .I2(\data_out_frame[17] [5]), 
            .I3(n37578), .O(n33875));
    defparam i3_4_lut_adj_908.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n19237));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_12_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n30311), .O(n2_adj_3928)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_909 (.I0(n37613), .I1(n37707), .I2(\data_out_frame[18] [0]), 
            .I3(GND_net), .O(n18200));
    defparam i2_3_lut_adj_909.LUT_INIT = 16'h9696;
    SB_CARRY add_44_12 (.CI(n30311), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n30312));
    SB_LUT4 add_44_11_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n30310), .O(n2_adj_3929)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_910 (.I0(n33845), .I1(n37673), .I2(\data_out_frame[18] [5]), 
            .I3(GND_net), .O(n33902));
    defparam i2_3_lut_adj_910.LUT_INIT = 16'h9696;
    SB_LUT4 i36207_2_lut (.I0(\data_out_frame[0] [0]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n42985));
    defparam i36207_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i33786_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n40910));
    defparam i33786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i19_3_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\data_out_frame[21] [0]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n19096));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n19220));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_911 (.I0(n18200), .I1(n33875), .I2(GND_net), 
            .I3(GND_net), .O(n37863));
    defparam i1_2_lut_adj_911.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n19095));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_adj_912 (.I0(n37492), .I1(\data_out_frame[18] [3]), 
            .I2(n39208), .I3(GND_net), .O(n33882));
    defparam i2_3_lut_adj_912.LUT_INIT = 16'h6969;
    SB_LUT4 i33810_4_lut (.I0(n19), .I1(\data_out_frame[22] [0]), .I2(byte_transmit_counter[1]), 
            .I3(byte_transmit_counter[0]), .O(n40934));
    defparam i33810_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i33787_4_lut (.I0(n40910), .I1(n42985), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[1]), .O(n40911));
    defparam i33787_4_lut.LUT_INIT = 16'ha0ac;
    SB_LUT4 i3_4_lut_adj_913 (.I0(\data_out_frame[13] [4]), .I1(n37601), 
            .I2(n18143), .I3(n17916), .O(n17638));
    defparam i3_4_lut_adj_913.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_914 (.I0(n18147), .I1(n17638), .I2(\data_out_frame[13] [5]), 
            .I3(n17979), .O(n10_adj_3930));
    defparam i4_4_lut_adj_914.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_915 (.I0(n37422), .I1(n10_adj_3930), .I2(n17916), 
            .I3(GND_net), .O(n37539));
    defparam i5_3_lut_adj_915.LUT_INIT = 16'h9696;
    SB_LUT4 i33785_3_lut (.I0(\data_out_frame[4][0] ), .I1(\data_out_frame[5] [0]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n40909));
    defparam i33785_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n19094));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i37374_3_lut (.I0(n46031), .I1(n45881), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n44499));
    defparam i37374_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_916 (.I0(\data_out_frame[17] [1]), .I1(n39027), 
            .I2(n37539), .I3(GND_net), .O(n37911));
    defparam i1_3_lut_adj_916.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_917 (.I0(n33815), .I1(n37911), .I2(GND_net), 
            .I3(GND_net), .O(n37890));
    defparam i1_2_lut_adj_917.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_918 (.I0(\data_out_frame[4][2] ), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n37561));
    defparam i1_2_lut_adj_918.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_919 (.I0(n37561), .I1(\data_out_frame[10] [7]), 
            .I2(\data_out_frame[6] [3]), .I3(n37884), .O(n10_adj_3931));
    defparam i4_4_lut_adj_919.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_920 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n37413));
    defparam i1_2_lut_adj_920.LUT_INIT = 16'h6666;
    SB_LUT4 i33811_3_lut (.I0(n45941), .I1(n40934), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n40935));
    defparam i33811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_921 (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n37634));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_921.LUT_INIT = 16'h6666;
    SB_LUT4 i37603_3_lut (.I0(n40912), .I1(n44499), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n44728));   // verilog/coms.v(104[34:55])
    defparam i37603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut_adj_922 (.I0(n37486), .I1(\data_out_frame[8] [4]), 
            .I2(\data_out_frame[6] [1]), .I3(n37763), .O(n10_adj_3932));   // verilog/coms.v(71[16:42])
    defparam i4_4_lut_adj_922.LUT_INIT = 16'h6996;
    SB_LUT4 i37604_4_lut (.I0(n44728), .I1(n40935), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(tx_data[0]));   // verilog/coms.v(104[34:55])
    defparam i37604_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i5_3_lut_adj_923 (.I0(\data_out_frame[6] [3]), .I1(n10_adj_3932), 
            .I2(\data_out_frame[8] [3]), .I3(GND_net), .O(n17782));   // verilog/coms.v(71[16:42])
    defparam i5_3_lut_adj_923.LUT_INIT = 16'h9696;
    SB_LUT4 i14281_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37354), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n19313));
    defparam i14281_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i23_4_lut (.I0(\data_out_frame[5] [3]), .I1(n37552), .I2(\data_out_frame[5] [4]), 
            .I3(n18209), .O(n54));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14282_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37354), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n19314));
    defparam i14282_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14283_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37354), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n19315));
    defparam i14283_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n19093));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n19092));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i21_4_lut (.I0(n37473), .I1(\data_out_frame[10] [6]), .I2(n37395), 
            .I3(\data_out_frame[6] [5]), .O(n52));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14284_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37354), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n19316));
    defparam i14284_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i22_4_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[11] [2]), .I3(\data_out_frame[12] [0]), 
            .O(n53));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(\data_out_frame[9] [6]), .I1(n37884), .I2(\data_out_frame[12] [2]), 
            .I3(n37786), .O(n51));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut (.I0(n17782), .I1(\data_out_frame[12] [1]), .I2(\data_out_frame[12] [3]), 
            .I3(n37935), .O(n48));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut (.I0(n37804), .I1(\data_out_frame[11] [5]), .I2(n37419), 
            .I3(\data_out_frame[10] [4]), .O(n50));
    defparam i19_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[11] [6]), 
            .I2(n37652), .I3(n18079), .O(n49));
    defparam i18_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i29_4_lut (.I0(n51), .I1(n53), .I2(n52), .I3(n54), .O(n60));
    defparam i29_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut (.I0(n37501), .I1(n48), .I2(\data_out_frame[12] [4]), 
            .I3(n1559), .O(n55));
    defparam i24_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut (.I0(n55), .I1(n60), .I2(n49), .I3(n50), .O(n37701));
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_924 (.I0(n16906), .I1(n37701), .I2(\data_out_frame[13] [0]), 
            .I3(GND_net), .O(n39220));
    defparam i2_3_lut_adj_924.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_925 (.I0(\data_out_frame[14] [5]), .I1(n16906), 
            .I2(GND_net), .I3(GND_net), .O(n32972));
    defparam i1_2_lut_adj_925.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n19091));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n19090));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n19089));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n19088));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n19087));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n19086));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n19085));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_926 (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[14] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n37530));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_926.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_927 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n37704));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_927.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n19084));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i14285_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37354), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n19317));
    defparam i14285_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n19083));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_928 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n17963));
    defparam i1_2_lut_adj_928.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n19082));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_929 (.I0(\data_out_frame[13] [2]), .I1(\data_out_frame[13] [4]), 
            .I2(n37704), .I3(\data_out_frame[13] [3]), .O(n39565));   // verilog/coms.v(83[17:28])
    defparam i3_4_lut_adj_929.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n19081));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_11 (.CI(n30310), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n30311));
    SB_LUT4 i14286_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37354), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n19318));
    defparam i14286_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14287_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37354), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n19319));
    defparam i14287_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_930 (.I0(\data_out_frame[13] [1]), .I1(n39565), 
            .I2(n37575), .I3(n32972), .O(n18));
    defparam i7_4_lut_adj_930.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_931 (.I0(\data_out_frame[12] [5]), .I1(n18), .I2(n37404), 
            .I3(\data_out_frame[14] [1]), .O(n20));
    defparam i9_4_lut_adj_931.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut (.I0(n15), .I1(n20), .I2(n39220), .I3(\data_out_frame[14] [2]), 
            .O(n33815));
    defparam i10_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i14288_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37354), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n19320));
    defparam i14288_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n19080));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_932 (.I0(n33815), .I1(n37687), .I2(\data_out_frame[15] [2]), 
            .I3(\data_out_frame[15] [1]), .O(n38802));
    defparam i3_4_lut_adj_932.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_933 (.I0(\data_in_frame[6] [2]), .I1(n18119), .I2(GND_net), 
            .I3(GND_net), .O(n17404));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_933.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_934 (.I0(\data_in_frame[16] [1]), .I1(n37517), 
            .I2(\data_in_frame[20] [5]), .I3(n33035), .O(n38540));
    defparam i3_4_lut_adj_934.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_935 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n37804));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_935.LUT_INIT = 16'h6666;
    SB_LUT4 add_44_10_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n30309), .O(n2_adj_3934)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_10_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n19079));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_936 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n37486));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_936.LUT_INIT = 16'h6666;
    SB_LUT4 i803_2_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1559));   // verilog/coms.v(69[16:27])
    defparam i803_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n19078));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_4_lut_adj_937 (.I0(n17860), .I1(n1559), .I2(n17325), .I3(n17422), 
            .O(n12_adj_3935));   // verilog/coms.v(74[16:43])
    defparam i5_4_lut_adj_937.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_938 (.I0(\data_out_frame[13] [0]), .I1(n12_adj_3935), 
            .I2(n37504), .I3(\data_out_frame[10] [6]), .O(n1642));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_938.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_939 (.I0(n37486), .I1(n17365), .I2(\data_out_frame[8] [6]), 
            .I3(n37804), .O(n10_adj_3936));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_939.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n19077));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_940 (.I0(\data_out_frame[13] [1]), .I1(n1595), 
            .I2(GND_net), .I3(GND_net), .O(n37504));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_940.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_941 (.I0(\data_out_frame[15] [2]), .I1(n1642), 
            .I2(GND_net), .I3(GND_net), .O(n37647));
    defparam i1_2_lut_adj_941.LUT_INIT = 16'h6666;
    SB_LUT4 i14217_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37342), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n19249));
    defparam i14217_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_942 (.I0(\data_out_frame[10] [2]), .I1(n37572), 
            .I2(n18079), .I3(n17817), .O(n17626));
    defparam i3_4_lut_adj_942.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_943 (.I0(n37655), .I1(n37875), .I2(\data_in_frame[1] [6]), 
            .I3(GND_net), .O(n17844));   // verilog/coms.v(68[16:27])
    defparam i2_3_lut_adj_943.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_944 (.I0(\data_out_frame[16] [6]), .I1(n17626), 
            .I2(GND_net), .I3(GND_net), .O(n37992));
    defparam i1_2_lut_adj_944.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_945 (.I0(n37647), .I1(n37504), .I2(\data_out_frame[15] [3]), 
            .I3(n6_adj_3937), .O(n33047));
    defparam i4_4_lut_adj_945.LUT_INIT = 16'h6996;
    SB_LUT4 i8_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n25));
    defparam i8_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_946 (.I0(n37643), .I1(n38695), .I2(n37866), .I3(\data_in_frame[21] [5]), 
            .O(n19_adj_3938));
    defparam i3_4_lut_adj_946.LUT_INIT = 16'hb77b;
    SB_CARRY add_44_10 (.CI(n30309), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n30310));
    SB_LUT4 i13_4_lut (.I0(n25), .I1(\data_out_frame[15] [0]), .I2(n38802), 
            .I3(n37422), .O(n30));
    defparam i13_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i14218_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37342), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n19250));
    defparam i14218_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n19076));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n19075));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n19074));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n19073));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i11_4_lut (.I0(\data_out_frame[9] [0]), .I1(n32972), .I2(n17764), 
            .I3(n37923), .O(n28));
    defparam i11_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n19072));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n19071));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n19070));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n19069));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n19068));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n19067));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n19066));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n19065));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n19269));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n19064));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n19268));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n19063));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12_4_lut (.I0(n37792), .I1(n37413), .I2(n37572), .I3(\data_out_frame[12] [3]), 
            .O(n29));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_947 (.I0(n37839), .I1(n37941), .I2(\data_out_frame[13] [5]), 
            .I3(n37634), .O(n27));
    defparam i10_4_lut_adj_947.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n19062));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i16_4_lut (.I0(n27), .I1(n29), .I2(n28), .I3(n30), .O(n39027));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n19061));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n19060));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_4_lut_adj_948 (.I0(\data_out_frame[11] [0]), .I1(n37766), 
            .I2(\data_out_frame[8] [5]), .I3(\data_out_frame[11] [1]), .O(n12_adj_3939));
    defparam i5_4_lut_adj_948.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_949 (.I0(\data_out_frame[8] [7]), .I1(n12_adj_3939), 
            .I2(n37923), .I3(\data_out_frame[10] [6]), .O(n16787));
    defparam i6_4_lut_adj_949.LUT_INIT = 16'h6996;
    SB_LUT4 i14219_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37342), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n19251));
    defparam i14219_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_950 (.I0(\data_out_frame[13] [2]), .I1(n16787), 
            .I2(GND_net), .I3(GND_net), .O(n37416));
    defparam i1_2_lut_adj_950.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_951 (.I0(\data_out_frame[9] [3]), .I1(n16915), 
            .I2(n17979), .I3(\data_out_frame[7] [1]), .O(n37575));
    defparam i3_4_lut_adj_951.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_952 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[8] [4]), .I3(GND_net), .O(n37766));
    defparam i2_3_lut_adj_952.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n19059));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n19058));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n19057));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n19056));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n19055));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n19054));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n19053));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n19052));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n19051));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n19050));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n19049));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n19048));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n19047));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n19046));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n19045));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n19044));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n19043));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i14220_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37342), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n19252));
    defparam i14220_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14221_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37342), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n19253));
    defparam i14221_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_953 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n18147));
    defparam i1_2_lut_adj_953.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_954 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[11] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n37935));
    defparam i1_2_lut_adj_954.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_955 (.I0(n37935), .I1(\data_out_frame[8] [7]), 
            .I2(\data_out_frame[6] [7]), .I3(n6_adj_3940), .O(n37404));
    defparam i4_4_lut_adj_955.LUT_INIT = 16'h6996;
    SB_LUT4 add_44_9_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n30308), .O(n2_adj_3941)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_956 (.I0(\data_out_frame[16] [1]), .I1(n37757), 
            .I2(\data_out_frame[13] [5]), .I3(n17988), .O(n10_adj_3942));
    defparam i4_4_lut_adj_956.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_957 (.I0(n37404), .I1(n10_adj_3942), .I2(\data_out_frame[15] [7]), 
            .I3(GND_net), .O(n37492));
    defparam i5_3_lut_adj_957.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_958 (.I0(\data_out_frame[4][0] ), .I1(\data_out_frame[6] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n17817));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_958.LUT_INIT = 16'h6666;
    SB_LUT4 i14222_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37342), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n19254));
    defparam i14222_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_959 (.I0(\data_out_frame[6] [2]), .I1(n1119), .I2(\data_out_frame[6] [0]), 
            .I3(n6_adj_3943), .O(n17325));   // verilog/coms.v(71[16:42])
    defparam i4_4_lut_adj_959.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_960 (.I0(\data_out_frame[10] [3]), .I1(n17325), 
            .I2(n17817), .I3(n6_adj_3944), .O(n16906));
    defparam i4_4_lut_adj_960.LUT_INIT = 16'h6996;
    SB_LUT4 i14223_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37342), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n19255));
    defparam i14223_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_961 (.I0(\data_out_frame[12] [5]), .I1(n16906), 
            .I2(\data_out_frame[14] [6]), .I3(GND_net), .O(n37380));
    defparam i2_3_lut_adj_961.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n19267));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_962 (.I0(\data_out_frame[17] [0]), .I1(\data_out_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_3945));
    defparam i1_2_lut_adj_962.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_adj_963 (.I0(n37380), .I1(n4_adj_3945), .I2(n37741), 
            .I3(n38435), .O(n37658));
    defparam i2_4_lut_adj_963.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_964 (.I0(\data_out_frame[16] [5]), .I1(n33067), 
            .I2(\data_out_frame[14] [5]), .I3(GND_net), .O(n37741));
    defparam i2_3_lut_adj_964.LUT_INIT = 16'h9696;
    SB_LUT4 i14224_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37342), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n19256));
    defparam i14224_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_965 (.I0(n37578), .I1(n17638), .I2(\data_out_frame[15] [5]), 
            .I3(GND_net), .O(n17969));
    defparam i2_3_lut_adj_965.LUT_INIT = 16'h9696;
    SB_CARRY add_44_9 (.CI(n30308), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n30309));
    SB_LUT4 i22_4_lut_adj_966 (.I0(\data_out_frame[17] [6]), .I1(n39208), 
            .I2(n17969), .I3(\data_out_frame[17] [5]), .O(n52_adj_3946));
    defparam i22_4_lut_adj_966.LUT_INIT = 16'h9669;
    SB_LUT4 i14273_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37354), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n19305));
    defparam i14273_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i20_4_lut_adj_967 (.I0(n37965), .I1(n37741), .I2(n37807), 
            .I3(n37658), .O(n50_adj_3948));
    defparam i20_4_lut_adj_967.LUT_INIT = 16'h6996;
    SB_LUT4 i14274_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37354), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n19306));
    defparam i14274_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14275_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37354), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n19307));
    defparam i14275_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21_4_lut_adj_968 (.I0(n37416), .I1(n17330), .I2(\data_out_frame[11] [3]), 
            .I3(\data_out_frame[15] [4]), .O(n51_adj_3949));
    defparam i21_4_lut_adj_968.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_969 (.I0(n39027), .I1(n33047), .I2(\data_out_frame[16] [3]), 
            .I3(n37992), .O(n49_adj_3950));
    defparam i19_4_lut_adj_969.LUT_INIT = 16'h9669;
    SB_LUT4 i16_4_lut_adj_970 (.I0(n37977), .I1(n37578), .I2(\data_out_frame[9] [1]), 
            .I3(\data_out_frame[15] [6]), .O(n46));
    defparam i16_4_lut_adj_970.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n19042));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_8_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n30307), .O(n2_adj_3951)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_8_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n19041));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n19040));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n19039));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n19038));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n19266));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n19037));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_8 (.CI(n30307), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n30308));
    SB_LUT4 i18_4_lut_adj_971 (.I0(n37890), .I1(\data_out_frame[16] [4]), 
            .I2(n37704), .I3(\data_out_frame[13] [5]), .O(n48_adj_3952));
    defparam i18_4_lut_adj_971.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_972 (.I0(n37766), .I1(\data_out_frame[14] [1]), 
            .I2(n32716), .I3(\data_out_frame[17] [7]), .O(n47));
    defparam i17_4_lut_adj_972.LUT_INIT = 16'h6996;
    SB_LUT4 i28_4_lut (.I0(n49_adj_3950), .I1(n51_adj_3949), .I2(n50_adj_3948), 
            .I3(n52_adj_3946), .O(n58));
    defparam i28_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i23_3_lut (.I0(\data_out_frame[17] [3]), .I1(n46), .I2(n37665), 
            .I3(GND_net), .O(n53_adj_3953));
    defparam i23_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 add_44_7_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n30306), .O(n2_adj_3954)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i29_4_lut_adj_973 (.I0(n53_adj_3953), .I1(n58), .I2(n47), 
            .I3(n48_adj_3952), .O(n39387));
    defparam i29_4_lut_adj_973.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_974 (.I0(\data_out_frame[18] [4]), .I1(\data_out_frame[18] [7]), 
            .I2(n37798), .I3(n32719), .O(n16_adj_3955));
    defparam i6_4_lut_adj_974.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_975 (.I0(n39387), .I1(n33882), .I2(n37863), .I3(n33902), 
            .O(n17_adj_3956));
    defparam i7_4_lut_adj_975.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_976 (.I0(n17_adj_3956), .I1(n16817), .I2(n16_adj_3955), 
            .I3(n17746), .O(n38620));
    defparam i9_4_lut_adj_976.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_977 (.I0(n37717), .I1(\data_out_frame[19] [7]), 
            .I2(\data_out_frame[19] [1]), .I3(n37720), .O(n10_adj_3957));
    defparam i4_4_lut_adj_977.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_978 (.I0(n33875), .I1(\data_out_frame[19] [6]), 
            .I2(n10_adj_3957), .I3(n38620), .O(n37479));
    defparam i1_4_lut_adj_978.LUT_INIT = 16'h9669;
    SB_LUT4 i14276_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37354), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n19308));
    defparam i14276_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14277_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37354), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n19309));
    defparam i14277_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14278_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37354), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n19310));
    defparam i14278_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_979 (.I0(\data_out_frame[18] [7]), .I1(n37658), 
            .I2(GND_net), .I3(GND_net), .O(n33008));
    defparam i1_2_lut_adj_979.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n19036));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n19035));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n19034));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n19033));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n19032));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n19265));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_7 (.CI(n30306), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n30307));
    SB_LUT4 i4_4_lut_adj_980 (.I0(n37665), .I1(n33941), .I2(n33008), .I3(n37479), 
            .O(n10_adj_3958));
    defparam i4_4_lut_adj_980.LUT_INIT = 16'h6996;
    SB_LUT4 add_44_6_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n30305), .O(n2_adj_3959)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_6_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n19031));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_3_lut_adj_981 (.I0(n33016), .I1(n10_adj_3958), .I2(\data_out_frame[20] [7]), 
            .I3(GND_net), .O(n38514));
    defparam i5_3_lut_adj_981.LUT_INIT = 16'h6969;
    SB_LUT4 i14279_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37354), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n19311));
    defparam i14279_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_6 (.CI(n30305), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n30306));
    SB_LUT4 add_44_5_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n30304), .O(n2_adj_3960)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_5_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n19030));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n19029));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n19028));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n19027));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n19219));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i24201_3_lut (.I0(\data_out_frame[4] [1]), .I1(ID1), .I2(n14536), 
            .I3(GND_net), .O(n19016));
    defparam i24201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14280_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37354), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n19312));
    defparam i14280_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_982 (.I0(\data_in_frame[21] [7]), .I1(n37830), 
            .I2(n37555), .I3(n17833), .O(n39798));   // verilog/coms.v(73[16:43])
    defparam i3_4_lut_adj_982.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_983 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n17418));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_983.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n19218));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 mux_1033_i2_3_lut (.I0(\data_in_frame[16] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n4658), .I3(GND_net), .O(n4660));
    defparam mux_1033_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_44_5 (.CI(n30304), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n30305));
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n19026));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_984 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n37473));
    defparam i1_2_lut_adj_984.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_985 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n37786));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_985.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n19025));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n19024));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n19023));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n19022));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i3_4_lut_adj_986 (.I0(\data_out_frame[10] [1]), .I1(n17725), 
            .I2(\data_out_frame[5] [4]), .I3(n17330), .O(n37440));   // verilog/coms.v(72[16:27])
    defparam i3_4_lut_adj_986.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_987 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[10] [1]), 
            .I2(\data_out_frame[10] [2]), .I3(n17764), .O(n37652));
    defparam i3_4_lut_adj_987.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_988 (.I0(\data_out_frame[10] [1]), .I1(n17742), 
            .I2(GND_net), .I3(GND_net), .O(n37941));
    defparam i1_2_lut_adj_988.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_989 (.I0(\data_out_frame[12] [3]), .I1(n37652), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_3961));
    defparam i1_2_lut_adj_989.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_990 (.I0(\data_out_frame[6] [0]), .I1(n18031), 
            .I2(n17742), .I3(n6_adj_3961), .O(n33067));
    defparam i4_4_lut_adj_990.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_991 (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[16] [4]), 
            .I2(\data_out_frame[14] [3]), .I3(GND_net), .O(n14_adj_3962));
    defparam i5_3_lut_adj_991.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_992 (.I0(n37810), .I1(n33891), .I2(n37941), .I3(n37944), 
            .O(n15_adj_3963));
    defparam i6_4_lut_adj_992.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut (.I0(n15_adj_3963), .I1(n37827), .I2(n14_adj_3962), 
            .I3(n37496), .O(n37673));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_993 (.I0(n33891), .I1(n33067), .I2(n37588), .I3(n39794), 
            .O(n16_adj_3964));
    defparam i6_4_lut_adj_993.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_994 (.I0(n17_adj_3965), .I1(\data_out_frame[12] [1]), 
            .I2(n16_adj_3964), .I3(n18073), .O(n38435));
    defparam i9_4_lut_adj_994.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1033_i15_3_lut (.I0(\data_in_frame[15] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n4658), .I3(GND_net), .O(n4673));
    defparam mux_1033_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n19021));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk32MHz), 
           .D(n19020));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 mux_1033_i14_3_lut (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n4658), .I3(GND_net), .O(n4672));
    defparam mux_1033_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1033_i13_3_lut (.I0(\data_in_frame[15] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n4658), .I3(GND_net), .O(n4671));
    defparam mux_1033_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1033_i12_3_lut (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n4658), .I3(GND_net), .O(n4670));
    defparam mux_1033_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1033_i11_3_lut (.I0(\data_in_frame[15] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n4658), .I3(GND_net), .O(n4669));
    defparam mux_1033_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1033_i10_3_lut (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n4658), .I3(GND_net), .O(n4668));
    defparam mux_1033_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_2_lut (.I0(Kp_23__N_893), .I1(\data_in_frame[4] [6]), .I2(GND_net), 
            .I3(GND_net), .O(n11));   // verilog/coms.v(69[16:27])
    defparam i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_995 (.I0(\data_in_frame[3] [2]), .I1(\data_in_frame[3] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n37817));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_995.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_996 (.I0(\data_in_frame[5] [3]), .I1(n37899), .I2(n37817), 
            .I3(n15612), .O(n17687));   // verilog/coms.v(83[17:28])
    defparam i3_4_lut_adj_996.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n19019));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_997 (.I0(\data_out_frame[5] [1]), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n37588));
    defparam i1_2_lut_adj_997.LUT_INIT = 16'h6666;
    SB_LUT4 add_44_4_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n30303), .O(n2_adj_3966)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_2_lut_adj_998 (.I0(n17979), .I1(n37496), .I2(GND_net), 
            .I3(GND_net), .O(n17648));
    defparam i1_2_lut_adj_998.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_999 (.I0(n17648), .I1(\data_out_frame[14] [2]), 
            .I2(n17988), .I3(n6_adj_3967), .O(n37944));   // verilog/coms.v(83[17:28])
    defparam i4_4_lut_adj_999.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1000 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n37601));
    defparam i1_2_lut_adj_1000.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n19018));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1001 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[13] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n37757));
    defparam i1_2_lut_adj_1001.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1002 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [0]), .I3(GND_net), .O(n37591));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_adj_1002.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1003 (.I0(\data_out_frame[6] [5]), .I1(n37965), 
            .I2(n1287), .I3(\data_out_frame[8] [4]), .O(n37920));
    defparam i3_4_lut_adj_1003.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1004 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[8] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17860));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1004.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i35 (.Q(\data_out_frame[4][2] ), .C(clk32MHz), 
           .D(n19017));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i366_2_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1119));   // verilog/coms.v(83[17:28])
    defparam i366_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(clk32MHz), 
           .D(n19016));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i6_4_lut_adj_1005 (.I0(n1185), .I1(\data_out_frame[7] [3]), 
            .I2(\data_out_frame[7] [1]), .I3(\data_out_frame[7] [2]), .O(n15_adj_3968));   // verilog/coms.v(83[17:63])
    defparam i6_4_lut_adj_1005.LUT_INIT = 16'h6996;
    SB_CARRY add_44_4 (.CI(n30303), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n30304));
    SB_LUT4 i8_4_lut_adj_1006 (.I0(n15_adj_3968), .I1(n18219), .I2(n14_adj_3969), 
            .I3(\data_out_frame[7] [7]), .O(n37395));   // verilog/coms.v(83[17:63])
    defparam i8_4_lut_adj_1006.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1007 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[6] [1]), 
            .I2(n37395), .I3(n17422), .O(n12_adj_3970));
    defparam i5_4_lut_adj_1007.LUT_INIT = 16'h6996;
    SB_LUT4 add_44_3_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n30302), .O(n2_adj_3971)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_3 (.CI(n30302), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n30303));
    SB_LUT4 add_44_2_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [0]), .I2(n164), 
            .I3(GND_net), .O(n2_adj_3902)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i6_4_lut_adj_1008 (.I0(n17764), .I1(n12_adj_3970), .I2(\data_out_frame[6] [0]), 
            .I3(\data_out_frame[6] [3]), .O(n18292));
    defparam i6_4_lut_adj_1008.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1009 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n37419));
    defparam i1_2_lut_adj_1009.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i33 (.Q(\data_out_frame[4][0] ), .C(clk32MHz), 
           .D(n19014));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i5 (.Q(\data_out_frame[0][4] ), .C(clk32MHz), 
           .D(n19013));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_out_frame_0___i4 (.Q(\data_out_frame[0][3] ), .C(clk32MHz), 
           .D(n19012));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n19011));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n19010));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n19009));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n164), 
            .CO(n30302));
    SB_LUT4 add_624_9_lut (.I0(n10308), .I1(byte_transmit_counter[7]), .I2(GND_net), 
            .I3(n30339), .O(n42885)) /* synthesis syn_instantiated=1 */ ;
    defparam add_624_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_624_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n30338), .O(n2236[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_624_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i531_2_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1287));   // verilog/coms.v(69[16:27])
    defparam i531_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n19008));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n19007));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n19006));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n19005));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1010 (.I0(\data_out_frame[8] [0]), .I1(n17725), 
            .I2(GND_net), .I3(GND_net), .O(n32986));
    defparam i1_2_lut_adj_1010.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1011 (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[8] [2]), 
            .I2(\data_out_frame[5] [6]), .I3(GND_net), .O(n17821));
    defparam i2_3_lut_adj_1011.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1012 (.I0(\data_out_frame[9] [4]), .I1(\data_out_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n37552));
    defparam i1_2_lut_adj_1012.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1013 (.I0(\data_in_frame[3] [2]), .I1(n37750), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[5] [4]), .O(n37914));   // verilog/coms.v(94[12:25])
    defparam i3_4_lut_adj_1013.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1014 (.I0(n18082), .I1(n17821), .I2(n32986), 
            .I3(n37677), .O(n10_adj_3972));
    defparam i4_4_lut_adj_1014.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1015 (.I0(n17365), .I1(n10_adj_3972), .I2(n18292), 
            .I3(GND_net), .O(n33891));
    defparam i5_3_lut_adj_1015.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n19004));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1016 (.I0(n37501), .I1(n37827), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_3973));
    defparam i1_2_lut_adj_1016.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n19003));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n19002));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i4_4_lut_adj_1017 (.I0(\data_out_frame[11] [7]), .I1(n33891), 
            .I2(n37552), .I3(n6_adj_3973), .O(n39794));
    defparam i4_4_lut_adj_1017.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1018 (.I0(\data_out_frame[12] [0]), .I1(n39794), 
            .I2(GND_net), .I3(GND_net), .O(n37810));
    defparam i1_2_lut_adj_1018.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1019 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n18219));
    defparam i1_2_lut_adj_1019.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n19001));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_624_8 (.CI(n30338), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n30339));
    SB_LUT4 add_624_7_lut (.I0(n10308), .I1(byte_transmit_counter[5]), .I2(GND_net), 
            .I3(n30337), .O(n42882)) /* synthesis syn_instantiated=1 */ ;
    defparam add_624_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_1020 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[7] [1]), 
            .I2(\data_out_frame[9] [3]), .I3(GND_net), .O(n37422));
    defparam i2_3_lut_adj_1020.LUT_INIT = 16'h9696;
    SB_LUT4 i395_2_lut (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1185));   // verilog/coms.v(69[16:27])
    defparam i395_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1021 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[6] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n16915));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_1021.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1022 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[11] [5]), 
            .I2(n37842), .I3(\data_out_frame[16] [2]), .O(n18_adj_3974));
    defparam i7_4_lut_adj_1022.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n19000));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n18999));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i5_2_lut (.I0(n37407), .I1(\data_out_frame[14] [0]), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_3975));
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n18998));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i9_4_lut_adj_1023 (.I0(\data_out_frame[9] [4]), .I1(n18_adj_3974), 
            .I2(n37520), .I3(n37977), .O(n20_adj_3976));
    defparam i9_4_lut_adj_1023.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1024 (.I0(n37920), .I1(n20_adj_3976), .I2(n16_adj_3975), 
            .I3(n37591), .O(n39208));
    defparam i10_4_lut_adj_1024.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1025 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[1] [1]), .I3(GND_net), .O(n6_adj_3977));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_3_lut_adj_1025.LUT_INIT = 16'h9696;
    SB_CARRY add_624_7 (.CI(n30337), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n30338));
    SB_LUT4 i3_4_lut_adj_1026 (.I0(n39794), .I1(n37920), .I2(n37757), 
            .I3(n37601), .O(n38809));
    defparam i3_4_lut_adj_1026.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1027 (.I0(n37944), .I1(n18082), .I2(\data_out_frame[9] [7]), 
            .I3(\data_out_frame[5] [6]), .O(n14_adj_3978));
    defparam i6_4_lut_adj_1027.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1028 (.I0(\data_out_frame[16] [3]), .I1(n14_adj_3978), 
            .I2(n10_adj_3979), .I3(n38809), .O(n33845));
    defparam i7_4_lut_adj_1028.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1029 (.I0(n33845), .I1(n39208), .I2(GND_net), 
            .I3(GND_net), .O(n16817));
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'h9999;
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n18997));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n18996));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n18995));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n18994));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n18993));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n18992));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_4_lut_adj_1030 (.I0(\data_out_frame[18] [6]), .I1(n38435), 
            .I2(n37673), .I3(\data_out_frame[16] [5]), .O(n37798));
    defparam i1_4_lut_adj_1030.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1031 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n37467));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_1031.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1032 (.I0(n6119), .I1(n6121), .I2(GND_net), .I3(GND_net), 
            .O(n18436));   // verilog/coms.v(110[11:16])
    defparam i1_2_lut_adj_1032.LUT_INIT = 16'h2222;
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n18991));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n18990));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_624_6_lut (.I0(n10308), .I1(byte_transmit_counter[4]), .I2(GND_net), 
            .I3(n30336), .O(n42884)) /* synthesis syn_instantiated=1 */ ;
    defparam add_624_6_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n18989));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n18988));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n18987));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n18986));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n18985));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n18984));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n18983));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n18982));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n18981));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n18980));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n18979));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n18978));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n18977));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n18976));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n18975));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n18974));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n18973));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n18972));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n18971));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n18970));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n18969));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n18968));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n18967));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i23 (.Q(gearBoxRatio[23]), .C(clk32MHz), .D(n18966));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i22 (.Q(gearBoxRatio[22]), .C(clk32MHz), .D(n18965));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i21 (.Q(gearBoxRatio[21]), .C(clk32MHz), .D(n18964));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i20 (.Q(gearBoxRatio[20]), .C(clk32MHz), .D(n18963));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i19 (.Q(gearBoxRatio[19]), .C(clk32MHz), .D(n18962));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i18 (.Q(gearBoxRatio[18]), .C(clk32MHz), .D(n18961));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i17 (.Q(gearBoxRatio[17]), .C(clk32MHz), .D(n18960));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i16 (.Q(gearBoxRatio[16]), .C(clk32MHz), .D(n18959));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i15 (.Q(gearBoxRatio[15]), .C(clk32MHz), .D(n18958));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i14 (.Q(gearBoxRatio[14]), .C(clk32MHz), .D(n18957));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i13 (.Q(gearBoxRatio[13]), .C(clk32MHz), .D(n18956));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i12 (.Q(gearBoxRatio[12]), .C(clk32MHz), .D(n18955));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i11 (.Q(gearBoxRatio[11]), .C(clk32MHz), .D(n18954));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i10 (.Q(gearBoxRatio[10]), .C(clk32MHz), .D(n18953));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i9 (.Q(gearBoxRatio[9]), .C(clk32MHz), .D(n18952));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i8 (.Q(gearBoxRatio[8]), .C(clk32MHz), .D(n18951));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i7 (.Q(gearBoxRatio[7]), .C(clk32MHz), .D(n18950));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i6 (.Q(gearBoxRatio[6]), .C(clk32MHz), .D(n18949));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i5 (.Q(gearBoxRatio[5]), .C(clk32MHz), .D(n18948));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i4 (.Q(gearBoxRatio[4]), .C(clk32MHz), .D(n18947));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i3 (.Q(gearBoxRatio[3]), .C(clk32MHz), .D(n18946));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_624_6 (.CI(n30336), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n30337));
    SB_LUT4 i2_3_lut_adj_1033 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [2]), .I3(GND_net), .O(n4_adj_3980));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_1033.LUT_INIT = 16'h9696;
    SB_DFF gearBoxRatio_i0_i2 (.Q(gearBoxRatio[2]), .C(clk32MHz), .D(n18945));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i1 (.Q(gearBoxRatio[1]), .C(clk32MHz), .D(n18944));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i14167_3_lut_4_lut (.I0(n8_adj_3912), .I1(n37361), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n19199));
    defparam i14167_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n18937));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n18936));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13632_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[10] [0]), 
            .I3(IntegralLimit[0]), .O(n18664));   // verilog/coms.v(258[9] 260[65])
    defparam i13632_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14321_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[5] [6]), 
            .I3(PWMLimit[22]), .O(n19353));   // verilog/coms.v(258[9] 260[65])
    defparam i14321_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n18935));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n18934));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n18933));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13763_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[19] [0]), 
            .I3(gearBoxRatio[0]), .O(n18795));   // verilog/coms.v(258[9] 260[65])
    defparam i13763_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13764_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[2] [0]), 
            .I3(\Kp[0] ), .O(n18796));   // verilog/coms.v(258[9] 260[65])
    defparam i13764_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1034 (.I0(n37545), .I1(n37610), .I2(\data_in_frame[21] [2]), 
            .I3(GND_net), .O(n38719));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1034.LUT_INIT = 16'h9696;
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n18932));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n18931));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n18930));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n18929));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13765_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[3] [0]), 
            .I3(\Ki[0] ), .O(n18797));   // verilog/coms.v(258[9] 260[65])
    defparam i13765_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13768_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[1] [0]), 
            .I3(control_mode[0]), .O(n18800));   // verilog/coms.v(258[9] 260[65])
    defparam i13768_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 add_624_5_lut (.I0(n10308), .I1(byte_transmit_counter[3]), .I2(GND_net), 
            .I3(n30335), .O(n42881)) /* synthesis syn_instantiated=1 */ ;
    defparam add_624_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13769_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[7] [0]), 
            .I3(PWMLimit[0]), .O(n18801));   // verilog/coms.v(258[9] 260[65])
    defparam i13769_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13883_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[10] [1]), 
            .I3(IntegralLimit[1]), .O(n18915));   // verilog/coms.v(258[9] 260[65])
    defparam i13883_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n18928));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n18927));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n18926));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1035 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17482));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1035.LUT_INIT = 16'h6666;
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n18925));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13884_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[10] [2]), 
            .I3(IntegralLimit[2]), .O(n18916));   // verilog/coms.v(258[9] 260[65])
    defparam i13884_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n18924));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n18923));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n18922));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13885_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[10] [3]), 
            .I3(IntegralLimit[3]), .O(n18917));   // verilog/coms.v(258[9] 260[65])
    defparam i13885_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n18921));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n18920));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n18919));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13886_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[10] [4]), 
            .I3(IntegralLimit[4]), .O(n18918));   // verilog/coms.v(258[9] 260[65])
    defparam i13886_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13887_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[10] [5]), 
            .I3(IntegralLimit[5]), .O(n18919));   // verilog/coms.v(258[9] 260[65])
    defparam i13887_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n18918));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n18917));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n18916));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n18915));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13888_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[10] [6]), 
            .I3(IntegralLimit[6]), .O(n18920));   // verilog/coms.v(258[9] 260[65])
    defparam i13888_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13889_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[10] [7]), 
            .I3(IntegralLimit[7]), .O(n18921));   // verilog/coms.v(258[9] 260[65])
    defparam i13889_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(clk32MHz), 
           .D(n18914));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(clk32MHz), 
           .D(n18913));   // verilog/coms.v(126[12] 289[6])
    SB_DFF byte_transmit_counter_i0_i2 (.Q(byte_transmit_counter[2]), .C(clk32MHz), 
           .D(n36219));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13890_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[9] [0]), 
            .I3(IntegralLimit[8]), .O(n18922));   // verilog/coms.v(258[9] 260[65])
    defparam i13890_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(clk32MHz), 
           .D(n36213));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13891_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[9] [1]), 
            .I3(IntegralLimit[9]), .O(n18923));   // verilog/coms.v(258[9] 260[65])
    defparam i13891_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_out_frame_0___i2 (.Q(\data_out_frame[0] [1]), .C(clk32MHz), 
           .D(n18910));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13892_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[9] [2]), 
            .I3(IntegralLimit[10]), .O(n18924));   // verilog/coms.v(258[9] 260[65])
    defparam i13892_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13893_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[9] [3]), 
            .I3(IntegralLimit[11]), .O(n18925));   // verilog/coms.v(258[9] 260[65])
    defparam i13893_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13894_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[9] [4]), 
            .I3(IntegralLimit[12]), .O(n18926));   // verilog/coms.v(258[9] 260[65])
    defparam i13894_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13895_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[9] [5]), 
            .I3(IntegralLimit[13]), .O(n18927));   // verilog/coms.v(258[9] 260[65])
    defparam i13895_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1036 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[4] [0]), .I3(n37860), .O(n18119));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_4_lut_adj_1036.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1037 (.I0(\FRAME_MATCHER.state_31__N_2492 [3]), .I1(n6121), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n14536));
    defparam i2_3_lut_adj_1037.LUT_INIT = 16'h0808;
    SB_CARRY add_624_5 (.CI(n30335), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n30336));
    SB_LUT4 i14168_3_lut_4_lut (.I0(n8_adj_3912), .I1(n37361), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n19200));
    defparam i14168_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13896_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[9] [6]), 
            .I3(IntegralLimit[14]), .O(n18928));   // verilog/coms.v(258[9] 260[65])
    defparam i13896_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13897_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[9] [7]), 
            .I3(IntegralLimit[15]), .O(n18929));   // verilog/coms.v(258[9] 260[65])
    defparam i13897_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE data_out_frame_0___i3 (.Q(\data_out_frame[0] [2]), .C(clk32MHz), 
            .E(VCC_net), .D(n18850));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i14161_3_lut_4_lut (.I0(n8_adj_3912), .I1(n37361), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n19193));
    defparam i14161_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13898_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[8] [0]), 
            .I3(IntegralLimit[16]), .O(n18930));   // verilog/coms.v(258[9] 260[65])
    defparam i13898_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13899_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[8] [1]), 
            .I3(IntegralLimit[17]), .O(n18931));   // verilog/coms.v(258[9] 260[65])
    defparam i13899_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14162_3_lut_4_lut (.I0(n8_adj_3912), .I1(n37361), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n19194));
    defparam i14162_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13900_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[8] [2]), 
            .I3(IntegralLimit[18]), .O(n18932));   // verilog/coms.v(258[9] 260[65])
    defparam i13900_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14163_3_lut_4_lut (.I0(n8_adj_3912), .I1(n37361), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n19195));
    defparam i14163_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_624_4_lut (.I0(n10308), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(n30334), .O(n42974)) /* synthesis syn_instantiated=1 */ ;
    defparam add_624_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13901_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[8] [3]), 
            .I3(IntegralLimit[19]), .O(n18933));   // verilog/coms.v(258[9] 260[65])
    defparam i13901_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13902_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[8] [4]), 
            .I3(IntegralLimit[20]), .O(n18934));   // verilog/coms.v(258[9] 260[65])
    defparam i13902_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14164_3_lut_4_lut (.I0(n8_adj_3912), .I1(n37361), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n19196));
    defparam i14164_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13903_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[8] [5]), 
            .I3(IntegralLimit[21]), .O(n18935));   // verilog/coms.v(258[9] 260[65])
    defparam i13903_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i22108_1_lut (.I0(n27114), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1972));
    defparam i22108_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13904_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[8] [6]), 
            .I3(IntegralLimit[22]), .O(n18936));   // verilog/coms.v(258[9] 260[65])
    defparam i13904_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13905_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[8] [7]), 
            .I3(IntegralLimit[23]), .O(n18937));   // verilog/coms.v(258[9] 260[65])
    defparam i13905_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14165_3_lut_4_lut (.I0(n8_adj_3912), .I1(n37361), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n19197));
    defparam i14165_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14166_3_lut_4_lut (.I0(n8_adj_3912), .I1(n37361), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n19198));
    defparam i14166_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13912_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[19] [1]), 
            .I3(gearBoxRatio[1]), .O(n18944));   // verilog/coms.v(258[9] 260[65])
    defparam i13912_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13913_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[19] [2]), 
            .I3(gearBoxRatio[2]), .O(n18945));   // verilog/coms.v(258[9] 260[65])
    defparam i13913_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2004_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(\FRAME_MATCHER.i [4]), .O(n10_adj_3982));
    defparam i2004_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i13940_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[2] [6]), 
            .I3(\Kp[6] ), .O(n18972));   // verilog/coms.v(258[9] 260[65])
    defparam i13940_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i21401_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n17031), .I3(\FRAME_MATCHER.i [31]), .O(n2857));
    defparam i21401_3_lut_4_lut.LUT_INIT = 16'h00f8;
    SB_LUT4 i13939_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[2] [5]), 
            .I3(\Kp[5] ), .O(n18971));   // verilog/coms.v(258[9] 260[65])
    defparam i13939_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 equal_105_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3912));
    defparam equal_105_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1038 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n37361), .I3(\FRAME_MATCHER.i [0]), .O(n37368));
    defparam i1_2_lut_3_lut_4_lut_adj_1038.LUT_INIT = 16'hf7ff;
    SB_LUT4 i13938_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[2] [4]), 
            .I3(\Kp[4] ), .O(n18970));   // verilog/coms.v(258[9] 260[65])
    defparam i13938_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13937_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[2] [3]), 
            .I3(\Kp[3] ), .O(n18969));   // verilog/coms.v(258[9] 260[65])
    defparam i13937_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1039 (.I0(\FRAME_MATCHER.state [2]), .I1(n17045), 
            .I2(GND_net), .I3(GND_net), .O(n17025));   // verilog/coms.v(244[5:25])
    defparam i1_2_lut_adj_1039.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1040 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n17183));   // verilog/coms.v(216[5:21])
    defparam i1_2_lut_adj_1040.LUT_INIT = 16'hbbbb;
    SB_LUT4 i17_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n164));   // verilog/coms.v(153[9:50])
    defparam i17_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_4_lut_adj_1041 (.I0(n17264), .I1(n17183), .I2(\FRAME_MATCHER.state [1]), 
            .I3(n17045), .O(n27114));
    defparam i2_4_lut_adj_1041.LUT_INIT = 16'haaa8;
    SB_LUT4 i1_2_lut_adj_1042 (.I0(\data_in_frame[14] [4]), .I1(n33852), 
            .I2(GND_net), .I3(GND_net), .O(n37476));
    defparam i1_2_lut_adj_1042.LUT_INIT = 16'h9999;
    SB_LUT4 i13936_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[2] [2]), 
            .I3(\Kp[2] ), .O(n18968));   // verilog/coms.v(258[9] 260[65])
    defparam i13936_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_adj_1043 (.I0(n18122), .I1(n17874), .I2(Kp_23__N_1353), 
            .I3(GND_net), .O(n37610));
    defparam i2_3_lut_adj_1043.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1044 (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[16] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n17778));   // verilog/coms.v(83[17:63])
    defparam i1_2_lut_adj_1044.LUT_INIT = 16'h6666;
    SB_LUT4 data_in_frame_16__7__I_0_3250_2_lut (.I0(\data_in_frame[16] [7]), 
            .I1(\data_in_frame[16] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1372));   // verilog/coms.v(76[16:27])
    defparam data_in_frame_16__7__I_0_3250_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1045 (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[17] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n37881));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_adj_1045.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1046 (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n18155));
    defparam i1_2_lut_adj_1046.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1047 (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[17] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n37723));
    defparam i1_2_lut_adj_1047.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1048 (.I0(\data_in_frame[1] [3]), .I1(n37795), 
            .I2(\data_in_frame[3] [4]), .I3(GND_net), .O(n17500));   // verilog/coms.v(71[16:34])
    defparam i2_3_lut_adj_1048.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1049 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n37893));
    defparam i1_2_lut_adj_1049.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1050 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[10] [4]), 
            .I2(\data_in_frame[10] [5]), .I3(GND_net), .O(n37848));   // verilog/coms.v(70[16:41])
    defparam i2_3_lut_adj_1050.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1051 (.I0(n17500), .I1(\data_in_frame[7] [7]), 
            .I2(\data_in_frame[10] [3]), .I3(GND_net), .O(n37950));   // verilog/coms.v(71[16:42])
    defparam i2_3_lut_adj_1051.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1052 (.I0(n37950), .I1(n37436), .I2(n37848), 
            .I3(\data_in_frame[12] [7]), .O(n14_adj_3983));   // verilog/coms.v(70[16:41])
    defparam i6_4_lut_adj_1052.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1053 (.I0(n17418), .I1(n14_adj_3983), .I2(n10_adj_3984), 
            .I3(n37594), .O(n17445));   // verilog/coms.v(70[16:41])
    defparam i7_4_lut_adj_1053.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1054 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[10] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n37769));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1054.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1055 (.I0(\data_in_frame[13] [1]), .I1(\data_in_frame[11] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n37980));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1055.LUT_INIT = 16'h6666;
    SB_LUT4 i8_4_lut_adj_1056 (.I0(n37845), .I1(\data_in_frame[17] [2]), 
            .I2(n17418), .I3(n37947), .O(n20_adj_3985));   // verilog/coms.v(69[16:27])
    defparam i8_4_lut_adj_1056.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1057 (.I0(\data_in_frame[19] [4]), .I1(n37980), 
            .I2(n37430), .I3(\data_in_frame[17] [3]), .O(n19_adj_3986));   // verilog/coms.v(69[16:27])
    defparam i7_4_lut_adj_1057.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1058 (.I0(n37769), .I1(n17696), .I2(n17492), 
            .I3(\data_in_frame[15] [2]), .O(n21));   // verilog/coms.v(69[16:27])
    defparam i9_4_lut_adj_1058.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1059 (.I0(\data_in[2] [6]), .I1(\data_in[1] [2]), 
            .I2(n17222), .I3(\data_in[3] [2]), .O(n18_adj_3987));
    defparam i7_4_lut_adj_1059.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_1060 (.I0(\data_in[1] [6]), .I1(n18_adj_3987), 
            .I2(\data_in[1] [3]), .I3(\data_in[2] [0]), .O(n20_adj_3988));
    defparam i9_4_lut_adj_1060.LUT_INIT = 16'hfffd;
    SB_LUT4 i13935_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[2] [1]), 
            .I3(\Kp[1] ), .O(n18967));   // verilog/coms.v(258[9] 260[65])
    defparam i13935_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1061 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n37342), .I3(\FRAME_MATCHER.i [0]), .O(n37348));
    defparam i1_2_lut_3_lut_4_lut_adj_1061.LUT_INIT = 16'hf7ff;
    SB_LUT4 i13934_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[17] [7]), 
            .I3(gearBoxRatio[23]), .O(n18966));   // verilog/coms.v(258[9] 260[65])
    defparam i13934_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i11_3_lut (.I0(n21), .I1(n19_adj_3986), .I2(n20_adj_3985), 
            .I3(GND_net), .O(n37866));   // verilog/coms.v(69[16:27])
    defparam i11_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1062 (.I0(\data_in_frame[19] [5]), .I1(n17445), 
            .I2(\data_in_frame[17] [3]), .I3(GND_net), .O(n37830));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_adj_1062.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1063 (.I0(n37830), .I1(n37866), .I2(\data_in_frame[15] [3]), 
            .I3(GND_net), .O(n37401));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_adj_1063.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1064 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[12] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3989));
    defparam i1_2_lut_adj_1064.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1065 (.I0(n17687), .I1(n37436), .I2(\data_in_frame[10] [2]), 
            .I3(GND_net), .O(n37929));
    defparam i2_3_lut_adj_1065.LUT_INIT = 16'h9696;
    SB_LUT4 data_in_frame_7__7__I_0_2_lut (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[7] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1083));   // verilog/coms.v(83[17:28])
    defparam data_in_frame_7__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1066 (.I0(\data_in_frame[10] [1]), .I1(\data_in_frame[7] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n37783));
    defparam i1_2_lut_adj_1066.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1067 (.I0(n37783), .I1(Kp_23__N_1083), .I2(n37929), 
            .I3(n5_adj_3989), .O(n37536));
    defparam i4_4_lut_adj_1067.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1068 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n37905));
    defparam i1_2_lut_adj_1068.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1069 (.I0(n17449), .I1(\data_in_frame[7] [4]), 
            .I2(n37780), .I3(n6_adj_3990), .O(n33852));
    defparam i4_4_lut_adj_1069.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1070 (.I0(\data_in_frame[14] [4]), .I1(\data_in_frame[14] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n37690));
    defparam i1_2_lut_adj_1070.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1071 (.I0(n37729), .I1(\data_in_frame[10] [1]), 
            .I2(n17449), .I3(n37908), .O(n10_adj_3991));
    defparam i4_4_lut_adj_1071.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1072 (.I0(n17696), .I1(n37536), .I2(GND_net), 
            .I3(GND_net), .O(n18006));
    defparam i1_2_lut_adj_1072.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1073 (.I0(n37914), .I1(n17482), .I2(n37747), 
            .I3(n17449), .O(n14_adj_3992));   // verilog/coms.v(94[12:25])
    defparam i6_4_lut_adj_1073.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1074 (.I0(\data_in_frame[6] [1]), .I1(n14_adj_3992), 
            .I2(n10_adj_3993), .I3(\data_in_frame[1] [6]), .O(n17696));   // verilog/coms.v(94[12:25])
    defparam i7_4_lut_adj_1074.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1075 (.I0(n17696), .I1(\data_in_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n37878));
    defparam i1_2_lut_adj_1075.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1076 (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[6] [1]), 
            .I2(\data_in_frame[16] [7]), .I3(n17425), .O(n15_adj_3994));   // verilog/coms.v(71[16:42])
    defparam i6_4_lut_adj_1076.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1077 (.I0(n15_adj_3994), .I1(n37950), .I2(n14_adj_3995), 
            .I3(n37597), .O(n37661));   // verilog/coms.v(71[16:42])
    defparam i8_4_lut_adj_1077.LUT_INIT = 16'h6996;
    SB_LUT4 i13933_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[17] [6]), 
            .I3(gearBoxRatio[22]), .O(n18965));   // verilog/coms.v(258[9] 260[65])
    defparam i13933_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13932_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[17] [5]), 
            .I3(gearBoxRatio[21]), .O(n18964));   // verilog/coms.v(258[9] 260[65])
    defparam i13932_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1078 (.I0(\data_in_frame[19] [1]), .I1(n37956), 
            .I2(n37661), .I3(\data_in_frame[18] [7]), .O(n10_adj_3996));
    defparam i4_4_lut_adj_1078.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1079 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[1] [0]), .I3(GND_net), .O(n15612));   // verilog/coms.v(94[12:25])
    defparam i2_3_lut_adj_1079.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1080 (.I0(\data_in_frame[1] [1]), .I1(\data_in_frame[3] [3]), 
            .I2(\data_in_frame[0] [7]), .I3(GND_net), .O(n37463));   // verilog/coms.v(83[17:28])
    defparam i2_3_lut_adj_1080.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1081 (.I0(\data_in_frame[0] [7]), .I1(Kp_23__N_858), 
            .I2(n37526), .I3(GND_net), .O(n37899));   // verilog/coms.v(69[16:69])
    defparam i2_3_lut_adj_1081.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut_adj_1082 (.I0(n37526), .I1(Kp_23__N_893), .I2(n3_adj_3997), 
            .I3(\data_in_frame[0] [3]), .O(n26));   // verilog/coms.v(83[17:28])
    defparam i11_4_lut_adj_1082.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1083 (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n37817), .I3(n17482), .O(n24));   // verilog/coms.v(83[17:28])
    defparam i9_4_lut_adj_1083.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1084 (.I0(n37386), .I1(\data_in_frame[2] [3]), 
            .I2(n37655), .I3(\data_in_frame[1] [5]), .O(n25_adj_3998));   // verilog/coms.v(83[17:28])
    defparam i10_4_lut_adj_1084.LUT_INIT = 16'h6996;
    SB_LUT4 i8_3_lut (.I0(n37463), .I1(n15612), .I2(n37631), .I3(GND_net), 
            .O(n23));   // verilog/coms.v(83[17:28])
    defparam i8_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i14_4_lut (.I0(n23), .I1(n25_adj_3998), .I2(n24), .I3(n26), 
            .O(n37710));   // verilog/coms.v(83[17:28])
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1085 (.I0(n37710), .I1(n37899), .I2(\data_in_frame[5] [1]), 
            .I3(GND_net), .O(n33070));
    defparam i2_3_lut_adj_1085.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1086 (.I0(\data_in_frame[7] [3]), .I1(\data_in_frame[12] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n37983));
    defparam i1_2_lut_adj_1086.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1087 (.I0(n33070), .I1(n33854), .I2(GND_net), 
            .I3(GND_net), .O(n33864));
    defparam i1_2_lut_adj_1087.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut (.I0(\data_in_frame[9] [7]), .I1(n17500), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1088 (.I0(n7), .I1(\data_in_frame[4] [7]), .I2(n33864), 
            .I3(n37983), .O(n37729));
    defparam i4_4_lut_adj_1088.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1089 (.I0(n37989), .I1(\data_in_frame[7] [6]), 
            .I2(n37905), .I3(\data_in_frame[12] [0]), .O(n14_adj_3999));
    defparam i6_4_lut_adj_1089.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1090 (.I0(\data_in_frame[14] [2]), .I1(n14_adj_3999), 
            .I2(n10_adj_4000), .I3(n37729), .O(n39322));
    defparam i7_4_lut_adj_1090.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_18__7__I_0_3252_2_lut (.I0(\data_in_frame[18] [7]), 
            .I1(\data_in_frame[18] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1353));   // verilog/coms.v(76[16:27])
    defparam data_in_frame_18__7__I_0_3252_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13931_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[17] [4]), 
            .I3(gearBoxRatio[20]), .O(n18963));   // verilog/coms.v(258[9] 260[65])
    defparam i13931_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13930_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[17] [3]), 
            .I3(gearBoxRatio[19]), .O(n18962));   // verilog/coms.v(258[9] 260[65])
    defparam i13930_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i17_4_lut_adj_1091 (.I0(n37769), .I1(n37795), .I2(\data_in_frame[7] [2]), 
            .I3(n37616), .O(n48_adj_4001));
    defparam i17_4_lut_adj_1091.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut_adj_1092 (.I0(n33886), .I1(\data_in_frame[6] [4]), 
            .I2(\data_in_frame[8] [0]), .I3(n17687), .O(n54_adj_4002));
    defparam i23_4_lut_adj_1092.LUT_INIT = 16'h9669;
    SB_LUT4 i21_4_lut_adj_1093 (.I0(n37783), .I1(n37747), .I2(n37773), 
            .I3(n37693), .O(n52_adj_4003));
    defparam i21_4_lut_adj_1093.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut_adj_1094 (.I0(n37597), .I1(\data_in_frame[2] [1]), 
            .I2(n37470), .I3(Kp_23__N_893), .O(n53_adj_4004));
    defparam i22_4_lut_adj_1094.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut_adj_1095 (.I0(\data_in_frame[9] [4]), .I1(n37887), 
            .I2(n37983), .I3(n37848), .O(n51_adj_4005));
    defparam i20_4_lut_adj_1095.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_1096 (.I0(n37714), .I1(\data_in_frame[5] [7]), 
            .I2(n37533), .I3(\data_in_frame[4] [1]), .O(n50_adj_4006));
    defparam i19_4_lut_adj_1096.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1097 (.I0(n33854), .I1(n37875), .I2(Kp_23__N_760), 
            .I3(n37780), .O(n49_adj_4007));
    defparam i18_4_lut_adj_1097.LUT_INIT = 16'h9669;
    SB_LUT4 i29_4_lut_adj_1098 (.I0(n51_adj_4005), .I1(n53_adj_4004), .I2(n52_adj_4003), 
            .I3(n54_adj_4002), .O(n60_adj_4008));
    defparam i29_4_lut_adj_1098.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut_adj_1099 (.I0(n5_adj_4009), .I1(n48_adj_4001), .I2(n37959), 
            .I3(n37433), .O(n55_adj_4010));
    defparam i24_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut_adj_1100 (.I0(n55_adj_4010), .I1(n60_adj_4008), .I2(n49_adj_4007), 
            .I3(n50_adj_4006), .O(n39467));
    defparam i30_4_lut_adj_1100.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1101 (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[17] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n37917));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1101.LUT_INIT = 16'h6666;
    SB_LUT4 i17_4_lut_adj_1102 (.I0(\data_in_frame[18] [3]), .I1(n37917), 
            .I2(Kp_23__N_1372), .I3(\data_in_frame[17] [0]), .O(n42));
    defparam i17_4_lut_adj_1102.LUT_INIT = 16'h6996;
    SB_LUT4 i6_3_lut (.I0(\data_in_frame[18] [2]), .I1(n33893), .I2(n37953), 
            .I3(GND_net), .O(n31_adj_4011));
    defparam i6_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i12_4_lut_adj_1103 (.I0(\data_in_frame[13] [4]), .I1(Kp_23__N_1406), 
            .I2(n39467), .I3(\data_in_frame[15] [6]), .O(n28_adj_4012));
    defparam i12_4_lut_adj_1103.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_1104 (.I0(n37968), .I1(\data_in_frame[13] [0]), 
            .I2(\data_in_frame[13] [3]), .I3(\data_in_frame[14] [2]), .O(n26_adj_4013));
    defparam i10_4_lut_adj_1104.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1105 (.I0(n37974), .I1(n37443), .I2(n37893), 
            .I3(\data_in_frame[14] [1]), .O(n27_adj_4014));
    defparam i11_4_lut_adj_1105.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1106 (.I0(n18006), .I1(n37690), .I2(\data_in_frame[13] [2]), 
            .I3(\data_in_frame[13] [1]), .O(n25_adj_4015));
    defparam i9_4_lut_adj_1106.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1107 (.I0(n37738), .I1(n37643), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4016));
    defparam i1_2_lut_adj_1107.LUT_INIT = 16'h6666;
    SB_LUT4 i15_4_lut (.I0(n25_adj_4015), .I1(n27_adj_4014), .I2(n26_adj_4013), 
            .I3(n28_adj_4012), .O(n39193));
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut (.I0(n37545), .I1(n37555), .I2(n37820), .I3(GND_net), 
            .O(n28_adj_4017));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i15_4_lut_adj_1108 (.I0(\data_in_frame[15] [2]), .I1(\data_in_frame[17] [5]), 
            .I2(\data_in_frame[17] [3]), .I3(Kp_23__N_1353), .O(n40_c));
    defparam i15_4_lut_adj_1108.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut_adj_1109 (.I0(n31_adj_4011), .I1(n42), .I2(n37726), 
            .I3(n37517), .O(n46_adj_4018));
    defparam i21_4_lut_adj_1109.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_1110 (.I0(n37723), .I1(n39193), .I2(n18155), 
            .I3(n26_adj_4016), .O(n44));
    defparam i19_4_lut_adj_1110.LUT_INIT = 16'h9669;
    SB_LUT4 i20_4_lut_adj_1111 (.I0(\data_in_frame[19] [7]), .I1(n40_c), 
            .I2(n28_adj_4017), .I3(n37401), .O(n45));
    defparam i20_4_lut_adj_1111.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1112 (.I0(n37760), .I1(n37956), .I2(\data_in_frame[16] [0]), 
            .I3(n37881), .O(n43));
    defparam i18_4_lut_adj_1112.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut_adj_1113 (.I0(n43), .I1(n45), .I2(n44), .I3(n46_adj_4018), 
            .O(n37669));
    defparam i24_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1114 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n37383));   // verilog/coms.v(94[12:25])
    defparam i1_2_lut_adj_1114.LUT_INIT = 16'h6666;
    SB_LUT4 i13929_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[17] [2]), 
            .I3(gearBoxRatio[18]), .O(n18961));   // verilog/coms.v(258[9] 260[65])
    defparam i13929_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13928_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[17] [1]), 
            .I3(gearBoxRatio[17]), .O(n18960));   // verilog/coms.v(258[9] 260[65])
    defparam i13928_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13927_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[17] [0]), 
            .I3(gearBoxRatio[16]), .O(n18959));   // verilog/coms.v(258[9] 260[65])
    defparam i13927_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13926_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[18] [7]), 
            .I3(gearBoxRatio[15]), .O(n18958));   // verilog/coms.v(258[9] 260[65])
    defparam i13926_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_2_lut (.I0(\data_in[2] [5]), .I1(\data_in[0] [1]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4019));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_adj_1115 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [4]), .I3(GND_net), .O(n6_adj_4020));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_1115.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1116 (.I0(\data_in_frame[9] [0]), .I1(n17844), 
            .I2(GND_net), .I3(GND_net), .O(n37926));   // verilog/coms.v(76[16:50])
    defparam i1_2_lut_adj_1116.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1117 (.I0(Kp_23__N_893), .I1(\data_in_frame[7] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n17827));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1117.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1118 (.I0(\data_in_frame[11] [2]), .I1(\data_in_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n37773));   // verilog/coms.v(76[16:50])
    defparam i1_2_lut_adj_1118.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1119 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[8] [6]), 
            .I2(\data_in_frame[6] [5]), .I3(GND_net), .O(n37430));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut_adj_1119.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1120 (.I0(\data_in_frame[9] [5]), .I1(n37902), 
            .I2(n37714), .I3(n33864), .O(n33843));
    defparam i3_4_lut_adj_1120.LUT_INIT = 16'h9669;
    SB_LUT4 i13925_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[18] [6]), 
            .I3(gearBoxRatio[14]), .O(n18957));   // verilog/coms.v(258[9] 260[65])
    defparam i13925_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 data_in_frame_13__7__I_0_2_lut (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1406));   // verilog/coms.v(68[16:27])
    defparam data_in_frame_13__7__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1121 (.I0(\data_in_frame[13] [5]), .I1(\data_in_frame[15] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n18228));
    defparam i1_2_lut_adj_1121.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1122 (.I0(n37430), .I1(n37773), .I2(\data_in_frame[6] [7]), 
            .I3(\data_in_frame[9] [1]), .O(n12_adj_4021));   // verilog/coms.v(76[16:50])
    defparam i5_4_lut_adj_1122.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1123 (.I0(n17827), .I1(n12_adj_4021), .I2(n37926), 
            .I3(\data_in_frame[4] [6]), .O(n18091));   // verilog/coms.v(76[16:50])
    defparam i6_4_lut_adj_1123.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1124 (.I0(n18091), .I1(\data_in_frame[16] [1]), 
            .I2(n17379), .I3(n37622), .O(n10_adj_4022));
    defparam i4_4_lut_adj_1124.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1125 (.I0(\data_in_frame[16] [0]), .I1(n10_adj_4022), 
            .I2(\data_in_frame[14] [0]), .I3(GND_net), .O(n33893));
    defparam i5_3_lut_adj_1125.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1126 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n37511));   // verilog/coms.v(230[9:81])
    defparam i1_2_lut_adj_1126.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1127 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[3] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n37631));   // verilog/coms.v(230[9:81])
    defparam i1_2_lut_adj_1127.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1128 (.I0(\data_in_frame[4] [3]), .I1(n37511), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[2] [1]), .O(n17863));   // verilog/coms.v(230[9:81])
    defparam i3_4_lut_adj_1128.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1129 (.I0(\data_in_frame[4] [1]), .I1(n37631), 
            .I2(\data_in_frame[1] [7]), .I3(\data_in_frame[2] [0]), .O(n17425));   // verilog/coms.v(230[9:81])
    defparam i3_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1130 (.I0(\data_in_frame[5] [7]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[1] [5]), .O(n37564));   // verilog/coms.v(94[12:25])
    defparam i3_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1131 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1] [2]), .I3(GND_net), .O(n37567));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1131.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1132 (.I0(\data_in_frame[8] [3]), .I1(\data_in_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n37851));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_1132.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1133 (.I0(n37567), .I1(n37776), .I2(\data_in_frame[6] [0]), 
            .I3(n37564), .O(n12_adj_4023));   // verilog/coms.v(74[16:43])
    defparam i5_4_lut_adj_1133.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1134 (.I0(\data_in_frame[8] [2]), .I1(n12_adj_4023), 
            .I2(n37851), .I3(\data_in_frame[3] [4]), .O(n17559));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_1134.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1135 (.I0(\data_in_frame[6] [4]), .I1(n17425), 
            .I2(n17863), .I3(\data_in_frame[8] [5]), .O(n37594));   // verilog/coms.v(69[16:27])
    defparam i3_4_lut_adj_1135.LUT_INIT = 16'h6996;
    SB_LUT4 i13924_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[18] [5]), 
            .I3(gearBoxRatio[13]), .O(n18956));   // verilog/coms.v(258[9] 260[65])
    defparam i13924_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13923_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[18] [4]), 
            .I3(gearBoxRatio[12]), .O(n18955));   // verilog/coms.v(258[9] 260[65])
    defparam i13923_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13922_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[18] [3]), 
            .I3(gearBoxRatio[11]), .O(n18954));   // verilog/coms.v(258[9] 260[65])
    defparam i13922_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13921_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[18] [2]), 
            .I3(gearBoxRatio[10]), .O(n18953));   // verilog/coms.v(258[9] 260[65])
    defparam i13921_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i10_4_lut_adj_1136 (.I0(n15_adj_4019), .I1(n20_adj_3988), .I2(\data_in[0] [5]), 
            .I3(\data_in[3] [7]), .O(n17055));
    defparam i10_4_lut_adj_1136.LUT_INIT = 16'hfeff;
    SB_LUT4 i13920_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[18] [1]), 
            .I3(gearBoxRatio[9]), .O(n18952));   // verilog/coms.v(258[9] 260[65])
    defparam i13920_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13919_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[18] [0]), 
            .I3(gearBoxRatio[8]), .O(n18951));   // verilog/coms.v(258[9] 260[65])
    defparam i13919_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13918_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[19] [7]), 
            .I3(gearBoxRatio[7]), .O(n18950));   // verilog/coms.v(258[9] 260[65])
    defparam i13918_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13947_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[3] [6]), 
            .I3(\Ki[6] ), .O(n18979));   // verilog/coms.v(258[9] 260[65])
    defparam i13947_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13946_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[3] [5]), 
            .I3(\Ki[5] ), .O(n18978));   // verilog/coms.v(258[9] 260[65])
    defparam i13946_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_CARRY add_624_4 (.CI(n30334), .I0(byte_transmit_counter[2]), .I1(GND_net), 
            .CO(n30335));
    SB_LUT4 i1_2_lut_4_lut_adj_1137 (.I0(n326), .I1(n200), .I2(n324), 
            .I3(\FRAME_MATCHER.state [31]), .O(n8_adj_4024));
    defparam i1_2_lut_4_lut_adj_1137.LUT_INIT = 16'hfe00;
    SB_LUT4 i13945_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[3] [4]), 
            .I3(\Ki[4] ), .O(n18977));   // verilog/coms.v(258[9] 260[65])
    defparam i13945_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13944_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[3] [3]), 
            .I3(\Ki[3] ), .O(n18976));   // verilog/coms.v(258[9] 260[65])
    defparam i13944_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13943_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[3] [2]), 
            .I3(\Ki[2] ), .O(n18975));   // verilog/coms.v(258[9] 260[65])
    defparam i13943_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13942_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[3] [1]), 
            .I3(\Ki[1] ), .O(n18974));   // verilog/coms.v(258[9] 260[65])
    defparam i13942_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_1138 (.I0(\data_in_frame[18] [7]), .I1(n12_adj_4025), 
            .I2(n37669), .I3(n18122), .O(n38781));
    defparam i6_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1139 (.I0(\data_in_frame[21] [3]), .I1(n37545), 
            .I2(n37820), .I3(GND_net), .O(n37939));
    defparam i1_3_lut_adj_1139.LUT_INIT = 16'h9696;
    SB_LUT4 i9_4_lut_adj_1140 (.I0(n17_adj_4026), .I1(\data_in_frame[17] [6]), 
            .I2(n16_adj_4027), .I3(\data_in_frame[20] [2]), .O(n39117));
    defparam i9_4_lut_adj_1140.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1141 (.I0(n37643), .I1(n38588), .I2(n37820), 
            .I3(\data_in_frame[21] [4]), .O(n22));
    defparam i6_4_lut_adj_1141.LUT_INIT = 16'hb77b;
    SB_LUT4 i33763_4_lut (.I0(n37939), .I1(n38781), .I2(n38719), .I3(n39798), 
            .O(n40829));
    defparam i33763_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i6_4_lut_adj_1142 (.I0(n17167), .I1(\data_in[3] [3]), .I2(\data_in[2] [1]), 
            .I3(\data_in[3] [6]), .O(n16_adj_4028));
    defparam i6_4_lut_adj_1142.LUT_INIT = 16'hffbf;
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_3971), .S(n3_adj_4029));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13941_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[2] [7]), 
            .I3(\Kp[7] ), .O(n18973));   // verilog/coms.v(258[9] 260[65])
    defparam i13941_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_3966), .S(n3_adj_4030));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i14312_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[6] [5]), 
            .I3(PWMLimit[13]), .O(n19344));   // verilog/coms.v(258[9] 260[65])
    defparam i14312_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14311_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[6] [4]), 
            .I3(PWMLimit[12]), .O(n19343));   // verilog/coms.v(258[9] 260[65])
    defparam i14311_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14310_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[6] [3]), 
            .I3(PWMLimit[11]), .O(n19342));   // verilog/coms.v(258[9] 260[65])
    defparam i14310_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14309_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[6] [2]), 
            .I3(PWMLimit[10]), .O(n19341));   // verilog/coms.v(258[9] 260[65])
    defparam i14309_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7_4_lut_adj_1143 (.I0(\data_in[2] [3]), .I1(n17055), .I2(\data_in[3] [5]), 
            .I3(\data_in[0] [7]), .O(n17_adj_4031));
    defparam i7_4_lut_adj_1143.LUT_INIT = 16'hffdf;
    SB_LUT4 i14308_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[6] [1]), 
            .I3(PWMLimit[9]), .O(n19340));   // verilog/coms.v(258[9] 260[65])
    defparam i14308_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14307_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[6] [0]), 
            .I3(PWMLimit[8]), .O(n19339));   // verilog/coms.v(258[9] 260[65])
    defparam i14307_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14306_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[7] [7]), 
            .I3(PWMLimit[7]), .O(n19338));   // verilog/coms.v(258[9] 260[65])
    defparam i14306_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_3960), .S(n3_adj_4032));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_3959), .S(n3_adj_4033));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2_adj_3954), .S(n3_adj_4034));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_3951), .S(n3_adj_4035));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_3941), .S(n3_adj_4036));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_3934), .S(n3_adj_4037));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_3929), .S(n3_adj_4038));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_3928), .S(n3_adj_4039));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_3917), .S(n3_adj_4040));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_3914), .S(n3_adj_4041));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_3913), .S(n3_adj_4042));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_3905), .S(n3_adj_4043));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_3904), .S(n3_adj_4044));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_3903), .S(n3_adj_4045));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2), .S(n3_adj_4046));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_4047), .S(n3_adj_4048));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_4049), .S(n3_adj_4050));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_4051), .S(n3_adj_4052));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_4053), .S(n3_adj_4054));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_4055), .S(n3_adj_4056));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_4057), .S(n3_adj_4058));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_4059), .S(n3_adj_4060));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_4061), .S(n3_adj_4062));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_4063), .S(n3_adj_4064));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_4065), .S(n3_adj_4066));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_4067), .S(n3_adj_4068));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_4069), .S(n3_adj_4070));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_4071), .S(n3_adj_4072));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_4073), .S(n3_adj_4074));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk32MHz), 
            .E(n18436), .D(n38745));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i14305_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[7] [6]), 
            .I3(PWMLimit[6]), .O(n19337));   // verilog/coms.v(258[9] 260[65])
    defparam i14305_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1144 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [6]), .I3(n37561), .O(n18143));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(byte_transmit_counter[1]), .O(n46028));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i14304_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[7] [5]), 
            .I3(PWMLimit[5]), .O(n19336));   // verilog/coms.v(258[9] 260[65])
    defparam i14304_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFFE data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk32MHz), 
            .E(n18436), .D(n38514));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk32MHz), 
            .E(n18436), .D(n39012));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk32MHz), 
            .E(n18436), .D(n38922));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk32MHz), 
            .E(n18436), .D(n37721));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk32MHz), 
            .E(n18436), .D(n38639));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk32MHz), 
            .E(n18436), .D(n38629));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk32MHz), 
            .E(n18436), .D(n38644));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk32MHz), 
            .E(n18436), .D(n38857));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk32MHz), 
            .E(n18436), .D(n37802));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk32MHz), 
            .E(n18436), .D(n37826));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk32MHz), 
            .E(n18436), .D(n37825));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk32MHz), 
            .E(n18436), .D(n37551));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk32MHz), 
            .E(n18436), .D(n17597));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk32MHz), 
            .E(n18436), .D(n38713));   // verilog/coms.v(126[12] 289[6])
    SB_DFFE data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk32MHz), 
            .E(n18436), .D(n39432));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i14303_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[7] [4]), 
            .I3(PWMLimit[4]), .O(n19335));   // verilog/coms.v(258[9] 260[65])
    defparam i14303_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .D(n18829));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state [1]), .C(clk32MHz), 
            .D(n36585), .S(n46228));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state[3] ), .C(clk32MHz), 
            .D(n36589), .S(n36609));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n36783), .S(n36679));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n36787), .S(n36599));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n36791), .S(n36601));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n36795), .S(n36659));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n36799), .S(n36657));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n36803), .S(n36655));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n36811), .S(n36651));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n36815), .S(n36649));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n36819), .S(n36647));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n36823), .S(n36645));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n36827), .S(n36643));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n7_adj_4075), .S(n8_adj_4076));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n36831), .S(n36603));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n7_adj_4077), .S(n8_adj_4078));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n7_adj_4079), .S(n8_adj_4080));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n36751), .S(n36579));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n7_adj_4081), .S(n36683));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n36807), .S(n36653));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n36763), .S(n36641));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n7_adj_4082), .S(n8_adj_4083));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n7_adj_4084), .S(n36639));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n36767), .S(n36693));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n36771), .S(n36637));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n7_adj_4085), .S(n8_adj_4086));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n36775), .S(n36635));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n7_adj_4087), .S(n8_adj_4088));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n36779), .S(n8_adj_4089));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n7_adj_4090), .S(n8_adj_4024));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n19217));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n46028_bdd_4_lut (.I0(n46028), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(byte_transmit_counter[1]), 
            .O(n46031));
    defparam n46028_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 data_in_frame_12__7__I_0_3248_2_lut (.I0(\data_in_frame[12] [7]), 
            .I1(\data_in_frame[12] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_760));   // verilog/coms.v(69[16:27])
    defparam data_in_frame_12__7__I_0_3248_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_38879 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(byte_transmit_counter[1]), .O(n46022));
    defparam byte_transmit_counter_0__bdd_4_lut_38879.LUT_INIT = 16'he4aa;
    SB_LUT4 n46022_bdd_4_lut (.I0(n46022), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(byte_transmit_counter[1]), 
            .O(n46025));
    defparam n46022_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_4_lut_adj_1145 (.I0(Kp_23__N_760), .I1(n37845), .I2(n17418), 
            .I3(n17844), .O(n12_adj_4091));   // verilog/coms.v(69[16:27])
    defparam i5_4_lut_adj_1145.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_38874 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(byte_transmit_counter[1]), .O(n46016));
    defparam byte_transmit_counter_0__bdd_4_lut_38874.LUT_INIT = 16'he4aa;
    SB_LUT4 n46016_bdd_4_lut (.I0(n46016), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(byte_transmit_counter[1]), 
            .O(n46019));
    defparam n46016_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1146 (.I0(n37594), .I1(n12_adj_4091), .I2(n17559), 
            .I3(\data_in_frame[19] [6]), .O(n37754));   // verilog/coms.v(69[16:27])
    defparam i6_4_lut_adj_1146.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_38869 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(byte_transmit_counter[1]), .O(n46010));
    defparam byte_transmit_counter_0__bdd_4_lut_38869.LUT_INIT = 16'he4aa;
    SB_LUT4 n46010_bdd_4_lut (.I0(n46010), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(byte_transmit_counter[1]), 
            .O(n46013));
    defparam n46010_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1147 (.I0(\data_in_frame[8] [6]), .I1(n17863), 
            .I2(GND_net), .I3(GND_net), .O(n37392));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_adj_1147.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_38864 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(byte_transmit_counter[1]), .O(n46004));
    defparam byte_transmit_counter_0__bdd_4_lut_38864.LUT_INIT = 16'he4aa;
    SB_LUT4 n46004_bdd_4_lut (.I0(n46004), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(byte_transmit_counter[1]), 
            .O(n46007));
    defparam n46004_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1148 (.I0(\data_in_frame[6] [4]), .I1(\data_in_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n37896));
    defparam i1_2_lut_adj_1148.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_38859 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(byte_transmit_counter[1]), .O(n45998));
    defparam byte_transmit_counter_0__bdd_4_lut_38859.LUT_INIT = 16'he4aa;
    SB_LUT4 n45998_bdd_4_lut (.I0(n45998), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(byte_transmit_counter[1]), 
            .O(n46001));
    defparam n45998_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut_adj_1149 (.I0(n33886), .I1(\data_in_frame[7] [1]), 
            .I2(n37698), .I3(\data_in_frame[11] [3]), .O(n18_adj_4092));
    defparam i7_4_lut_adj_1149.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_38854 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(byte_transmit_counter[1]), .O(n45992));
    defparam byte_transmit_counter_0__bdd_4_lut_38854.LUT_INIT = 16'he4aa;
    SB_LUT4 n45992_bdd_4_lut (.I0(n45992), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(byte_transmit_counter[1]), 
            .O(n45995));
    defparam n45992_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_2_lut_adj_1150 (.I0(\data_in_frame[7] [0]), .I1(\data_in_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4093));
    defparam i5_2_lut_adj_1150.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_38849 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(byte_transmit_counter[1]), .O(n45986));
    defparam byte_transmit_counter_0__bdd_4_lut_38849.LUT_INIT = 16'he4aa;
    SB_LUT4 i14302_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[7] [3]), 
            .I3(PWMLimit[3]), .O(n19334));   // verilog/coms.v(258[9] 260[65])
    defparam i14302_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14301_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[7] [2]), 
            .I3(PWMLimit[2]), .O(n19333));   // verilog/coms.v(258[9] 260[65])
    defparam i14301_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_adj_1151 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[4] [1]), .I3(GND_net), .O(n18209));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1151.LUT_INIT = 16'h9696;
    SB_LUT4 i14300_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[7] [1]), 
            .I3(PWMLimit[1]), .O(n19332));   // verilog/coms.v(258[9] 260[65])
    defparam i14300_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14299_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[1] [7]), 
            .I3(control_mode[7]), .O(n19331));   // verilog/coms.v(258[9] 260[65])
    defparam i14299_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14298_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[1] [6]), 
            .I3(control_mode[6]), .O(n19330));   // verilog/coms.v(258[9] 260[65])
    defparam i14298_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14297_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[1] [5]), 
            .I3(control_mode[5]), .O(n19329));   // verilog/coms.v(258[9] 260[65])
    defparam i14297_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 n45986_bdd_4_lut (.I0(n45986), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(byte_transmit_counter[1]), 
            .O(n45989));
    defparam n45986_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i9_4_lut_adj_1152 (.I0(n17_adj_4031), .I1(\data_in[0] [2]), 
            .I2(n16_adj_4028), .I3(\data_in[3] [1]), .O(n63_adj_3909));
    defparam i9_4_lut_adj_1152.LUT_INIT = 16'hfbff;
    SB_LUT4 i14296_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[1] [4]), 
            .I3(control_mode[4]), .O(n19328));   // verilog/coms.v(258[9] 260[65])
    defparam i14296_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14295_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[1] [3]), 
            .I3(control_mode[3]), .O(n19327));   // verilog/coms.v(258[9] 260[65])
    defparam i14295_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14294_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[1] [2]), 
            .I3(control_mode[2]), .O(n19326));   // verilog/coms.v(258[9] 260[65])
    defparam i14294_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14289_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[1] [1]), 
            .I3(control_mode[1]), .O(n19321));   // verilog/coms.v(258[9] 260[65])
    defparam i14289_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14322_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[5] [7]), 
            .I3(PWMLimit[23]), .O(n19354));   // verilog/coms.v(258[9] 260[65])
    defparam i14322_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 add_624_3_lut (.I0(n10308), .I1(byte_transmit_counter[1]), .I2(GND_net), 
            .I3(n30333), .O(n42973)) /* synthesis syn_instantiated=1 */ ;
    defparam add_624_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i14153_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37361), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n19185));
    defparam i14153_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14320_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[5] [5]), 
            .I3(PWMLimit[21]), .O(n19352));   // verilog/coms.v(258[9] 260[65])
    defparam i14320_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13948_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[3] [7]), 
            .I3(\Ki[7] ), .O(n18980));   // verilog/coms.v(258[9] 260[65])
    defparam i13948_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14319_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[5] [4]), 
            .I3(PWMLimit[20]), .O(n19351));   // verilog/coms.v(258[9] 260[65])
    defparam i14319_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_1153 (.I0(\data_in[3] [0]), .I1(n17247), .I2(n17055), 
            .I3(\data_in[2] [2]), .O(n16_adj_4094));
    defparam i6_4_lut_adj_1153.LUT_INIT = 16'hfffe;
    SB_LUT4 i14318_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[5] [3]), 
            .I3(PWMLimit[19]), .O(n19350));   // verilog/coms.v(258[9] 260[65])
    defparam i14318_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i7_4_lut_adj_1154 (.I0(\data_in[2] [4]), .I1(\data_in[1] [0]), 
            .I2(\data_in[1] [5]), .I3(\data_in[0] [3]), .O(n17_adj_4095));
    defparam i7_4_lut_adj_1154.LUT_INIT = 16'hfffd;
    SB_LUT4 i14317_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[5] [2]), 
            .I3(PWMLimit[18]), .O(n19349));   // verilog/coms.v(258[9] 260[65])
    defparam i14317_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14154_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37361), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n19186));
    defparam i14154_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14316_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[5] [1]), 
            .I3(PWMLimit[17]), .O(n19348));   // verilog/coms.v(258[9] 260[65])
    defparam i14316_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 add_44_22_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n30321), .O(n2_adj_4051)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_22_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n19216));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_adj_1155 (.I0(\data_in_frame[1] [2]), .I1(n37914), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4009));   // verilog/coms.v(94[12:25])
    defparam i1_2_lut_adj_1155.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1156 (.I0(\data_in_frame[3] [5]), .I1(n37564), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4096));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1156.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n19215));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n19214));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i14315_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[5] [0]), 
            .I3(PWMLimit[16]), .O(n19347));   // verilog/coms.v(258[9] 260[65])
    defparam i14315_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n19213));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(clk32MHz), 
           .D(n19200));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n19212));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n19264));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_624_3 (.CI(n30333), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n30334));
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n19263));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i14314_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[6] [7]), 
            .I3(PWMLimit[15]), .O(n19346));   // verilog/coms.v(258[9] 260[65])
    defparam i14314_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14313_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[6] [6]), 
            .I3(PWMLimit[14]), .O(n19345));   // verilog/coms.v(258[9] 260[65])
    defparam i14313_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9_4_lut_adj_1157 (.I0(\data_in_frame[9] [2]), .I1(n18_adj_4092), 
            .I2(Kp_23__N_820), .I3(n37926), .O(n20_adj_4097));
    defparam i9_4_lut_adj_1157.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_38844 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(byte_transmit_counter[1]), .O(n45980));
    defparam byte_transmit_counter_0__bdd_4_lut_38844.LUT_INIT = 16'he4aa;
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n19262));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n19261));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n19260));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n19259));   // verilog/coms.v(126[12] 289[6])
    SB_DFFSR tx_transmit_3227 (.Q(r_SM_Main_2__N_3323[0]), .C(clk32MHz), 
            .D(n43083), .R(n38178));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n19211));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n19210));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n19209));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n19208));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i13914_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[19] [3]), 
            .I3(gearBoxRatio[3]), .O(n18946));   // verilog/coms.v(258[9] 260[65])
    defparam i13914_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i14155_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37361), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n19187));
    defparam i14155_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13915_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[19] [4]), 
            .I3(gearBoxRatio[4]), .O(n18947));   // verilog/coms.v(258[9] 260[65])
    defparam i13915_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13916_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[19] [5]), 
            .I3(gearBoxRatio[5]), .O(n18948));   // verilog/coms.v(258[9] 260[65])
    defparam i13916_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n19240));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i12_4_lut_adj_1158 (.I0(n17500), .I1(n5_adj_4009), .I2(n17900), 
            .I3(n7_adj_4098), .O(n28_adj_4099));   // verilog/coms.v(230[9:81])
    defparam i12_4_lut_adj_1158.LUT_INIT = 16'hfffd;
    SB_LUT4 i13917_3_lut_4_lut (.I0(Kp_23__N_718), .I1(n63_adj_3981), .I2(\data_in_frame[19] [6]), 
            .I3(gearBoxRatio[6]), .O(n18949));   // verilog/coms.v(258[9] 260[65])
    defparam i13917_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9_4_lut_adj_1159 (.I0(n17_adj_4095), .I1(\data_in[0] [6]), 
            .I2(n16_adj_4094), .I3(\data_in[1] [4]), .O(n63_c));
    defparam i9_4_lut_adj_1159.LUT_INIT = 16'hfbff;
    SB_LUT4 i2_3_lut_adj_1160 (.I0(\data_in_frame[18] [4]), .I1(n37726), 
            .I2(\data_in_frame[20] [6]), .I3(GND_net), .O(n39620));
    defparam i2_3_lut_adj_1160.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1161 (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[20] [0]), 
            .I2(\data_in_frame[17] [4]), .I3(GND_net), .O(n7_adj_4100));   // verilog/coms.v(69[16:27])
    defparam i1_3_lut_adj_1161.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1162 (.I0(n37754), .I1(n7_adj_4100), .I2(\data_in_frame[19] [7]), 
            .I3(n8_adj_4101), .O(n39166));   // verilog/coms.v(69[16:27])
    defparam i5_4_lut_adj_1162.LUT_INIT = 16'h6996;
    SB_LUT4 i21406_4_lut (.I0(n10_adj_3982), .I1(\FRAME_MATCHER.i [31]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(n17208), .O(n3761));   // verilog/coms.v(249[9:58])
    defparam i21406_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i14156_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37361), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n19188));
    defparam i14156_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14157_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37361), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n19189));
    defparam i14157_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21485_2_lut (.I0(byte_transmit_counter[1]), .I1(byte_transmit_counter[2]), 
            .I2(GND_net), .I3(GND_net), .O(n26492));
    defparam i21485_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i14158_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37361), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n19190));
    defparam i14158_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_624_2_lut (.I0(GND_net), .I1(byte_transmit_counter[0]), 
            .I2(tx_transmit_N_3215), .I3(GND_net), .O(n2236[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_624_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_624_2 (.CI(GND_net), .I0(byte_transmit_counter[0]), .I1(tx_transmit_N_3215), 
            .CO(n30333));
    SB_LUT4 i33726_4_lut (.I0(n38953), .I1(n33880), .I2(n10), .I3(n33893), 
            .O(n40790));
    defparam i33726_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i10_4_lut_adj_1163 (.I0(n19_adj_3938), .I1(\data_in_frame[21] [1]), 
            .I2(n38540), .I3(n37669), .O(n26_adj_4102));
    defparam i10_4_lut_adj_1163.LUT_INIT = 16'hbfef;
    SB_LUT4 i14_4_lut_adj_1164 (.I0(n39620), .I1(n40829), .I2(n22), .I3(n39117), 
            .O(n30_adj_4103));
    defparam i14_4_lut_adj_1164.LUT_INIT = 16'hfbff;
    SB_LUT4 i1_4_lut_adj_1165 (.I0(n37610), .I1(n39166), .I2(n37669), 
            .I3(\data_in_frame[21] [0]), .O(n17_adj_4104));
    defparam i1_4_lut_adj_1165.LUT_INIT = 16'hedde;
    SB_LUT4 i10_4_lut_adj_1166 (.I0(n37896), .I1(n20_adj_4097), .I2(n16_adj_4093), 
            .I3(n37392), .O(Kp_23__N_1433));
    defparam i10_4_lut_adj_1166.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1167 (.I0(n17_adj_4104), .I1(n30_adj_4103), .I2(n26_adj_4102), 
            .I3(n40790), .O(n31_adj_4105));
    defparam i15_4_lut_adj_1167.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_adj_1168 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n17833));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1168.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1169 (.I0(byte_transmit_counter[6]), .I1(byte_transmit_counter[5]), 
            .I2(n27441), .I3(byte_transmit_counter[7]), .O(n20_adj_4106));
    defparam i3_4_lut_adj_1169.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1170 (.I0(\FRAME_MATCHER.state [31]), .I1(\FRAME_MATCHER.state [24]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4107));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_adj_1170.LUT_INIT = 16'heeee;
    SB_LUT4 i4_4_lut_adj_1171 (.I0(\FRAME_MATCHER.state [27]), .I1(\FRAME_MATCHER.state [20]), 
            .I2(\FRAME_MATCHER.state [23]), .I3(n6_adj_4107), .O(n33677));   // verilog/coms.v(126[12] 289[6])
    defparam i4_4_lut_adj_1171.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1172 (.I0(\FRAME_MATCHER.state [29]), .I1(\FRAME_MATCHER.state [15]), 
            .I2(\FRAME_MATCHER.state [11]), .I3(\FRAME_MATCHER.state [13]), 
            .O(n30_adj_4108));   // verilog/coms.v(206[5:16])
    defparam i11_4_lut_adj_1172.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1173 (.I0(\FRAME_MATCHER.state [12]), .I1(n30_adj_4108), 
            .I2(\FRAME_MATCHER.state [21]), .I3(\FRAME_MATCHER.state [28]), 
            .O(n34));   // verilog/coms.v(206[5:16])
    defparam i15_4_lut_adj_1173.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1174 (.I0(\FRAME_MATCHER.state [22]), .I1(\FRAME_MATCHER.state [25]), 
            .I2(\FRAME_MATCHER.state [30]), .I3(\FRAME_MATCHER.state [14]), 
            .O(n32));   // verilog/coms.v(206[5:16])
    defparam i13_4_lut_adj_1174.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1175 (.I0(\FRAME_MATCHER.state [18]), .I1(\FRAME_MATCHER.state [16]), 
            .I2(\FRAME_MATCHER.state [9]), .I3(\FRAME_MATCHER.state [17]), 
            .O(n33));   // verilog/coms.v(206[5:16])
    defparam i14_4_lut_adj_1175.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1176 (.I0(n17031), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_4109));
    defparam i1_2_lut_adj_1176.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1177 (.I0(\FRAME_MATCHER.state [19]), .I1(\FRAME_MATCHER.state [8]), 
            .I2(\FRAME_MATCHER.state [10]), .I3(\FRAME_MATCHER.state [26]), 
            .O(n31_adj_4110));   // verilog/coms.v(206[5:16])
    defparam i12_4_lut_adj_1177.LUT_INIT = 16'hfffe;
    SB_LUT4 i21400_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n4_adj_4109), .I3(\FRAME_MATCHER.i [1]), .O(n740));   // verilog/coms.v(157[9:60])
    defparam i21400_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i31032_2_lut (.I0(n17265), .I1(n26317), .I2(GND_net), .I3(GND_net), 
            .O(n38092));
    defparam i31032_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_3_lut_adj_1178 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17199), .I3(GND_net), .O(n17201));   // verilog/coms.v(253[5:27])
    defparam i1_2_lut_3_lut_adj_1178.LUT_INIT = 16'hfefe;
    SB_LUT4 add_44_33_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n30332), .O(n2_adj_4073)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i10_4_lut_adj_1179 (.I0(n17425), .I1(n17687), .I2(n17636), 
            .I3(n33070), .O(n26_adj_4111));   // verilog/coms.v(230[9:81])
    defparam i10_4_lut_adj_1179.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_3_lut_adj_1180 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17266), .I3(GND_net), .O(n63_adj_3981));   // verilog/coms.v(253[5:27])
    defparam i1_2_lut_3_lut_adj_1180.LUT_INIT = 16'hfefe;
    SB_LUT4 i14159_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37361), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n19191));
    defparam i14159_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n19207));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1181 (.I0(\data_in_frame[3] [0]), .I1(n37750), 
            .I2(n37607), .I3(\data_in_frame[2] [6]), .O(n37489));   // verilog/coms.v(69[16:69])
    defparam i1_2_lut_3_lut_4_lut_adj_1181.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n19206));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n19205));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i14160_3_lut_4_lut (.I0(n8_adj_3933), .I1(n37361), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n19192));
    defparam i14160_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n19204));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 equal_106_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3933));   // verilog/coms.v(154[7:23])
    defparam equal_106_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i3_3_lut_adj_1182 (.I0(n63_adj_3981), .I1(n27114), .I2(n17265), 
            .I3(GND_net), .O(n8_adj_4112));
    defparam i3_3_lut_adj_1182.LUT_INIT = 16'h8080;
    SB_LUT4 i4_4_lut_adj_1183 (.I0(n17200), .I1(n8_adj_4112), .I2(n17170), 
            .I3(n17045), .O(n2664));
    defparam i4_4_lut_adj_1183.LUT_INIT = 16'h8880;
    SB_LUT4 i17_4_lut_adj_1184 (.I0(\FRAME_MATCHER.i [17]), .I1(\FRAME_MATCHER.i [26]), 
            .I2(\FRAME_MATCHER.i [14]), .I3(\FRAME_MATCHER.i [23]), .O(n42_adj_4113));
    defparam i17_4_lut_adj_1184.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1185 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [24]), 
            .I2(\FRAME_MATCHER.i [15]), .I3(\FRAME_MATCHER.i [16]), .O(n40_adj_4114));
    defparam i15_4_lut_adj_1185.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1186 (.I0(\FRAME_MATCHER.i [28]), .I1(\FRAME_MATCHER.i [12]), 
            .I2(\FRAME_MATCHER.i [11]), .I3(\FRAME_MATCHER.i [30]), .O(n41));
    defparam i16_4_lut_adj_1186.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1187 (.I0(\FRAME_MATCHER.state [2]), .I1(n17045), 
            .I2(n17263), .I3(GND_net), .O(n17265));   // verilog/coms.v(206[5:16])
    defparam i1_2_lut_3_lut_adj_1187.LUT_INIT = 16'hfdfd;
    SB_LUT4 i14_4_lut_adj_1188 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [22]), .I3(\FRAME_MATCHER.i [25]), .O(n39));
    defparam i14_4_lut_adj_1188.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1189 (.I0(\FRAME_MATCHER.state [2]), .I1(n17045), 
            .I2(\FRAME_MATCHER.state [1]), .I3(GND_net), .O(n17266));   // verilog/coms.v(206[5:16])
    defparam i1_2_lut_3_lut_adj_1189.LUT_INIT = 16'hfdfd;
    SB_LUT4 i13_3_lut (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [18]), 
            .I2(\FRAME_MATCHER.i [8]), .I3(GND_net), .O(n38));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i12_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(\FRAME_MATCHER.i [10]), 
            .I2(GND_net), .I3(GND_net), .O(n37));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i23_4_lut_adj_1190 (.I0(n39), .I1(n41), .I2(n40_adj_4114), 
            .I3(n42_adj_4113), .O(n48_adj_4115));
    defparam i23_4_lut_adj_1190.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1191 (.I0(\FRAME_MATCHER.i [19]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [9]), .I3(\FRAME_MATCHER.i [27]), .O(n43_adj_4116));
    defparam i18_4_lut_adj_1191.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut_adj_1192 (.I0(n43_adj_4116), .I1(n48_adj_4115), .I2(n37), 
            .I3(n38), .O(n17208));
    defparam i24_4_lut_adj_1192.LUT_INIT = 16'hfffe;
    SB_LUT4 i33761_4_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [2]), .I2(\data_in[0] [3]), 
            .I3(\data_in[1] [0]), .O(n40827));
    defparam i33761_4_lut.LUT_INIT = 16'h8000;
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(clk32MHz), 
           .D(n36597));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_32_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n30331), .O(n2_adj_4071)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_32_lut.LUT_INIT = 16'h8228;
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n18801));   // verilog/coms.v(126[12] 289[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n18800));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n18799));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n19199));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 n45980_bdd_4_lut (.I0(n45980), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(byte_transmit_counter[1]), 
            .O(n45983));
    defparam n45980_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1193 (.I0(\data_in[2] [4]), .I1(\data_in[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4117));
    defparam i1_2_lut_adj_1193.LUT_INIT = 16'heeee;
    SB_CARRY add_44_32 (.CI(n30331), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n30332));
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n19203));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 equal_107_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3947));   // verilog/coms.v(154[7:23])
    defparam equal_107_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_adj_1194 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[15] [7]), 
            .I2(n37839), .I3(GND_net), .O(n6_adj_3925));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1194.LUT_INIT = 16'h9696;
    SB_LUT4 add_44_31_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n30330), .O(n2_adj_4069)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_31_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n18798));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n18797));   // verilog/coms.v(126[12] 289[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n18796));   // verilog/coms.v(126[12] 289[6])
    SB_DFF gearBoxRatio_i0_i0 (.Q(gearBoxRatio[0]), .C(clk32MHz), .D(n18795));   // verilog/coms.v(126[12] 289[6])
    SB_DFF LED_3230 (.Q(LED_c), .C(clk32MHz), .D(n38165));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1195 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[15] [7]), 
            .I2(\data_out_frame[15] [5]), .I3(n17963), .O(n37687));   // verilog/coms.v(76[16:27])
    defparam i2_3_lut_4_lut_adj_1195.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1196 (.I0(n33854), .I1(n22_adj_4118), .I2(n11), 
            .I3(\data_in_frame[4] [7]), .O(n27_adj_4119));   // verilog/coms.v(230[9:81])
    defparam i11_4_lut_adj_1196.LUT_INIT = 16'hfdfe;
    SB_LUT4 i9_4_lut_adj_1197 (.I0(n33886), .I1(n17863), .I2(n17844), 
            .I3(n18119), .O(n25_adj_4120));   // verilog/coms.v(230[9:81])
    defparam i9_4_lut_adj_1197.LUT_INIT = 16'hfffe;
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n19175));   // verilog/coms.v(126[12] 289[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n19353));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_31 (.CI(n30330), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n30331));
    SB_LUT4 i7_4_lut_adj_1198 (.I0(n9_adj_4117), .I1(n40827), .I2(\data_in[3] [0]), 
            .I3(\data_in[0] [6]), .O(n17167));
    defparam i7_4_lut_adj_1198.LUT_INIT = 16'hffbf;
    SB_LUT4 i18_4_lut_adj_1199 (.I0(n31_adj_4110), .I1(n33), .I2(n32), 
            .I3(n34), .O(n37209));   // verilog/coms.v(206[5:16])
    defparam i18_4_lut_adj_1199.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut_adj_1200 (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4121));
    defparam i2_2_lut_adj_1200.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1201 (.I0(\data_in[0] [2]), .I1(\data_in[3] [5]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_4122));
    defparam i6_4_lut_adj_1201.LUT_INIT = 16'hfeff;
    SB_LUT4 i7_4_lut_adj_1202 (.I0(\data_in[3] [6]), .I1(n14_adj_4122), 
            .I2(n10_adj_4121), .I3(\data_in[2] [1]), .O(n17247));
    defparam i7_4_lut_adj_1202.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_4_lut_adj_1203 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_4123));
    defparam i4_4_lut_adj_1203.LUT_INIT = 16'hfdff;
    SB_LUT4 i5_3_lut_adj_1204 (.I0(\data_in[2] [7]), .I1(n10_adj_4123), 
            .I2(\data_in[3] [4]), .I3(GND_net), .O(n17222));
    defparam i5_3_lut_adj_1204.LUT_INIT = 16'hdfdf;
    SB_LUT4 i33744_2_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n40809));
    defparam i33744_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i8_4_lut_adj_1205 (.I0(n17222), .I1(\data_in[2] [6]), .I2(\data_in[3] [7]), 
            .I3(n17247), .O(n21_adj_4124));
    defparam i8_4_lut_adj_1205.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1206 (.I0(\data_in_frame[13] [4]), .I1(Kp_23__N_1433), 
            .I2(GND_net), .I3(GND_net), .O(n37398));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1206.LUT_INIT = 16'h6666;
    SB_LUT4 i7_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[0] [1]), .I2(\data_in[1] [6]), 
            .I3(GND_net), .O(n20_adj_4125));
    defparam i7_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i3_4_lut_adj_1207 (.I0(\FRAME_MATCHER.state [4]), .I1(\FRAME_MATCHER.state [7]), 
            .I2(\FRAME_MATCHER.state [6]), .I3(\FRAME_MATCHER.state [5]), 
            .O(n37378));
    defparam i3_4_lut_adj_1207.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_2_lut (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n37386));   // verilog/coms.v(94[12:25])
    defparam i24_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1208 (.I0(n37378), .I1(n37209), .I2(n33677), 
            .I3(GND_net), .O(n17045));   // verilog/coms.v(206[5:16])
    defparam i2_3_lut_adj_1208.LUT_INIT = 16'hfefe;
    SB_LUT4 add_44_30_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n30329), .O(n2_adj_4067)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_30 (.CI(n30329), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n30330));
    SB_LUT4 add_44_29_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n30328), .O(n2_adj_4065)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i11_4_lut_adj_1209 (.I0(n21_adj_4124), .I1(n17167), .I2(n40809), 
            .I3(\data_in[1] [3]), .O(n24_adj_4126));
    defparam i11_4_lut_adj_1209.LUT_INIT = 16'hefff;
    SB_LUT4 i12_4_lut_adj_1210 (.I0(\data_in[3] [2]), .I1(n24_adj_4126), 
            .I2(n20_adj_4125), .I3(\data_in[2] [0]), .O(n63));
    defparam i12_4_lut_adj_1210.LUT_INIT = 16'hfdff;
    SB_CARRY add_44_29 (.CI(n30328), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n30329));
    SB_LUT4 i2_3_lut_adj_1211 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n17199), .I3(GND_net), .O(n17200));   // verilog/coms.v(195[5:24])
    defparam i2_3_lut_adj_1211.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_3_lut_adj_1212 (.I0(\FRAME_MATCHER.state [2]), .I1(n63_c), 
            .I2(n63_adj_3909), .I3(GND_net), .O(n20639));   // verilog/coms.v(110[11:16])
    defparam i1_3_lut_adj_1212.LUT_INIT = 16'hb3b3;
    SB_LUT4 i1_2_lut_adj_1213 (.I0(n37489), .I1(n37710), .I2(GND_net), 
            .I3(GND_net), .O(n33828));
    defparam i1_2_lut_adj_1213.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(clk32MHz), 
           .D(n19258));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_28_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n30327), .O(n2_adj_4063)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_28 (.CI(n30327), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n30328));
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n19257));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n19256));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1214 (.I0(n37413), .I1(n10_adj_3931), .I2(\data_out_frame[6] [7]), 
            .I3(\data_out_frame[13] [3]), .O(n37578));
    defparam i1_2_lut_4_lut_adj_1214.LUT_INIT = 16'h6996;
    SB_LUT4 select_357_Select_2_i5_4_lut (.I0(n2857), .I1(n17268), .I2(n63), 
            .I3(n20639), .O(n5));
    defparam select_357_Select_2_i5_4_lut.LUT_INIT = 16'h3222;
    SB_LUT4 i1_rep_207_2_lut (.I0(n63), .I1(n20639), .I2(GND_net), .I3(GND_net), 
            .O(n46559));   // verilog/coms.v(110[11:16])
    defparam i1_rep_207_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_adj_1215 (.I0(n37413), .I1(n10_adj_3931), .I2(\data_out_frame[6] [7]), 
            .I3(n16787), .O(n37508));
    defparam i1_2_lut_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n19255));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n19254));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n19253));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n19252));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_27_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n30326), .O(n2_adj_4061)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_27 (.CI(n30326), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n30327));
    SB_LUT4 i1_3_lut_adj_1216 (.I0(\data_in_frame[5] [2]), .I1(\data_in_frame[3] [1]), 
            .I2(n37489), .I3(GND_net), .O(n17636));
    defparam i1_3_lut_adj_1216.LUT_INIT = 16'h9696;
    SB_LUT4 Kp_23__I_0_2_lut (.I0(n31_adj_4105), .I1(Kp_23__N_1745), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_718));   // verilog/coms.v(258[9] 260[65])
    defparam Kp_23__I_0_2_lut.LUT_INIT = 16'h4444;
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n19251));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_26_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n30325), .O(n2_adj_4059)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_26 (.CI(n30325), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n30326));
    SB_LUT4 i1_4_lut_4_lut_adj_1217 (.I0(n63), .I1(n740), .I2(n38092), 
            .I3(n17202), .O(n5_adj_3));   // verilog/coms.v(157[6] 159[9])
    defparam i1_4_lut_4_lut_adj_1217.LUT_INIT = 16'h0a2a;
    SB_LUT4 add_44_25_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n30324), .O(n2_adj_4057)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i21318_2_lut_3_lut (.I0(n63), .I1(n740), .I2(n93[1]), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_2460 [1]));   // verilog/coms.v(157[6] 159[9])
    defparam i21318_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n19250));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n19249));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n19248));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n19247));   // verilog/coms.v(126[12] 289[6])
    SB_CARRY add_44_25 (.CI(n30324), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n30325));
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n19246));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_24_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n30323), .O(n2_adj_4055)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i33794_3_lut_4_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[1]), 
            .I2(n40965), .I3(n40963), .O(n40918));
    defparam i33794_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_CARRY add_44_24 (.CI(n30323), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n30324));
    SB_LUT4 i33791_3_lut_4_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[1]), 
            .I2(n40956), .I3(n40954), .O(n40915));
    defparam i33791_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n19245));   // verilog/coms.v(126[12] 289[6])
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n18664));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n19239));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n19202));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 add_44_23_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n30322), .O(n2_adj_4053)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_23 (.CI(n30322), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n30323));
    SB_LUT4 i33788_3_lut_4_lut (.I0(byte_transmit_counter[2]), .I1(byte_transmit_counter[1]), 
            .I2(n40911), .I3(n40909), .O(n40912));
    defparam i33788_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 add_44_20_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n30319), .O(n2_adj_4047)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15_4_lut_adj_1218 (.I0(n25_adj_4120), .I1(n27_adj_4119), .I2(n26_adj_4111), 
            .I3(n28_adj_4099), .O(n31));   // verilog/coms.v(230[9:81])
    defparam i15_4_lut_adj_1218.LUT_INIT = 16'hfffe;
    SB_CARRY add_44_22 (.CI(n30321), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n30322));
    SB_LUT4 i15_2_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_4129));
    defparam i15_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_4_lut_adj_1219 (.I0(n37687), .I1(n10_adj_3923), .I2(n33049), 
            .I3(n37872), .O(n6_adj_3919));
    defparam i1_2_lut_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_LUT4 add_44_21_lut (.I0(n1972), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n30320), .O(n2_adj_4049)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_3_lut_adj_1220 (.I0(n33070), .I1(\data_in_frame[7] [1]), 
            .I2(\data_in_frame[9] [3]), .I3(GND_net), .O(n37854));
    defparam i2_3_lut_adj_1220.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1221 (.I0(\data_in_frame[6] [7]), .I1(n17900), 
            .I2(GND_net), .I3(GND_net), .O(n17853));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1221.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1222 (.I0(\data_in_frame[9] [4]), .I1(n17636), 
            .I2(n33828), .I3(\data_in_frame[5] [0]), .O(n37619));
    defparam i3_4_lut_adj_1222.LUT_INIT = 16'h9669;
    SB_CARRY add_44_21 (.CI(n30320), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n30321));
    SB_LUT4 i1_2_lut_4_lut_adj_1223 (.I0(n37687), .I1(n10_adj_3923), .I2(n33049), 
            .I3(n32717), .O(n33941));
    defparam i1_2_lut_4_lut_adj_1223.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1224 (.I0(\data_out_frame[15] [1]), .I1(n33822), 
            .I2(n33047), .I3(GND_net), .O(n37869));
    defparam i1_2_lut_3_lut_adj_1224.LUT_INIT = 16'h6969;
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n19201));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n19244));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n19243));   // verilog/coms.v(126[12] 289[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n19242));   // verilog/coms.v(126[12] 289[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1225 (.I0(\data_out_frame[15] [1]), .I1(n33822), 
            .I2(n33049), .I3(GND_net), .O(n37665));
    defparam i1_2_lut_3_lut_adj_1225.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1226 (.I0(\data_out_frame[19] [1]), .I1(n33008), 
            .I2(n32717), .I3(\data_out_frame[19] [2]), .O(n38922));
    defparam i2_3_lut_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1227 (.I0(n37640), .I1(n37863), .I2(n37801), 
            .I3(n37666), .O(n38857));
    defparam i2_3_lut_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1228 (.I0(n37640), .I1(n37863), .I2(n37666), 
            .I3(\data_out_frame[20] [1]), .O(n37826));
    defparam i1_2_lut_3_lut_4_lut_adj_1228.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1229 (.I0(n37640), .I1(n37863), .I2(n37549), 
            .I3(\data_out_frame[20] [1]), .O(n37825));
    defparam i1_2_lut_3_lut_4_lut_adj_1229.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1230 (.I0(n33882), .I1(n17671), .I2(n37482), 
            .I3(GND_net), .O(n6_adj_3915));
    defparam i1_2_lut_3_lut_adj_1230.LUT_INIT = 16'h6969;
    SB_LUT4 i15539_4_lut (.I0(\data_out_frame[0] [1]), .I1(n6119), .I2(n18435), 
            .I3(ID1), .O(n18910));
    defparam i15539_4_lut.LUT_INIT = 16'h3a0a;
    SB_LUT4 i11_3_lut_adj_1231 (.I0(byte_transmit_counter[1]), .I1(n42973), 
            .I2(n18381), .I3(GND_net), .O(n36213));   // verilog/coms.v(100[12:33])
    defparam i11_3_lut_adj_1231.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_3_lut_adj_1232 (.I0(byte_transmit_counter[2]), .I1(n42974), 
            .I2(n18381), .I3(GND_net), .O(n36219));   // verilog/coms.v(100[12:33])
    defparam i11_3_lut_adj_1232.LUT_INIT = 16'hcaca;
    SB_LUT4 i15448_3_lut (.I0(byte_transmit_counter[3]), .I1(n42881), .I2(n18381), 
            .I3(GND_net), .O(n18913));
    defparam i15448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15452_3_lut (.I0(byte_transmit_counter[4]), .I1(n42884), .I2(n18381), 
            .I3(GND_net), .O(n18914));
    defparam i15452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1233 (.I0(n33882), .I1(n17671), .I2(\data_out_frame[20] [4]), 
            .I3(GND_net), .O(n33079));
    defparam i1_2_lut_3_lut_adj_1233.LUT_INIT = 16'h6969;
    SB_LUT4 i305_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17199), .I3(n14748), .O(n326));   // verilog/coms.v(113[11:12])
    defparam i305_2_lut_3_lut_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1234 (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(\FRAME_MATCHER.state[0] ), .I2(n17266), .I3(n14721), .O(n200));   // verilog/coms.v(216[5:21])
    defparam i1_2_lut_3_lut_4_lut_adj_1234.LUT_INIT = 16'h0400;
    SB_LUT4 i31038_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n17045), 
            .I2(n17263), .I3(n3761), .O(n38098));
    defparam i31038_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1235 (.I0(\data_out_frame[11] [5]), .I1(n17979), 
            .I2(n37496), .I3(n37575), .O(n32950));
    defparam i1_2_lut_3_lut_4_lut_adj_1235.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1236 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[5] [5]), .I3(n17821), .O(n6_adj_3944));
    defparam i1_2_lut_3_lut_4_lut_adj_1236.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1237 (.I0(n93[1]), .I1(n63), .I2(n37376), 
            .I3(GND_net), .O(n36585));   // verilog/coms.v(143[4] 146[7])
    defparam i1_2_lut_3_lut_adj_1237.LUT_INIT = 16'hb0b0;
    SB_LUT4 i1_3_lut_4_lut (.I0(n63), .I1(n20661), .I2(n3761), .I3(n17264), 
            .O(n301));   // verilog/coms.v(143[7:84])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i1_2_lut_adj_1238 (.I0(\data_in_frame[11] [5]), .I1(\data_in_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4130));
    defparam i1_2_lut_adj_1238.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_38839 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(byte_transmit_counter[1]), .O(n45974));
    defparam byte_transmit_counter_0__bdd_4_lut_38839.LUT_INIT = 16'he4aa;
    SB_LUT4 n45974_bdd_4_lut (.I0(n45974), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(byte_transmit_counter[1]), 
            .O(n45977));
    defparam n45974_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_4_lut_adj_1239 (.I0(n37619), .I1(n17853), .I2(n37854), 
            .I3(n6_adj_4130), .O(n37986));
    defparam i4_4_lut_adj_1239.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1240 (.I0(\data_in_frame[7] [5]), .I1(n37887), 
            .I2(n37971), .I3(\data_in_frame[13] [7]), .O(n14_adj_4131));
    defparam i6_4_lut_adj_1240.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_38834 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(byte_transmit_counter[1]), .O(n45968));
    defparam byte_transmit_counter_0__bdd_4_lut_38834.LUT_INIT = 16'he4aa;
    SB_LUT4 n45968_bdd_4_lut (.I0(n45968), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(byte_transmit_counter[1]), 
            .O(n45971));
    defparam n45968_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut_adj_1241 (.I0(\data_in_frame[14] [1]), .I1(n14_adj_4131), 
            .I2(n10_adj_4132), .I3(n37986), .O(n37523));
    defparam i7_4_lut_adj_1241.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_38829 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(byte_transmit_counter[1]), .O(n45962));
    defparam byte_transmit_counter_0__bdd_4_lut_38829.LUT_INIT = 16'he4aa;
    SB_LUT4 n45962_bdd_4_lut (.I0(n45962), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(byte_transmit_counter[1]), 
            .O(n44437));
    defparam n45962_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_38824 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(byte_transmit_counter[1]), .O(n45956));
    defparam byte_transmit_counter_0__bdd_4_lut_38824.LUT_INIT = 16'he4aa;
    SB_LUT4 n45956_bdd_4_lut (.I0(n45956), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(byte_transmit_counter[1]), 
            .O(n40996));
    defparam n45956_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_38819 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(byte_transmit_counter[1]), .O(n45950));
    defparam byte_transmit_counter_0__bdd_4_lut_38819.LUT_INIT = 16'he4aa;
    SB_LUT4 n45950_bdd_4_lut (.I0(n45950), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(byte_transmit_counter[1]), 
            .O(n45953));
    defparam n45950_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut_adj_1242 (.I0(n37533), .I1(n33886), .I2(n17827), 
            .I3(n10_adj_4133), .O(n16_adj_4134));
    defparam i7_4_lut_adj_1242.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_38814 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(byte_transmit_counter[1]), .O(n45944));
    defparam byte_transmit_counter_0__bdd_4_lut_38814.LUT_INIT = 16'he4aa;
    SB_LUT4 n45944_bdd_4_lut (.I0(n45944), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(byte_transmit_counter[1]), 
            .O(n45947));
    defparam n45944_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1243 (.I0(n33864), .I1(n18295), .I2(n17853), 
            .I3(\data_in_frame[9] [3]), .O(n15_adj_4135));
    defparam i6_4_lut_adj_1243.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_38809 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(byte_transmit_counter[1]), .O(n45938));
    defparam byte_transmit_counter_0__bdd_4_lut_38809.LUT_INIT = 16'he4aa;
    SB_LUT4 n45938_bdd_4_lut (.I0(n45938), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(byte_transmit_counter[1]), 
            .O(n45941));
    defparam n45938_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_4_lut_adj_1244 (.I0(n15_adj_4135), .I1(n37523), .I2(n16_adj_4134), 
            .I3(\data_in_frame[14] [0]), .O(n33880));
    defparam i2_4_lut_adj_1244.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1245 (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[16] [2]), 
            .I2(n33880), .I3(n17874), .O(n37726));
    defparam i1_4_lut_adj_1245.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_2__bdd_4_lut (.I0(byte_transmit_counter[2]), 
            .I1(n40996), .I2(n44437), .I3(byte_transmit_counter[3]), .O(n45926));
    defparam byte_transmit_counter_2__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n45926_bdd_4_lut (.I0(n45926), .I1(n40946), .I2(n40945), .I3(byte_transmit_counter[3]), 
            .O(n45929));
    defparam n45926_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_in_frame[1] [2]), .I1(n37914), 
            .I2(n17636), .I3(\data_in_frame[10] [0]), .O(n10_adj_4000));
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9383_2_lut_4_lut (.I0(Kp_23__N_1745), .I1(n31_adj_4105), .I2(n31), 
            .I3(\FRAME_MATCHER.state [1]), .O(n12503));
    defparam i9383_2_lut_4_lut.LUT_INIT = 16'h0a22;
    SB_LUT4 i1_2_lut_3_lut_adj_1246 (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[0] [0]), 
            .I2(Kp_23__N_839), .I3(GND_net), .O(n33430));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_3_lut_adj_1246.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1247 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n3_adj_3997));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1247.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1248 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[1] [3]), 
            .I2(n37470), .I3(n6_adj_3977), .O(Kp_23__N_858));   // verilog/coms.v(71[16:34])
    defparam i4_4_lut_adj_1248.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1249 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(Kp_23__N_858), .I3(\data_in_frame[1] [0]), .O(n37526));   // verilog/coms.v(68[16:69])
    defparam i3_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1250 (.I0(\data_in_frame[5] [6]), .I1(\data_in_frame[4] [0]), 
            .I2(\data_in_frame[10] [3]), .I3(Kp_23__N_1083), .O(n12_adj_4136));   // verilog/coms.v(94[12:25])
    defparam i5_4_lut_adj_1250.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1251 (.I0(\data_in_frame[12] [4]), .I1(n12_adj_4136), 
            .I2(\data_in_frame[8] [2]), .I3(\data_in_frame[10] [2]), .O(n37747));   // verilog/coms.v(94[12:25])
    defparam i6_4_lut_adj_1251.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1252 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n37470));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_adj_1252.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1253 (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n37597));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_adj_1253.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1254 (.I0(n17636), .I1(\data_in_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n37908));
    defparam i1_2_lut_adj_1254.LUT_INIT = 16'h6666;
    SB_LUT4 i3_3_lut_adj_1255 (.I0(n5_adj_3989), .I1(n37908), .I2(\data_in_frame[10] [0]), 
            .I3(GND_net), .O(n37780));
    defparam i3_3_lut_adj_1255.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1256 (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[4] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4137));
    defparam i1_2_lut_adj_1256.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1257 (.I0(n37699), .I1(n18001), .I2(n37619), 
            .I3(n6_adj_4137), .O(n37989));
    defparam i4_4_lut_adj_1257.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1258 (.I0(\data_in_frame[7] [4]), .I1(n37989), 
            .I2(GND_net), .I3(GND_net), .O(n37714));
    defparam i1_2_lut_adj_1258.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1259 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[4] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n37875));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_1259.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1260 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[2] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n37655));   // verilog/coms.v(68[16:27])
    defparam i1_2_lut_adj_1260.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1261 (.I0(\data_in_frame[7] [3]), .I1(\data_in_frame[4] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n18001));
    defparam i1_2_lut_adj_1261.LUT_INIT = 16'h6666;
    SB_LUT4 i15626_4_lut_4_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state[0] ), 
            .O(n16726));   // verilog/coms.v(110[11:16])
    defparam i15626_4_lut_4_lut.LUT_INIT = 16'h2026;
    SB_LUT4 i1_2_lut_adj_1262 (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n37968));
    defparam i1_2_lut_adj_1262.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1263 (.I0(\data_in_frame[15] [4]), .I1(n17928), 
            .I2(GND_net), .I3(GND_net), .O(n37732));
    defparam i1_2_lut_adj_1263.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1264 (.I0(\data_in_frame[8] [4]), .I1(\data_in_frame[11] [0]), 
            .I2(\data_in_frame[8] [6]), .I3(\data_in_frame[8] [7]), .O(n10_adj_4138));   // verilog/coms.v(69[16:27])
    defparam i4_4_lut_adj_1264.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1265 (.I0(\data_in_frame[10] [6]), .I1(n10_adj_4138), 
            .I2(\data_in_frame[8] [5]), .I3(GND_net), .O(n37433));   // verilog/coms.v(69[16:27])
    defparam i5_3_lut_adj_1265.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1266 (.I0(\data_in_frame[13] [2]), .I1(n37776), 
            .I2(n37433), .I3(n17840), .O(n17542));   // verilog/coms.v(69[16:27])
    defparam i3_4_lut_adj_1266.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1267 (.I0(n39322), .I1(n33850), .I2(\data_in_frame[14] [3]), 
            .I3(GND_net), .O(n37628));
    defparam i2_3_lut_adj_1267.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1268 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n37616));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1268.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1269 (.I0(n17492), .I1(n17900), .I2(\data_in_frame[6] [6]), 
            .I3(GND_net), .O(n18295));
    defparam i2_3_lut_adj_1269.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1270 (.I0(n37769), .I1(n37896), .I2(\data_in_frame[13] [3]), 
            .I3(n17425), .O(n12_adj_4139));   // verilog/coms.v(69[16:27])
    defparam i5_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1271 (.I0(n18091), .I1(n12_adj_4139), .I2(n37932), 
            .I3(n17840), .O(n17928));   // verilog/coms.v(69[16:27])
    defparam i6_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1272 (.I0(n37410), .I1(n37760), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1562));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1272.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [1]), .I3(n38088), .O(n6121));
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h0054;
    SB_LUT4 i4_4_lut_adj_1273 (.I0(n37398), .I1(n37476), .I2(\data_in_frame[16] [0]), 
            .I3(Kp_23__N_1562), .O(n10_adj_4140));   // verilog/coms.v(73[16:43])
    defparam i4_4_lut_adj_1273.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1274 (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[15] [5]), 
            .I2(n10_adj_4140), .I3(n17928), .O(n37953));
    defparam i1_4_lut_adj_1274.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1275 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[8] [3]), 
            .I2(\data_in_frame[6] [2]), .I3(GND_net), .O(n37959));   // verilog/coms.v(70[16:41])
    defparam i2_3_lut_adj_1275.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1276 (.I0(\data_in_frame[10] [5]), .I1(n37959), 
            .I2(n8_adj_4096), .I3(\data_in_frame[8] [4]), .O(n37789));   // verilog/coms.v(72[16:43])
    defparam i3_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1277 (.I0(n37789), .I1(n37932), .I2(\data_in_frame[10] [7]), 
            .I3(n37392), .O(n12_adj_4141));   // verilog/coms.v(72[16:43])
    defparam i5_4_lut_adj_1277.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1278 (.I0(\data_in_frame[11] [7]), .I1(\data_in_frame[9] [5]), 
            .I2(\data_in_frame[9] [6]), .I3(\data_in_frame[12] [0]), .O(n37887));
    defparam i1_2_lut_3_lut_4_lut_adj_1278.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1279 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [2]), .I3(n6_adj_4020), .O(Kp_23__N_893));   // verilog/coms.v(94[12:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1280 (.I0(\data_in_frame[12] [7]), .I1(n12_adj_4141), 
            .I2(n37980), .I3(n17404), .O(n18140));   // verilog/coms.v(72[16:43])
    defparam i6_4_lut_adj_1280.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1281 (.I0(n18023), .I1(\data_in_frame[18] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n32943));
    defparam i1_2_lut_adj_1281.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1282 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[0] [2]), .I3(n4_adj_4142), .O(n37698));   // verilog/coms.v(94[12:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1282.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[4] [6]), 
            .I2(n10_adj_4143), .I3(\data_in_frame[8] [7]), .O(n18023));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1283 (.I0(\data_in_frame[15] [3]), .I1(n18228), 
            .I2(n18140), .I3(n6_adj_4144), .O(n37738));
    defparam i4_4_lut_adj_1283.LUT_INIT = 16'h6996;
    SB_LUT4 data_in_frame_4__7__I_0_3240_2_lut (.I0(\data_in_frame[4] [7]), 
            .I1(\data_in_frame[4] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_820));   // verilog/coms.v(69[16:27])
    defparam data_in_frame_4__7__I_0_3240_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1284 (.I0(\data_in_frame[8] [5]), .I1(n17492), 
            .I2(\data_in_frame[6] [5]), .I3(GND_net), .O(n37932));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_3_lut_adj_1284.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1285 (.I0(n17492), .I1(n17900), .I2(\data_in_frame[6] [6]), 
            .I3(n37616), .O(n17840));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_4_lut_adj_1285.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1286 (.I0(\data_in_frame[16] [5]), .I1(\data_in_frame[16] [4]), 
            .I2(\data_in_frame[16] [3]), .I3(GND_net), .O(n37410));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_adj_1286.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1287 (.I0(n17492), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n37450));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_1287.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1288 (.I0(n37410), .I1(n37760), .I2(n16859), 
            .I3(n32982), .O(n37857));
    defparam i2_3_lut_4_lut_adj_1288.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1289 (.I0(\data_in_frame[7] [2]), .I1(n37698), 
            .I2(GND_net), .I3(GND_net), .O(n37699));
    defparam i1_2_lut_adj_1289.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1290 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[14] [6]), 
            .I2(\data_in_frame[15] [0]), .I3(GND_net), .O(n37947));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_1290.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1291 (.I0(n63), .I1(n63_c), .I2(n63_adj_3909), 
            .I3(\FRAME_MATCHER.state[0] ), .O(n40));   // verilog/coms.v(143[7:84])
    defparam i1_2_lut_3_lut_4_lut_adj_1291.LUT_INIT = 16'hff7f;
    SB_LUT4 i4_4_lut_adj_1292 (.I0(\data_in_frame[9] [1]), .I1(n37450), 
            .I2(\data_in_frame[11] [3]), .I3(\data_in_frame[11] [4]), .O(n10_adj_4146));   // verilog/coms.v(83[17:70])
    defparam i4_4_lut_adj_1292.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1293 (.I0(\data_in_frame[7] [0]), .I1(n10_adj_4146), 
            .I2(n17863), .I3(GND_net), .O(n37693));   // verilog/coms.v(83[17:70])
    defparam i5_3_lut_adj_1293.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1294 (.I0(n37693), .I1(n37699), .I2(n11), .I3(n37854), 
            .O(n10_adj_4143));
    defparam i4_4_lut_adj_1294.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1295 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[7] [2]), 
            .I2(n37698), .I3(GND_net), .O(n37533));
    defparam i1_2_lut_3_lut_adj_1295.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1296 (.I0(\data_in_frame[1] [2]), .I1(n37914), 
            .I2(n17636), .I3(GND_net), .O(n37971));
    defparam i1_2_lut_3_lut_adj_1296.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1297 (.I0(\data_in_frame[14] [0]), .I1(n37986), 
            .I2(\data_in_frame[13] [5]), .I3(\data_in_frame[15] [7]), .O(n37443));   // verilog/coms.v(72[16:43])
    defparam i3_4_lut_adj_1297.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1298 (.I0(\data_in_frame[13] [7]), .I1(n37443), 
            .I2(n33843), .I3(n18023), .O(n16859));   // verilog/coms.v(72[16:43])
    defparam i3_4_lut_adj_1298.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1299 (.I0(\data_in_frame[18] [3]), .I1(n16859), 
            .I2(GND_net), .I3(GND_net), .O(n33035));
    defparam i1_2_lut_adj_1299.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i16_3_lut (.I0(\data_out_frame[16] [6]), 
            .I1(\data_out_frame[17] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4147));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1300 (.I0(n17687), .I1(\data_in_frame[7] [3]), 
            .I2(\data_in_frame[4] [7]), .I3(GND_net), .O(n37902));
    defparam i1_2_lut_3_lut_adj_1300.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[3] [4]), 
            .I2(\data_in_frame[3] [5]), .I3(n37567), .O(n17449));   // verilog/coms.v(83[17:28])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i17_3_lut (.I0(\data_out_frame[18] [6]), 
            .I1(\data_out_frame[19] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4148));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35976_2_lut (.I0(\data_out_frame[22] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n42810));
    defparam i35976_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i19_3_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\data_out_frame[21] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_4149));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i16_3_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\data_out_frame[17] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4150));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1301 (.I0(n326), .I1(n200), .I2(n324), 
            .I3(\FRAME_MATCHER.state [30]), .O(n8_adj_4089));
    defparam i1_2_lut_4_lut_adj_1301.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1302 (.I0(n63), .I1(n63_c), .I2(n63_adj_3909), 
            .I3(n2857), .O(n14721));   // verilog/coms.v(143[7:84])
    defparam i1_2_lut_3_lut_4_lut_adj_1302.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_4_lut_adj_1303 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(n33843), .I3(\data_in_frame[11] [4]), .O(n10_adj_4133));
    defparam i1_2_lut_4_lut_adj_1303.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i17_3_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\data_out_frame[19] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4151));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1304 (.I0(\data_in_frame[16] [4]), .I1(n39322), 
            .I2(n33850), .I3(\data_in_frame[14] [3]), .O(n17874));
    defparam i1_2_lut_4_lut_adj_1304.LUT_INIT = 16'h9669;
    SB_LUT4 i36236_2_lut (.I0(\data_out_frame[22] [5]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n42811));
    defparam i36236_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i19_3_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\data_out_frame[21] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_4152));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut_adj_1305 (.I0(n37878), .I1(n37776), .I2(\data_in_frame[12] [6]), 
            .I3(\data_in_frame[17] [1]), .O(n18_adj_4153));   // verilog/coms.v(74[16:43])
    defparam i7_4_lut_adj_1305.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i16_3_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\data_out_frame[17] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4154));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i17_3_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\data_out_frame[19] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4155));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36215_2_lut (.I0(\data_out_frame[22] [4]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n42818));
    defparam i36215_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i19_3_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\data_out_frame[21] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_4156));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31104_3_lut_4_lut (.I0(n63), .I1(n20661), .I2(LED_c), .I3(n17201), 
            .O(n38165));   // verilog/coms.v(143[7:84])
    defparam i31104_3_lut_4_lut.LUT_INIT = 16'hf700;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i16_3_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\data_out_frame[17] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4157));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i17_3_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\data_out_frame[19] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4158));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36510_2_lut (.I0(\data_out_frame[22] [7]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n42987));
    defparam i36510_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i19_3_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\data_out_frame[21] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_4159));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i16_3_lut (.I0(\data_out_frame[16] [3]), 
            .I1(\data_out_frame[17] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n16_adj_4160));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i17_3_lut (.I0(\data_out_frame[18] [3]), 
            .I1(\data_out_frame[19] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n17_adj_4161));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36229_2_lut (.I0(\data_out_frame[22] [3]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n42819));
    defparam i36229_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i19_3_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\data_out_frame[21] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_4162));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i301_3_lut_4_lut (.I0(n63), .I1(n20661), .I2(n26317), .I3(n17265), 
            .O(n322));   // verilog/coms.v(143[7:84])
    defparam i301_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i33821_3_lut (.I0(\data_out_frame[0][4] ), .I1(byte_transmit_counter[0]), 
            .I2(byte_transmit_counter[1]), .I3(GND_net), .O(n40945));
    defparam i33821_3_lut.LUT_INIT = 16'hc2c2;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4163));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33822_4_lut (.I0(\data_out_frame[5] [4]), .I1(n5_adj_4163), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n40946));
    defparam i33822_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i6_3_lut_4_lut (.I0(\data_in_frame[2] [4]), .I1(n37383), .I2(\data_in_frame[0] [7]), 
            .I3(\data_in_frame[1] [1]), .O(n22_adj_4164));   // verilog/coms.v(94[12:25])
    defparam i6_3_lut_4_lut.LUT_INIT = 16'h9009;
    SB_LUT4 i2_2_lut_4_lut_adj_1306 (.I0(n33070), .I1(n33854), .I2(n17687), 
            .I3(n18001), .O(n10_adj_4132));
    defparam i2_2_lut_4_lut_adj_1306.LUT_INIT = 16'h6996;
    SB_LUT4 i303_2_lut_3_lut_4_lut (.I0(n63), .I1(n63_c), .I2(n63_adj_3909), 
            .I3(n2664), .O(n324));   // verilog/coms.v(143[7:84])
    defparam i303_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i2008_3_lut (.I0(n31_adj_4105), .I1(n31), .I2(\FRAME_MATCHER.state [1]), 
            .I3(GND_net), .O(n14340));
    defparam i2008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1307 (.I0(\data_in_frame[2] [4]), .I1(n37383), 
            .I2(\data_in_frame[4] [5]), .I3(n4_adj_3980), .O(n17900));   // verilog/coms.v(94[12:25])
    defparam i2_3_lut_4_lut_adj_1307.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1308 (.I0(n39322), .I1(n37523), .I2(n37628), 
            .I3(n33295), .O(n32982));
    defparam i2_3_lut_4_lut_adj_1308.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1309 (.I0(n39322), .I1(n37523), .I2(\data_in_frame[16] [3]), 
            .I3(\data_in_frame[18] [4]), .O(n37517));
    defparam i2_3_lut_4_lut_adj_1309.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1310 (.I0(\data_in_frame[11] [7]), .I1(n37905), 
            .I2(\data_in_frame[7] [7]), .I3(n10_adj_3991), .O(n33850));
    defparam i5_3_lut_4_lut_adj_1310.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1311 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [31]), 
            .I3(GND_net), .O(n7_adj_4090));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1311.LUT_INIT = 16'he0e0;
    SB_LUT4 i5_2_lut_4_lut (.I0(n37476), .I1(\data_in_frame[16] [6]), .I2(n33087), 
            .I3(n17844), .O(n16_adj_4165));
    defparam i5_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1312 (.I0(n37476), .I1(\data_in_frame[16] [6]), 
            .I2(n33087), .I3(\data_in_frame[19] [0]), .O(n18122));
    defparam i1_2_lut_4_lut_adj_1312.LUT_INIT = 16'h6996;
    SB_LUT4 i14143_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37361), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n19175));
    defparam i14143_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14144_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37361), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n19176));
    defparam i14144_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14137_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37361), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n19169));
    defparam i14137_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14138_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37361), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n19170));
    defparam i14138_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14139_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37361), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n19171));
    defparam i14139_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14140_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37361), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n19172));
    defparam i14140_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14141_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37361), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n19173));
    defparam i14141_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14142_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37361), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n19174));
    defparam i14142_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1313 (.I0(n63), .I1(n63_c), .I2(n63_adj_3909), 
            .I3(n740), .O(n14748));   // verilog/coms.v(143[7:84])
    defparam i1_2_lut_3_lut_4_lut_adj_1313.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1314 (.I0(\data_out_frame[20] [3]), .I1(n17671), 
            .I2(n37604), .I3(n37549), .O(n37551));
    defparam i1_2_lut_3_lut_4_lut_adj_1314.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1315 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [30]), 
            .I3(GND_net), .O(n36779));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1315.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1316 (.I0(\data_out_frame[20] [3]), .I1(n17671), 
            .I2(n37604), .I3(n33079), .O(n17597));
    defparam i1_2_lut_3_lut_4_lut_adj_1316.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1317 (.I0(n37640), .I1(n18200), .I2(n33875), 
            .I3(n37801), .O(n37802));
    defparam i1_2_lut_3_lut_4_lut_adj_1317.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1318 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n26281), .O(n37361));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1318.LUT_INIT = 16'hfeff;
    SB_LUT4 i2_3_lut_4_lut_adj_1319 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n26281), .O(n37342));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1319.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_3_lut_adj_1320 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [29]), 
            .I3(GND_net), .O(n7_adj_4087));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1320.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1321 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n17263));   // verilog/coms.v(206[5:16])
    defparam i1_2_lut_3_lut_adj_1321.LUT_INIT = 16'hbfbf;
    SB_LUT4 mux_1033_i8_3_lut (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n4658), .I3(GND_net), .O(n4666));
    defparam mux_1033_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1322 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n17170));   // verilog/coms.v(206[5:16])
    defparam i1_2_lut_3_lut_adj_1322.LUT_INIT = 16'hfbfb;
    SB_LUT4 equal_108_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4166));   // verilog/coms.v(154[7:23])
    defparam equal_108_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 equal_109_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // verilog/coms.v(154[7:23])
    defparam equal_109_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i14263_3_lut_4_lut (.I0(n8), .I1(n37354), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n19295));
    defparam i14263_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14264_3_lut_4_lut (.I0(n8), .I1(n37354), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n19296));
    defparam i14264_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14257_3_lut_4_lut (.I0(n8), .I1(n37354), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n19289));
    defparam i14257_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1033_i7_3_lut (.I0(\data_in_frame[16] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n4658), .I3(GND_net), .O(n4665));
    defparam mux_1033_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14258_3_lut_4_lut (.I0(n8), .I1(n37354), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n19290));
    defparam i14258_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1323 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [28]), 
            .I3(GND_net), .O(n36775));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1323.LUT_INIT = 16'he0e0;
    SB_LUT4 i14259_3_lut_4_lut (.I0(n8), .I1(n37354), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n19291));
    defparam i14259_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14260_3_lut_4_lut (.I0(n8), .I1(n37354), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n19292));
    defparam i14260_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14261_3_lut_4_lut (.I0(n8), .I1(n37354), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n19293));
    defparam i14261_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1324 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [27]), 
            .I3(GND_net), .O(n7_adj_4085));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1324.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n19_adj_4162), .I2(n42819), .I3(byte_transmit_counter[2]), 
            .O(n45920));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 mux_1033_i18_3_lut (.I0(\data_in_frame[14] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n4658), .I3(GND_net), .O(n4676));
    defparam mux_1033_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14262_3_lut_4_lut (.I0(n8), .I1(n37354), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n19294));
    defparam i14262_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1325 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n17208), .I3(\FRAME_MATCHER.i [4]), .O(n17031));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1325.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1326 (.I0(\FRAME_MATCHER.i [3]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [4]), .I3(n26281), .O(n37354));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1326.LUT_INIT = 16'hefff;
    SB_LUT4 i14249_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37354), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n19281));
    defparam i14249_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14250_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37354), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n19282));
    defparam i14250_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14251_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37354), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n19283));
    defparam i14251_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14252_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37354), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n19284));
    defparam i14252_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14253_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37354), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n19285));
    defparam i14253_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14254_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37354), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n19286));
    defparam i14254_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14255_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37354), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n19287));
    defparam i14255_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14256_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37354), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n19288));
    defparam i14256_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_95_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_3907));   // verilog/coms.v(154[7:23])
    defparam equal_95_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 equal_94_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4167));   // verilog/coms.v(154[7:23])
    defparam equal_94_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 mux_1033_i17_3_lut (.I0(\data_in_frame[14] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n4658), .I3(GND_net), .O(n4675));
    defparam mux_1033_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1033_i16_3_lut (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n4658), .I3(GND_net), .O(n4674));
    defparam mux_1033_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1327 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [26]), 
            .I3(GND_net), .O(n36771));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1327.LUT_INIT = 16'he0e0;
    SB_LUT4 mux_1033_i20_3_lut (.I0(\data_in_frame[14] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n4658), .I3(GND_net), .O(n4678));
    defparam mux_1033_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1328 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [25]), 
            .I3(GND_net), .O(n36767));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1328.LUT_INIT = 16'he0e0;
    SB_LUT4 mux_1033_i19_3_lut (.I0(\data_in_frame[14] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n4658), .I3(GND_net), .O(n4677));
    defparam mux_1033_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1329 (.I0(\data_out_frame[19] [1]), .I1(\data_out_frame[18] [7]), 
            .I2(n37658), .I3(\data_out_frame[19] [0]), .O(n4_c));
    defparam i1_2_lut_3_lut_4_lut_adj_1329.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1330 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [24]), 
            .I3(GND_net), .O(n7_adj_4084));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1330.LUT_INIT = 16'he0e0;
    SB_LUT4 mux_1033_i22_3_lut (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n4658), .I3(GND_net), .O(n4680));
    defparam mux_1033_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1331 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [23]), 
            .I3(GND_net), .O(n7_adj_4082));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1331.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_adj_1332 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[3] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n37860));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_adj_1332.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1333 (.I0(n17559), .I1(n18_adj_4153), .I2(\data_in_frame[19] [2]), 
            .I3(\data_in_frame[6] [3]), .O(n20_adj_4168));   // verilog/coms.v(74[16:43])
    defparam i9_4_lut_adj_1333.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1334 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[15] [4]), 
            .I2(\data_in_frame[15] [3]), .I3(\data_in_frame[15] [2]), .O(n37974));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1334.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1335 (.I0(\data_in_frame[15] [5]), .I1(\data_in_frame[15] [4]), 
            .I2(n18023), .I3(\data_in_frame[18] [0]), .O(n6_adj_4144));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1335.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1336 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17266), .I3(GND_net), .O(n17268));   // verilog/coms.v(216[5:21])
    defparam i1_2_lut_3_lut_adj_1336.LUT_INIT = 16'hfbfb;
    SB_LUT4 i1_2_lut_3_lut_adj_1337 (.I0(\data_in_frame[1] [0]), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[0] [6]), .I3(GND_net), .O(n37750));   // verilog/coms.v(69[16:69])
    defparam i1_2_lut_3_lut_adj_1337.LUT_INIT = 16'h9696;
    SB_LUT4 i33738_2_lut_3_lut_4_lut (.I0(\data_in_frame[2] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(n4_adj_3980), .O(n40802));   // verilog/coms.v(74[16:27])
    defparam i33738_2_lut_3_lut_4_lut.LUT_INIT = 16'hff96;
    SB_LUT4 i1_2_lut_3_lut_adj_1338 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [22]), 
            .I3(GND_net), .O(n36763));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1338.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1339 (.I0(\data_in_frame[3] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n37386), .I3(n37710), .O(n4_adj_4142));   // verilog/coms.v(69[16:69])
    defparam i1_2_lut_3_lut_4_lut_adj_1339.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1340 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [21]), 
            .I3(GND_net), .O(n36807));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1340.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1341 (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n17199), .I3(GND_net), .O(n17202));   // verilog/coms.v(152[5:27])
    defparam i1_2_lut_3_lut_adj_1341.LUT_INIT = 16'hfbfb;
    SB_LUT4 mux_1033_i21_3_lut (.I0(\data_in_frame[14] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n4658), .I3(GND_net), .O(n4679));
    defparam mux_1033_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1342 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [20]), 
            .I3(GND_net), .O(n7_adj_4081));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1342.LUT_INIT = 16'he0e0;
    SB_LUT4 i14265_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37354), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n19297));
    defparam i14265_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1033_i24_3_lut (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n4658), .I3(GND_net), .O(n4682));
    defparam mux_1033_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14266_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37354), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n19298));
    defparam i14266_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1033_i23_3_lut (.I0(\data_in_frame[14] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n4658), .I3(GND_net), .O(n4681));
    defparam mux_1033_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i14267_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37354), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n19299));
    defparam i14267_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14268_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37354), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n19300));
    defparam i14268_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14269_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37354), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n19301));
    defparam i14269_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14270_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37354), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n19302));
    defparam i14270_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14271_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37354), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n19303));
    defparam i14271_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14272_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37354), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n19304));
    defparam i14272_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i22430_3_lut_4_lut (.I0(byte_transmit_counter[1]), .I1(byte_transmit_counter[2]), 
            .I2(byte_transmit_counter[4]), .I3(byte_transmit_counter[3]), 
            .O(n27441));
    defparam i22430_3_lut_4_lut.LUT_INIT = 16'hf080;
    SB_LUT4 n45920_bdd_4_lut (.I0(n45920), .I1(n17_adj_4161), .I2(n16_adj_4160), 
            .I3(byte_transmit_counter[2]), .O(n45923));
    defparam n45920_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1343 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [19]), 
            .I3(GND_net), .O(n36751));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1343.LUT_INIT = 16'he0e0;
    SB_LUT4 i10_4_lut_adj_1344 (.I0(n37947), .I1(n20_adj_4168), .I2(n16_adj_4165), 
            .I3(n37789), .O(n37820));   // verilog/coms.v(74[16:43])
    defparam i10_4_lut_adj_1344.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1345 (.I0(n37209), .I1(n37378), .I2(n33677), 
            .I3(GND_net), .O(n27475));   // verilog/coms.v(126[12] 289[6])
    defparam i2_3_lut_adj_1345.LUT_INIT = 16'hfefe;
    SB_LUT4 i15450_3_lut (.I0(byte_transmit_counter[5]), .I1(n42882), .I2(n18381), 
            .I3(GND_net), .O(n20482));
    defparam i15450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1346 (.I0(Kp_23__N_1745), .I1(n27475), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4169));
    defparam i1_2_lut_adj_1346.LUT_INIT = 16'hdddd;
    SB_LUT4 i5532_2_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10308));
    defparam i5532_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1347 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [18]), 
            .I3(GND_net), .O(n7_adj_4079));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1347.LUT_INIT = 16'he0e0;
    SB_LUT4 i15612_4_lut (.I0(Kp_23__N_718), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(\FRAME_MATCHER.state [1]), .I3(\FRAME_MATCHER.state [2]), 
            .O(n20642));   // verilog/coms.v(110[11:16])
    defparam i15612_4_lut.LUT_INIT = 16'hcacf;
    SB_LUT4 i1_2_lut_3_lut_adj_1348 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [17]), 
            .I3(GND_net), .O(n7_adj_4077));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1348.LUT_INIT = 16'he0e0;
    SB_LUT4 i4_4_lut_adj_1349 (.I0(\FRAME_MATCHER.state[0] ), .I1(n14340), 
            .I2(n47_adj_4129), .I3(n6_adj_4169), .O(n39863));
    defparam i4_4_lut_adj_1349.LUT_INIT = 16'hffef;
    SB_LUT4 i2_4_lut_adj_1350 (.I0(n16726), .I1(n27475), .I2(n20642), 
            .I3(n4658), .O(n18381));
    defparam i2_4_lut_adj_1350.LUT_INIT = 16'h2220;
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_in_frame[13] [4]), .I1(Kp_23__N_1433), 
            .I2(n37974), .I3(GND_net), .O(n8_adj_4101));   // verilog/coms.v(69[16:27])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i15454_3_lut (.I0(byte_transmit_counter[7]), .I1(n42885), .I2(n18381), 
            .I3(GND_net), .O(n19325));
    defparam i15454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31028_2_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(n27475), .I2(GND_net), 
            .I3(GND_net), .O(n38088));
    defparam i31028_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mux_1033_i9_3_lut (.I0(\data_in_frame[15] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n4658), .I3(GND_net), .O(n4667));
    defparam mux_1033_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1351 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n37607));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1351.LUT_INIT = 16'h6666;
    SB_LUT4 i33750_3_lut (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [0]), 
            .I2(ID0), .I3(GND_net), .O(n40815));
    defparam i33750_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 i33748_3_lut (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [2]), 
            .I2(ID2), .I3(GND_net), .O(n40813));
    defparam i33748_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 i5_4_lut_adj_1352 (.I0(\data_in_frame[0] [1]), .I1(n40815), 
            .I2(\data_in_frame[0] [7]), .I3(ID1), .O(n13));
    defparam i5_4_lut_adj_1352.LUT_INIT = 16'h0201;
    SB_LUT4 i7_4_lut_adj_1353 (.I0(n13), .I1(n40813), .I2(\data_in_frame[0] [6]), 
            .I3(\data_in_frame[0] [3]), .O(Kp_23__N_1746));
    defparam i7_4_lut_adj_1353.LUT_INIT = 16'h0002;
    SB_LUT4 i6_2_lut_3_lut (.I0(\data_in_frame[3] [5]), .I1(n37564), .I2(n17492), 
            .I3(GND_net), .O(n22_adj_4118));   // verilog/coms.v(230[9:81])
    defparam i6_2_lut_3_lut.LUT_INIT = 16'hf6f6;
    SB_LUT4 i3_4_lut_adj_1354 (.I0(\data_in_frame[0] [1]), .I1(n37607), 
            .I2(n37386), .I3(n37383), .O(Kp_23__N_839));   // verilog/coms.v(94[12:25])
    defparam i3_4_lut_adj_1354.LUT_INIT = 16'h6996;
    SB_LUT4 select_327_Select_31_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [31]), .I3(GND_net), .O(n3_adj_4074));
    defparam select_327_Select_31_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_38791 (.I0(byte_transmit_counter[1]), 
            .I1(n19_adj_4159), .I2(n42987), .I3(byte_transmit_counter[2]), 
            .O(n45914));
    defparam byte_transmit_counter_1__bdd_4_lut_38791.LUT_INIT = 16'he4aa;
    SB_LUT4 select_327_Select_30_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [30]), .I3(GND_net), .O(n3_adj_4072));
    defparam select_327_Select_30_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_1355 (.I0(\data_in_frame[0] [0]), .I1(Kp_23__N_839), 
            .I2(GND_net), .I3(GND_net), .O(n37514));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_adj_1355.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1356 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n39564));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_1356.LUT_INIT = 16'h9696;
    SB_LUT4 select_327_Select_29_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [29]), .I3(GND_net), .O(n3_adj_4070));
    defparam select_327_Select_29_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_327_Select_28_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [28]), .I3(GND_net), .O(n3_adj_4068));
    defparam select_327_Select_28_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_327_Select_27_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [27]), .I3(GND_net), .O(n3_adj_4066));
    defparam select_327_Select_27_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i10_4_lut_adj_1357 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[1] [3]), .I3(n39564), .O(n26_adj_4170));
    defparam i10_4_lut_adj_1357.LUT_INIT = 16'h0080;
    SB_LUT4 i1_2_lut_3_lut_adj_1358 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [16]), 
            .I3(GND_net), .O(n36831));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1358.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_3_lut_adj_1359 (.I0(Kp_23__N_839), .I1(Kp_23__N_1746), .I2(\data_in_frame[2] [1]), 
            .I3(GND_net), .O(n17_adj_4171));
    defparam i1_3_lut_adj_1359.LUT_INIT = 16'h4848;
    SB_LUT4 i12_4_lut_adj_1360 (.I0(n12_adj_3918), .I1(n3_adj_3997), .I2(n33430), 
            .I3(n6_adj_4020), .O(n28_adj_4172));
    defparam i12_4_lut_adj_1360.LUT_INIT = 16'h0020;
    SB_LUT4 select_327_Select_26_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [26]), .I3(GND_net), .O(n3_adj_4064));
    defparam select_327_Select_26_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i13_4_lut_adj_1361 (.I0(n17_adj_4171), .I1(n26_adj_4170), .I2(\data_in_frame[1] [6]), 
            .I3(\data_in_frame[1] [5]), .O(n29_adj_4173));
    defparam i13_4_lut_adj_1361.LUT_INIT = 16'h8000;
    SB_LUT4 i15_4_lut_adj_1362 (.I0(n29_adj_4173), .I1(n40802), .I2(n28_adj_4172), 
            .I3(n22_adj_4164), .O(\FRAME_MATCHER.state_31__N_2492 [3]));
    defparam i15_4_lut_adj_1362.LUT_INIT = 16'h2000;
    SB_LUT4 i2_4_lut_adj_1363 (.I0(\FRAME_MATCHER.state[3] ), .I1(n38088), 
            .I2(\FRAME_MATCHER.state [2]), .I3(\FRAME_MATCHER.state [1]), 
            .O(n6119));
    defparam i2_4_lut_adj_1363.LUT_INIT = 16'h0102;
    SB_LUT4 i2_3_lut_4_lut_adj_1364 (.I0(n33850), .I1(\data_in_frame[14] [4]), 
            .I2(\data_in_frame[14] [3]), .I3(n33852), .O(n33295));
    defparam i2_3_lut_4_lut_adj_1364.LUT_INIT = 16'h6996;
    SB_LUT4 select_327_Select_25_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [25]), .I3(GND_net), .O(n3_adj_4062));
    defparam select_327_Select_25_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1365 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [15]), 
            .I3(GND_net), .O(n7_adj_4075));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1365.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_4_lut_adj_1366 (.I0(n12503), .I1(n6121), .I2(n6119), .I3(\FRAME_MATCHER.state_31__N_2492 [3]), 
            .O(n18435));
    defparam i2_4_lut_adj_1366.LUT_INIT = 16'hc808;
    SB_LUT4 i1_2_lut_3_lut_adj_1367 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [14]), 
            .I3(GND_net), .O(n36827));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1367.LUT_INIT = 16'he0e0;
    SB_LUT4 select_327_Select_24_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [24]), .I3(GND_net), .O(n3_adj_4060));
    defparam select_327_Select_24_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_327_Select_23_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [23]), .I3(GND_net), .O(n3_adj_4058));
    defparam select_327_Select_23_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_327_Select_22_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [22]), .I3(GND_net), .O(n3_adj_4056));
    defparam select_327_Select_22_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1368 (.I0(\data_in_frame[6] [2]), .I1(n18119), 
            .I2(\data_in_frame[8] [4]), .I3(GND_net), .O(n37845));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_1368.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1369 (.I0(n17425), .I1(\data_in_frame[6] [2]), 
            .I2(n18119), .I3(GND_net), .O(n37776));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_3_lut_adj_1369.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1370 (.I0(\data_in_frame[13] [4]), .I1(\data_in_frame[13] [5]), 
            .I2(\data_in_frame[15] [6]), .I3(GND_net), .O(n17379));   // verilog/coms.v(72[16:43])
    defparam i1_2_lut_3_lut_adj_1370.LUT_INIT = 16'h9696;
    SB_LUT4 select_327_Select_21_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [21]), .I3(GND_net), .O(n3_adj_4054));
    defparam select_327_Select_21_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_327_Select_20_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [20]), .I3(GND_net), .O(n3_adj_4052));
    defparam select_327_Select_20_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1371 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[13] [6]), 
            .I2(n33843), .I3(GND_net), .O(n37622));
    defparam i1_2_lut_3_lut_adj_1371.LUT_INIT = 16'h9696;
    SB_LUT4 select_327_Select_19_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [19]), .I3(GND_net), .O(n3_adj_4050));
    defparam select_327_Select_19_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_327_Select_18_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [18]), .I3(GND_net), .O(n3_adj_4048));
    defparam select_327_Select_18_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1372 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [13]), 
            .I3(GND_net), .O(n36823));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1372.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_2_lut_4_lut_adj_1373 (.I0(n6_adj_4020), .I1(\data_in_frame[3] [0]), 
            .I2(n37750), .I3(n37710), .O(n33854));
    defparam i2_2_lut_4_lut_adj_1373.LUT_INIT = 16'h6996;
    SB_LUT4 select_327_Select_17_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [17]), .I3(GND_net), .O(n3_adj_4046));
    defparam select_327_Select_17_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_327_Select_16_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [16]), .I3(GND_net), .O(n3_adj_4045));
    defparam select_327_Select_16_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_327_Select_15_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [15]), .I3(GND_net), .O(n3_adj_4044));
    defparam select_327_Select_15_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1374 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [12]), 
            .I3(GND_net), .O(n36819));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1374.LUT_INIT = 16'he0e0;
    SB_LUT4 select_327_Select_14_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [14]), .I3(GND_net), .O(n3_adj_4043));
    defparam select_327_Select_14_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_327_Select_13_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [13]), .I3(GND_net), .O(n3_adj_4042));
    defparam select_327_Select_13_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_327_Select_12_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [12]), .I3(GND_net), .O(n3_adj_4041));
    defparam select_327_Select_12_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_327_Select_11_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [11]), .I3(GND_net), .O(n3_adj_4040));
    defparam select_327_Select_11_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_327_Select_10_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [10]), .I3(GND_net), .O(n3_adj_4039));
    defparam select_327_Select_10_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_327_Select_9_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [9]), .I3(GND_net), .O(n3_adj_4038));
    defparam select_327_Select_9_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_327_Select_8_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [8]), .I3(GND_net), .O(n3_adj_4037));
    defparam select_327_Select_8_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_4_lut_adj_1375 (.I0(n326), .I1(n200), .I2(n324), 
            .I3(\FRAME_MATCHER.state [29]), .O(n8_adj_4088));
    defparam i1_2_lut_4_lut_adj_1375.LUT_INIT = 16'hfe00;
    SB_LUT4 select_327_Select_7_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [7]), .I3(GND_net), .O(n3_adj_4036));
    defparam select_327_Select_7_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 n45914_bdd_4_lut (.I0(n45914), .I1(n17_adj_4158), .I2(n16_adj_4157), 
            .I3(byte_transmit_counter[2]), .O(n45917));
    defparam n45914_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1376 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [11]), 
            .I3(GND_net), .O(n36815));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1376.LUT_INIT = 16'he0e0;
    SB_LUT4 select_327_Select_6_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [6]), .I3(GND_net), .O(n3_adj_4035));
    defparam select_327_Select_6_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i4_4_lut_adj_1377 (.I0(\data_in_frame[19] [3]), .I1(n37881), 
            .I2(n37536), .I3(\data_in_frame[14] [5]), .O(n10_adj_4174));   // verilog/coms.v(76[16:27])
    defparam i4_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 select_327_Select_5_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [5]), .I3(GND_net), .O(n3_adj_4034));
    defparam select_327_Select_5_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_327_Select_4_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [4]), .I3(GND_net), .O(n3_adj_4033));
    defparam select_327_Select_4_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_327_Select_3_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n3_adj_4032));
    defparam select_327_Select_3_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_38786 (.I0(byte_transmit_counter[1]), 
            .I1(n19_adj_4156), .I2(n42818), .I3(byte_transmit_counter[2]), 
            .O(n45908));
    defparam byte_transmit_counter_1__bdd_4_lut_38786.LUT_INIT = 16'he4aa;
    SB_LUT4 i5_3_lut_4_lut_adj_1378 (.I0(n17696), .I1(\data_in_frame[17] [0]), 
            .I2(n10_adj_3996), .I3(\data_in_frame[16] [5]), .O(n37545));
    defparam i5_3_lut_4_lut_adj_1378.LUT_INIT = 16'h6996;
    SB_LUT4 select_327_Select_2_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [2]), .I3(GND_net), .O(n3_adj_4030));
    defparam select_327_Select_2_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_3_lut_4_lut_adj_1379 (.I0(\data_in_frame[15] [4]), .I1(n17928), 
            .I2(n37754), .I3(\data_in_frame[17] [5]), .O(n37555));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_4_lut_adj_1379.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1380 (.I0(n33850), .I1(n37690), .I2(n33852), 
            .I3(n33087), .O(n37956));
    defparam i1_2_lut_4_lut_adj_1380.LUT_INIT = 16'h6996;
    SB_LUT4 select_327_Select_1_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [1]), .I3(GND_net), .O(n3_adj_4029));
    defparam select_327_Select_1_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 select_327_Select_0_i3_2_lut_3_lut (.I0(n27114), .I1(n17201), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n3));
    defparam select_327_Select_0_i3_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i14241_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37354), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n19273));
    defparam i14241_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14242_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37354), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n19274));
    defparam i14242_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1381 (.I0(\data_in_frame[6] [2]), .I1(\data_in_frame[12] [5]), 
            .I2(\data_in_frame[8] [3]), .I3(\data_in_frame[10] [4]), .O(n14_adj_3995));   // verilog/coms.v(71[16:42])
    defparam i5_3_lut_4_lut_adj_1381.LUT_INIT = 16'h6996;
    SB_LUT4 i14243_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37354), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n19275));
    defparam i14243_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14244_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37354), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n19276));
    defparam i14244_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n45908_bdd_4_lut (.I0(n45908), .I1(n17_adj_4155), .I2(n16_adj_4154), 
            .I3(byte_transmit_counter[2]), .O(n45911));
    defparam n45908_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_3_lut_adj_1382 (.I0(n37661), .I1(n10_adj_4174), .I2(n17445), 
            .I3(GND_net), .O(n37643));   // verilog/coms.v(76[16:27])
    defparam i5_3_lut_adj_1382.LUT_INIT = 16'h9696;
    SB_LUT4 i14245_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37354), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n19277));
    defparam i14245_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14246_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37354), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n19278));
    defparam i14246_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14247_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37354), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n19279));
    defparam i14247_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14248_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37354), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n19280));
    defparam i14248_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_38781 (.I0(byte_transmit_counter[1]), 
            .I1(n19_adj_4152), .I2(n42811), .I3(byte_transmit_counter[2]), 
            .O(n45902));
    defparam byte_transmit_counter_1__bdd_4_lut_38781.LUT_INIT = 16'he4aa;
    SB_LUT4 i14121_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37361), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n19153));
    defparam i14121_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14122_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37361), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n19154));
    defparam i14122_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14123_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37361), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n19155));
    defparam i14123_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14124_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37361), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n19156));
    defparam i14124_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14125_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37361), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n19157));
    defparam i14125_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_3_lut_adj_1383 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[3] [7]), 
            .I2(\data_in_frame[6] [0]), .I3(GND_net), .O(n10_adj_3993));   // verilog/coms.v(94[12:25])
    defparam i2_2_lut_3_lut_adj_1383.LUT_INIT = 16'h9696;
    SB_LUT4 i14126_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37361), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n19158));
    defparam i14126_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1384 (.I0(\data_in_frame[14] [5]), .I1(n17696), 
            .I2(n37536), .I3(GND_net), .O(n33087));
    defparam i1_2_lut_3_lut_adj_1384.LUT_INIT = 16'h9696;
    SB_LUT4 i14127_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37361), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n19159));
    defparam i14127_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14128_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37361), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n19160));
    defparam i14128_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n45902_bdd_4_lut (.I0(n45902), .I1(n17_adj_4151), .I2(n16_adj_4150), 
            .I3(byte_transmit_counter[2]), .O(n45905));
    defparam n45902_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1385 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [5]), .I3(\data_in_frame[0] [6]), .O(n14_adj_4175));
    defparam i6_4_lut_adj_1385.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_4_lut_adj_1386 (.I0(\data_in_frame[9] [6]), .I1(n17687), 
            .I2(n37436), .I3(\data_in_frame[10] [2]), .O(n6_adj_3990));
    defparam i1_2_lut_4_lut_adj_1386.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1387 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [10]), 
            .I3(GND_net), .O(n36811));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1387.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_4_lut_adj_1388 (.I0(\data_in_frame[4] [4]), .I1(\data_in_frame[0] [0]), 
            .I2(n37511), .I3(n4_adj_3980), .O(n17492));   // verilog/coms.v(72[16:43])
    defparam i2_3_lut_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1389 (.I0(\data_in_frame[14] [7]), .I1(\data_in_frame[15] [1]), 
            .I2(\data_in_frame[6] [3]), .I3(GND_net), .O(n10_adj_3984));   // verilog/coms.v(70[16:41])
    defparam i2_2_lut_3_lut_adj_1389.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1033_i6_3_lut (.I0(\data_in_frame[16] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n4658), .I3(GND_net), .O(n4664));
    defparam mux_1033_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1390 (.I0(\data_in_frame[3] [5]), .I1(n37564), 
            .I2(\data_in_frame[6] [0]), .I3(\data_in_frame[8] [1]), .O(n37436));   // verilog/coms.v(70[16:41])
    defparam i1_2_lut_4_lut_adj_1390.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1033_i5_3_lut (.I0(\data_in_frame[16] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n4658), .I3(GND_net), .O(n4663));
    defparam mux_1033_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1391 (.I0(\data_in_frame[5] [5]), .I1(\data_in_frame[1] [1]), 
            .I2(\data_in_frame[3] [3]), .I3(\data_in_frame[0] [7]), .O(n37795));   // verilog/coms.v(71[16:34])
    defparam i1_2_lut_4_lut_adj_1391.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1392 (.I0(\data_in_frame[16] [7]), .I1(\data_in_frame[16] [6]), 
            .I2(\data_in_frame[16] [2]), .I3(\data_in_frame[16] [1]), .O(n37760));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_4_lut_adj_1392.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1033_i4_3_lut (.I0(\data_in_frame[16] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n4658), .I3(GND_net), .O(n4662));
    defparam mux_1033_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21274_2_lut_3_lut (.I0(n27114), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n26281));
    defparam i21274_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_3_lut_adj_1393 (.I0(\FRAME_MATCHER.state [2]), .I1(n17045), 
            .I2(n17263), .I3(GND_net), .O(n17264));   // verilog/coms.v(244[5:25])
    defparam i1_2_lut_3_lut_adj_1393.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1394 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_4176));   // verilog/coms.v(110[11:16])
    defparam i1_2_lut_adj_1394.LUT_INIT = 16'heeee;
    SB_LUT4 i31117_4_lut (.I0(n27475), .I1(\FRAME_MATCHER.state[3] ), .I2(\FRAME_MATCHER.state [2]), 
            .I3(n44_adj_4176), .O(n38178));
    defparam i31117_4_lut.LUT_INIT = 16'heeea;
    SB_LUT4 i35957_3_lut (.I0(n27475), .I1(\FRAME_MATCHER.state [1]), .I2(\FRAME_MATCHER.state[0] ), 
            .I3(GND_net), .O(n43081));
    defparam i35957_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 mux_715_i1_4_lut (.I0(Kp_23__N_718), .I1(n3086[0]), .I2(\FRAME_MATCHER.state [1]), 
            .I3(\FRAME_MATCHER.state[0] ), .O(n3139[0]));   // verilog/coms.v(147[4] 288[11])
    defparam mux_715_i1_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i35959_4_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(n3139[0]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(n43081), .O(n43083));   // verilog/coms.v(147[4] 288[11])
    defparam i35959_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i1_2_lut_3_lut_adj_1395 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [9]), 
            .I3(GND_net), .O(n36803));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1395.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_38776 (.I0(byte_transmit_counter[1]), 
            .I1(n19_adj_4149), .I2(n42810), .I3(byte_transmit_counter[2]), 
            .O(n45896));
    defparam byte_transmit_counter_1__bdd_4_lut_38776.LUT_INIT = 16'he4aa;
    SB_LUT4 n45896_bdd_4_lut (.I0(n45896), .I1(n17_adj_4148), .I2(n16_adj_4147), 
            .I3(byte_transmit_counter[2]), .O(n45899));
    defparam n45896_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_4_lut_adj_1396 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(\data_in_frame[0] [1]), .O(n13_adj_4177));
    defparam i5_4_lut_adj_1396.LUT_INIT = 16'h8000;
    SB_LUT4 i36242_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n43367));   // verilog/coms.v(104[34:55])
    defparam i36242_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4178));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33806_4_lut (.I0(n5_adj_4178), .I1(n43367), .I2(n26492), 
            .I3(byte_transmit_counter[0]), .O(n40930));
    defparam i33806_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i33808_4_lut (.I0(n40930), .I1(n45917), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n40932));
    defparam i33808_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i33807_3_lut (.I0(n45977), .I1(n45971), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n40931));
    defparam i33807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36237_2_lut (.I0(byte_transmit_counter[2]), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n43362));   // verilog/coms.v(104[34:55])
    defparam i36237_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_3_lut_adj_1397 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [8]), 
            .I3(GND_net), .O(n36799));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1397.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1398 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [7]), 
            .I3(GND_net), .O(n36795));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1398.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4179));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33803_4_lut (.I0(n5_adj_4179), .I1(n43362), .I2(n26492), 
            .I3(byte_transmit_counter[0]), .O(n40927));
    defparam i33803_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i33805_4_lut (.I0(n40927), .I1(n45899), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n40929));
    defparam i33805_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i33804_3_lut (.I0(n45989), .I1(n45983), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n40928));
    defparam i33804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1399 (.I0(\FRAME_MATCHER.state [1]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n17045), .I3(GND_net), .O(n17199));   // verilog/coms.v(195[5:24])
    defparam i1_2_lut_3_lut_adj_1399.LUT_INIT = 16'hfefe;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(byte_transmit_counter[1]), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n43357));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4180));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33800_4_lut (.I0(n5_adj_4180), .I1(byte_transmit_counter[0]), 
            .I2(n26492), .I3(n43357), .O(n40924));
    defparam i33800_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i33802_4_lut (.I0(n40924), .I1(n45905), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n40926));
    defparam i33802_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i33801_3_lut (.I0(n46001), .I1(n45995), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n40925));
    defparam i33801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37612_4_lut (.I0(n45929), .I1(n45911), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(tx_data[4]));   // verilog/coms.v(104[34:55])
    defparam i37612_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i36220_2_lut (.I0(\data_out_frame[0][3] ), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n42914));   // verilog/coms.v(104[34:55])
    defparam i36220_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(n42914), .I2(byte_transmit_counter[2]), .I3(byte_transmit_counter[0]), 
            .O(n6_adj_4181));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf0c;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n5_adj_4182));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33797_3_lut (.I0(n5_adj_4182), .I1(n6_adj_4181), .I2(n26492), 
            .I3(GND_net), .O(n40921));
    defparam i33797_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i33799_4_lut (.I0(n40921), .I1(n45923), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(n40923));
    defparam i33799_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i33798_3_lut (.I0(n46013), .I1(n46007), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n40922));
    defparam i33798_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13767_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37361), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n18799));
    defparam i13767_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14114_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37361), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n19146));
    defparam i14114_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14115_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37361), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n19147));
    defparam i14115_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14116_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37361), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n19148));
    defparam i14116_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14117_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37361), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n19149));
    defparam i14117_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i36308_2_lut (.I0(\data_out_frame[0] [2]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n42930));
    defparam i36308_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i33840_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n40964));
    defparam i33840_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i19_3_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\data_out_frame[21] [2]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_4183));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33816_4_lut (.I0(n19_adj_4183), .I1(\data_out_frame[22] [2]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n40940));
    defparam i33816_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i33841_4_lut (.I0(n40964), .I1(n42930), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n40965));
    defparam i33841_4_lut.LUT_INIT = 16'ha0ac;
    SB_LUT4 i33839_3_lut (.I0(\data_out_frame[4][2] ), .I1(\data_out_frame[5] [2]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n40963));
    defparam i33839_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37364_3_lut (.I0(n46019), .I1(n45893), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n44489));
    defparam i37364_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_38804 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(byte_transmit_counter[1]), .O(n45890));
    defparam byte_transmit_counter_0__bdd_4_lut_38804.LUT_INIT = 16'he4aa;
    SB_LUT4 i33817_3_lut (.I0(n45953), .I1(n40940), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n40941));
    defparam i33817_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37609_3_lut (.I0(n40918), .I1(n44489), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n44734));   // verilog/coms.v(104[34:55])
    defparam i37609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37610_4_lut (.I0(n44734), .I1(n40941), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(tx_data[2]));   // verilog/coms.v(104[34:55])
    defparam i37610_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14118_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37361), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n19150));
    defparam i14118_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14119_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37361), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n19151));
    defparam i14119_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14120_3_lut_4_lut (.I0(n8_adj_3907), .I1(n37361), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n19152));
    defparam i14120_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14207_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37342), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n19239));
    defparam i14207_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14208_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37342), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n19240));
    defparam i14208_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i36105_2_lut (.I0(\data_out_frame[0] [1]), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n42938));
    defparam i36105_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i33831_3_lut (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[7] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n40955));
    defparam i33831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i19_3_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\data_out_frame[21] [1]), .I2(byte_transmit_counter[0]), 
            .I3(GND_net), .O(n19_adj_4184));   // verilog/coms.v(104[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33813_4_lut (.I0(n19_adj_4184), .I1(\data_out_frame[22] [1]), 
            .I2(byte_transmit_counter[1]), .I3(byte_transmit_counter[0]), 
            .O(n40937));
    defparam i33813_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i33832_4_lut (.I0(n40955), .I1(n42938), .I2(byte_transmit_counter[2]), 
            .I3(byte_transmit_counter[0]), .O(n40956));
    defparam i33832_4_lut.LUT_INIT = 16'hafac;
    SB_LUT4 i33830_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n40954));
    defparam i33830_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37366_3_lut (.I0(n46025), .I1(n45887), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n44491));
    defparam i37366_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1400 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [6]), 
            .I3(GND_net), .O(n36791));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1400.LUT_INIT = 16'he0e0;
    SB_LUT4 i33814_3_lut (.I0(n45947), .I1(n40937), .I2(byte_transmit_counter[2]), 
            .I3(GND_net), .O(n40938));
    defparam i33814_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37607_3_lut (.I0(n40915), .I1(n44491), .I2(byte_transmit_counter[3]), 
            .I3(GND_net), .O(n44732));   // verilog/coms.v(104[34:55])
    defparam i37607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37608_4_lut (.I0(n44732), .I1(n40938), .I2(byte_transmit_counter[4]), 
            .I3(byte_transmit_counter[3]), .O(tx_data[1]));   // verilog/coms.v(104[34:55])
    defparam i37608_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i14205_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37342), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n19237));
    defparam i14205_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14206_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37342), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n19238));
    defparam i14206_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n45890_bdd_4_lut (.I0(n45890), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(byte_transmit_counter[1]), 
            .O(n45893));
    defparam n45890_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i14201_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37342), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n19233));
    defparam i14201_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14202_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37342), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n19234));
    defparam i14202_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14203_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37342), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n19235));
    defparam i14203_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14204_3_lut_4_lut (.I0(n8_adj_4166), .I1(n37342), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n19236));
    defparam i14204_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1401 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [5]), 
            .I3(GND_net), .O(n36787));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1401.LUT_INIT = 16'he0e0;
    SB_LUT4 i14193_3_lut_4_lut (.I0(n8), .I1(n37342), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n19225));
    defparam i14193_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1402 (.I0(n322), .I1(n301), .I2(\FRAME_MATCHER.state [4]), 
            .I3(GND_net), .O(n36783));   // verilog/coms.v(113[11:12])
    defparam i1_2_lut_3_lut_adj_1402.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut_adj_1403 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [28]), .O(n36635));
    defparam i1_2_lut_4_lut_adj_1403.LUT_INIT = 16'hba00;
    SB_LUT4 i1_2_lut_4_lut_adj_1404 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [26]), .O(n36637));
    defparam i1_2_lut_4_lut_adj_1404.LUT_INIT = 16'hba00;
    SB_LUT4 i14194_3_lut_4_lut (.I0(n8), .I1(n37342), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n19226));
    defparam i14194_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14195_3_lut_4_lut (.I0(n8), .I1(n37342), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n19227));
    defparam i14195_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14196_3_lut_4_lut (.I0(n8), .I1(n37342), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n19228));
    defparam i14196_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14197_3_lut_4_lut (.I0(n8), .I1(n37342), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n19229));
    defparam i14197_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14198_3_lut_4_lut (.I0(n8), .I1(n37342), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n19230));
    defparam i14198_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14199_3_lut_4_lut (.I0(n8), .I1(n37342), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n19231));
    defparam i14199_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14200_3_lut_4_lut (.I0(n8), .I1(n37342), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n19232));
    defparam i14200_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 Kp_23__I_831_3_lut (.I0(Kp_23__N_1746), .I1(n13_adj_4177), .I2(n14_adj_4175), 
            .I3(GND_net), .O(Kp_23__N_1745));   // verilog/coms.v(232[12:65])
    defparam Kp_23__I_831_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i14210_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37342), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n19242));
    defparam i14210_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14211_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37342), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n19243));
    defparam i14211_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14212_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37342), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n19244));
    defparam i14212_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14213_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37342), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n19245));
    defparam i14213_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1405 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [25]), .O(n36693));
    defparam i1_2_lut_4_lut_adj_1405.LUT_INIT = 16'hba00;
    SB_LUT4 i1_2_lut_4_lut_adj_1406 (.I0(n326), .I1(n200), .I2(n324), 
            .I3(\FRAME_MATCHER.state [27]), .O(n8_adj_4086));
    defparam i1_2_lut_4_lut_adj_1406.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1407 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [24]), .O(n36639));
    defparam i1_2_lut_4_lut_adj_1407.LUT_INIT = 16'hba00;
    SB_LUT4 i1_2_lut_4_lut_adj_1408 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [22]), .O(n36641));
    defparam i1_2_lut_4_lut_adj_1408.LUT_INIT = 16'hba00;
    SB_LUT4 i14214_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37342), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n19246));
    defparam i14214_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14215_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37342), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n19247));
    defparam i14215_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14216_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37342), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n19248));
    defparam i14216_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_4_lut_adj_1409 (.I0(\data_in_frame[18] [5]), .I1(n37410), 
            .I2(\data_in_frame[20] [7]), .I3(n32982), .O(n12_adj_4025));
    defparam i5_4_lut_adj_1409.LUT_INIT = 16'h6996;
    SB_LUT4 i14209_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37342), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n19241));
    defparam i14209_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14145_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37361), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n19177));
    defparam i14145_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14146_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37361), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n19178));
    defparam i14146_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14147_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37361), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n19179));
    defparam i14147_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1410 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [21]), .O(n36653));
    defparam i1_2_lut_4_lut_adj_1410.LUT_INIT = 16'hba00;
    SB_LUT4 i14148_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37361), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n19180));
    defparam i14148_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14149_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37361), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n19181));
    defparam i14149_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14150_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37361), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n19182));
    defparam i14150_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14151_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37361), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n19183));
    defparam i14151_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1411 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [20]), .O(n36683));
    defparam i1_2_lut_4_lut_adj_1411.LUT_INIT = 16'hba00;
    SB_LUT4 i14152_3_lut_4_lut (.I0(n8_adj_3947), .I1(n37361), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n19184));
    defparam i14152_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1412 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [19]), .O(n36579));
    defparam i1_2_lut_4_lut_adj_1412.LUT_INIT = 16'hba00;
    SB_LUT4 i1_2_lut_3_lut_adj_1413 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[3] [5]), 
            .I2(n37567), .I3(GND_net), .O(n7_adj_4098));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1413.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1414 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [16]), .O(n36603));
    defparam i1_2_lut_4_lut_adj_1414.LUT_INIT = 16'hba00;
    SB_LUT4 i2_3_lut_4_lut_adj_1415 (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(n37798), .I3(n17664), .O(n38745));
    defparam i2_3_lut_4_lut_adj_1415.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1416 (.I0(\data_out_frame[18] [4]), .I1(n33845), 
            .I2(n39208), .I3(GND_net), .O(n17664));
    defparam i1_2_lut_3_lut_adj_1416.LUT_INIT = 16'h6969;
    SB_LUT4 i2_2_lut_4_lut_adj_1417 (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[6] [7]), .I3(\data_out_frame[12] [1]), .O(n10_adj_3979));
    defparam i2_2_lut_4_lut_adj_1417.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1418 (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[6] [7]), .I3(GND_net), .O(n37842));
    defparam i1_2_lut_3_lut_adj_1418.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1419 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(n37422), .I3(\data_out_frame[13] [6]), .O(n37407));
    defparam i2_3_lut_4_lut_adj_1419.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1420 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[12] [0]), .I3(n39794), .O(n37977));
    defparam i1_2_lut_4_lut_adj_1420.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1421 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[8] [5]), .I3(GND_net), .O(n37677));
    defparam i1_2_lut_3_lut_adj_1421.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1422 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[7] [6]), .I3(\data_out_frame[7] [7]), .O(n17725));
    defparam i1_2_lut_4_lut_adj_1422.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1423 (.I0(n17764), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[9] [3]), .I3(\data_out_frame[9] [2]), .O(n37827));
    defparam i1_2_lut_4_lut_adj_1423.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1424 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[9] [2]), .I3(GND_net), .O(n18073));
    defparam i1_2_lut_3_lut_adj_1424.LUT_INIT = 16'h9696;
    SB_LUT4 i14185_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37342), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n19217));
    defparam i14185_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14186_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37342), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n19218));
    defparam i14186_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1425 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [14]), .O(n36643));
    defparam i1_2_lut_4_lut_adj_1425.LUT_INIT = 16'hba00;
    SB_LUT4 i2_3_lut_4_lut_adj_1426 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[8] [3]), 
            .I2(\data_out_frame[8] [4]), .I3(\data_out_frame[8] [5]), .O(n17365));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1426.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1427 (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[8] [0]), 
            .I2(n17725), .I3(GND_net), .O(n6_adj_3967));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_3_lut_adj_1427.LUT_INIT = 16'h9696;
    SB_LUT4 i14187_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37342), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n19219));
    defparam i14187_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1428 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [13]), .O(n36645));
    defparam i1_2_lut_4_lut_adj_1428.LUT_INIT = 16'hba00;
    SB_LUT4 i1_2_lut_3_lut_adj_1429 (.I0(\data_in_frame[5] [0]), .I1(n37489), 
            .I2(n37710), .I3(GND_net), .O(n33886));
    defparam i1_2_lut_3_lut_adj_1429.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1430 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[7] [5]), 
            .I2(\data_out_frame[9] [6]), .I3(\data_out_frame[8] [0]), .O(n17330));   // verilog/coms.v(83[17:28])
    defparam i1_2_lut_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1431 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[5] [5]), .I3(GND_net), .O(n18031));
    defparam i1_2_lut_3_lut_adj_1431.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1432 (.I0(n326), .I1(n200), .I2(n324), 
            .I3(\FRAME_MATCHER.state [23]), .O(n8_adj_4083));
    defparam i1_2_lut_4_lut_adj_1432.LUT_INIT = 16'hfe00;
    SB_LUT4 i14188_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37342), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n19220));
    defparam i14188_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1433 (.I0(n326), .I1(n200), .I2(n324), 
            .I3(\FRAME_MATCHER.state [18]), .O(n8_adj_4080));
    defparam i1_2_lut_4_lut_adj_1433.LUT_INIT = 16'hfe00;
    SB_LUT4 i14189_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37342), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n19221));
    defparam i14189_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14190_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37342), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n19222));
    defparam i14190_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14191_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37342), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n19223));
    defparam i14191_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1434 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [12]), .O(n36647));
    defparam i1_2_lut_4_lut_adj_1434.LUT_INIT = 16'hba00;
    SB_LUT4 i14192_3_lut_4_lut (.I0(n8_adj_4167), .I1(n37342), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n19224));
    defparam i14192_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1435 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [11]), .O(n36649));
    defparam i1_2_lut_4_lut_adj_1435.LUT_INIT = 16'hba00;
    SB_LUT4 i2_3_lut_4_lut_adj_1436 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[5] [5]), .I3(\data_out_frame[9] [7]), .O(n17742));
    defparam i2_3_lut_4_lut_adj_1436.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1437 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[5] [4]), .I3(GND_net), .O(n17764));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1437.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1438 (.I0(\data_out_frame[16] [0]), .I1(n37404), 
            .I2(n10_adj_3942), .I3(\data_out_frame[15] [7]), .O(n37807));
    defparam i1_2_lut_4_lut_adj_1438.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1439 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [10]), .O(n36651));
    defparam i1_2_lut_4_lut_adj_1439.LUT_INIT = 16'hba00;
    SB_LUT4 i1_2_lut_4_lut_adj_1440 (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(\data_out_frame[6] [5]), .I3(\data_out_frame[9] [1]), .O(n6_adj_3940));
    defparam i1_2_lut_4_lut_adj_1440.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1441 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[9] [1]), .I3(GND_net), .O(n37814));
    defparam i1_2_lut_3_lut_adj_1441.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1442 (.I0(n17979), .I1(n37496), .I2(n37575), 
            .I3(GND_net), .O(n32716));
    defparam i1_2_lut_3_lut_adj_1442.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1443 (.I0(\data_out_frame[17] [4]), .I1(\data_out_frame[13] [2]), 
            .I2(n16787), .I3(GND_net), .O(n6_adj_3937));
    defparam i1_2_lut_3_lut_adj_1443.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1444 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [9]), .O(n36655));
    defparam i1_2_lut_4_lut_adj_1444.LUT_INIT = 16'hba00;
    SB_LUT4 i1_2_lut_4_lut_adj_1445 (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[7] [6]), .I3(\data_out_frame[7] [7]), .O(n37572));
    defparam i1_2_lut_4_lut_adj_1445.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1446 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[7] [7]), .I3(GND_net), .O(n18082));   // verilog/coms.v(73[16:27])
    defparam i1_2_lut_3_lut_adj_1446.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1447 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[8] [0]), 
            .I2(\data_out_frame[6] [0]), .I3(\data_out_frame[8] [2]), .O(n18079));   // verilog/coms.v(71[16:42])
    defparam i2_3_lut_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1448 (.I0(n326), .I1(n200), .I2(n324), 
            .I3(\FRAME_MATCHER.state [17]), .O(n8_adj_4078));
    defparam i1_2_lut_4_lut_adj_1448.LUT_INIT = 16'hfe00;
    SB_LUT4 i5_3_lut_4_lut_adj_1449 (.I0(\data_out_frame[4][0] ), .I1(\data_out_frame[6] [1]), 
            .I2(n10_adj_3936), .I3(\data_out_frame[12] [7]), .O(n1595));   // verilog/coms.v(70[16:27])
    defparam i5_3_lut_4_lut_adj_1449.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1450 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [8]), .O(n36657));
    defparam i1_2_lut_4_lut_adj_1450.LUT_INIT = 16'hba00;
    SB_LUT4 i2_3_lut_4_lut_adj_1451 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(n17742), .I3(\data_out_frame[7] [4]), .O(n37501));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1451.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1452 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [7]), .O(n36659));
    defparam i1_2_lut_4_lut_adj_1452.LUT_INIT = 16'hba00;
    SB_LUT4 i4_2_lut_4_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[14] [3]), 
            .I2(\data_out_frame[14] [6]), .I3(\data_out_frame[14] [7]), 
            .O(n15));
    defparam i4_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1453 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [2]), 
            .I2(\data_out_frame[11] [6]), .I3(\data_out_frame[9] [5]), .O(n37520));   // verilog/coms.v(72[16:27])
    defparam i2_3_lut_4_lut_adj_1453.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_38767 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(byte_transmit_counter[1]), .O(n45884));
    defparam byte_transmit_counter_0__bdd_4_lut_38767.LUT_INIT = 16'he4aa;
    SB_LUT4 i5_3_lut_4_lut_adj_1454 (.I0(\data_in_frame[20] [4]), .I1(n10_adj_3924), 
            .I2(\data_in_frame[18] [3]), .I3(n16859), .O(n38695));
    defparam i5_3_lut_4_lut_adj_1454.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1455 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(n1119), .I3(\data_out_frame[5] [1]), .O(n14_adj_3969));   // verilog/coms.v(83[17:70])
    defparam i5_3_lut_4_lut_adj_1455.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1456 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(\data_out_frame[8] [7]), .I3(\data_out_frame[11] [3]), .O(n17916));   // verilog/coms.v(83[17:70])
    defparam i1_2_lut_3_lut_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 n45884_bdd_4_lut (.I0(n45884), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(byte_transmit_counter[1]), 
            .O(n45887));
    defparam n45884_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1457 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [6]), .O(n36601));
    defparam i1_2_lut_4_lut_adj_1457.LUT_INIT = 16'hba00;
    SB_LUT4 i6_4_lut_adj_1458 (.I0(n33880), .I1(n32943), .I2(n37857), 
            .I3(n17542), .O(n16_adj_4027));
    defparam i6_4_lut_adj_1458.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1459 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[6] [4]), 
            .I2(n37763), .I3(GND_net), .O(n17422));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1459.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1460 (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[4][0] ), .I3(n18209), .O(n37923));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1460.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1461 (.I0(\data_out_frame[4] [1]), .I1(n1287), 
            .I2(\data_out_frame[8] [5]), .I3(\data_out_frame[11] [1]), .O(n37884));
    defparam i2_3_lut_4_lut_adj_1461.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1462 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[4][0] ), 
            .I2(n37792), .I3(GND_net), .O(n6_adj_3943));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_adj_1462.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1463 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[4][0] ), 
            .I2(\data_out_frame[4][2] ), .I3(GND_net), .O(n37763));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_adj_1463.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_38762 (.I0(byte_transmit_counter[0]), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(byte_transmit_counter[1]), .O(n45878));
    defparam byte_transmit_counter_0__bdd_4_lut_38762.LUT_INIT = 16'he4aa;
    SB_LUT4 n45878_bdd_4_lut (.I0(n45878), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(byte_transmit_counter[1]), 
            .O(n45881));
    defparam n45878_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut_3_lut_4_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[14] [3]), 
            .I2(\data_out_frame[9] [4]), .I3(n37786), .O(n17_adj_3965));
    defparam i7_4_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1464 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[8] [3]), 
            .I2(\data_out_frame[8] [1]), .I3(n18292), .O(n37965));   // verilog/coms.v(71[16:42])
    defparam i2_3_lut_4_lut_adj_1464.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1465 (.I0(n326), .I1(n200), .I2(n324), 
            .I3(\FRAME_MATCHER.state [15]), .O(n8_adj_4076));
    defparam i1_2_lut_4_lut_adj_1465.LUT_INIT = 16'hfe00;
    SB_LUT4 i7_4_lut_adj_1466 (.I0(Kp_23__N_1433), .I1(n37732), .I2(n37953), 
            .I3(n17379), .O(n17_adj_4026));
    defparam i7_4_lut_adj_1466.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1467 (.I0(n324), .I1(n17183), .I2(n9), 
            .I3(\FRAME_MATCHER.state [5]), .O(n36599));
    defparam i1_2_lut_4_lut_adj_1467.LUT_INIT = 16'hba00;
    SB_LUT4 i1_2_lut_4_lut_adj_1468 (.I0(\data_out_frame[11] [5]), .I1(n17648), 
            .I2(n37575), .I3(n18143), .O(n32979));
    defparam i1_2_lut_4_lut_adj_1468.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1469 (.I0(n17638), .I1(\data_out_frame[13] [1]), 
            .I2(n1595), .I3(GND_net), .O(n37962));
    defparam i1_2_lut_3_lut_adj_1469.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1470 (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[16] [6]), 
            .I2(n17626), .I3(GND_net), .O(n37744));
    defparam i1_2_lut_3_lut_adj_1470.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1471 (.I0(\data_out_frame[17] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(n1642), .I3(GND_net), .O(n37872));
    defparam i1_2_lut_3_lut_adj_1471.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1472 (.I0(\data_out_frame[19] [5]), .I1(\data_out_frame[19] [4]), 
            .I2(n37869), .I3(n33049), .O(n38629));
    defparam i2_3_lut_4_lut_adj_1472.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_adj_1473 (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[8] [3]), 
            .I2(\data_out_frame[10] [4]), .I3(GND_net), .O(n37792));   // verilog/coms.v(71[16:42])
    defparam i1_2_lut_3_lut_adj_1473.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1474 (.I0(\data_out_frame[19] [7]), .I1(n17969), 
            .I2(n37707), .I3(GND_net), .O(n37640));
    defparam i1_2_lut_3_lut_adj_1474.LUT_INIT = 16'h9696;
    SB_LUT4 i14129_3_lut_4_lut (.I0(n8), .I1(n37361), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n19161));
    defparam i14129_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1475 (.I0(n33902), .I1(n33882), .I2(\data_out_frame[20] [5]), 
            .I3(\data_out_frame[20] [6]), .O(n39432));
    defparam i2_3_lut_4_lut_adj_1475.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1476 (.I0(\FRAME_MATCHER.state [1]), .I1(n63_c), 
            .I2(n63_adj_3909), .I3(GND_net), .O(n93[1]));   // verilog/coms.v(126[12] 289[6])
    defparam i1_2_lut_3_lut_adj_1476.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1477 (.I0(n2664), .I1(n17265), .I2(n26317), 
            .I3(GND_net), .O(n37376));
    defparam i1_2_lut_3_lut_adj_1477.LUT_INIT = 16'habab;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1478 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[7] [3]), .I3(\data_out_frame[9] [4]), .O(n37496));
    defparam i1_2_lut_3_lut_4_lut_adj_1478.LUT_INIT = 16'h6996;
    SB_LUT4 i14130_3_lut_4_lut (.I0(n8), .I1(n37361), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n19162));
    defparam i14130_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_4_lut_adj_1479 (.I0(\data_in_frame[17] [7]), .I1(Kp_23__N_1562), 
            .I2(n16859), .I3(n32982), .O(n8_adj_3906));
    defparam i2_2_lut_4_lut_adj_1479.LUT_INIT = 16'h6996;
    uart_tx tx (.n18758(n18758), .clk32MHz(clk32MHz), .n18755(n18755), 
            .n18752(n18752), .n18749(n18749), .n19426(n19426), .r_SM_Main({r_SM_Main}), 
            .n18746(n18746), .n18767(n18767), .n18764(n18764), .n18761(n18761), 
            .n18744(n18744), .n18747(n18747), .\r_SM_Main_2__N_3323[0] (r_SM_Main_2__N_3323[0]), 
            .\r_SM_Main_2__N_3320[1] (\r_SM_Main_2__N_3320[1] ), .n18750(n18750), 
            .tx_data({tx_data}), .n18753(n18753), .n18756(n18756), .n18759(n18759), 
            .n18762(n18762), .n18765(n18765), .n18896(n18896), .VCC_net(VCC_net), 
            .GND_net(GND_net), .n18898(n18898), .n18816(n18816), .n18815(n18815), 
            .tx_active(tx_active), .n18814(n18814), .tx_o(tx_o), .n20(n20_adj_4106), 
            .tx_transmit_N_3215(tx_transmit_N_3215), .n26317(n26317), .n45935(n45935), 
            .tx_enable(tx_enable), .n18402(n18402), .n12501(n12501), .n18897(n18897)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(105[10:70])
    uart_rx rx (.n36985(n36985), .r_Clock_Count({\r_Clock_Count[7] , \r_Clock_Count[6] , 
            \r_Clock_Count[5] , \r_Clock_Count[4] , \r_Clock_Count[3] , 
            \r_Clock_Count[2] , \r_Clock_Count[1] , Open_0}), .clk32MHz(clk32MHz), 
            .n36987(n36987), .n36989(n36989), .n36919(n36919), .n36743(n36743), 
            .n36695(n36695), .n36983(n36983), .n18780(n18780), .r_Bit_Index({r_Bit_Index}), 
            .n18777(n18777), .n19419(n19419), .rx_data({rx_data}), .n27445(n27445), 
            .r_SM_Main({Open_1, \r_SM_Main[1]_adj_4 , Open_2}), .VCC_net(VCC_net), 
            .rx_data_ready(rx_data_ready), .GND_net(GND_net), .n95(n95), 
            .n16(n16), .\r_SM_Main[2] (\r_SM_Main[2]_adj_5 ), .r_Rx_Data(r_Rx_Data), 
            .PIN_13_N_105(PIN_13_N_105), .n37215(n37215), .n37220(n37220), 
            .n37217(n37217), .n37216(n37216), .n37218(n37218), .n37219(n37219), 
            .n37214(n37214), .n18943(n18943), .n18806(n18806), .n18793(n18793), 
            .n18786(n18786), .n18785(n18785), .n18784(n18784), .n18783(n18783), 
            .n18782(n18782), .n18781(n18781), .n42920(n42920), .n20874(n20874), 
            .n42919(n42919), .n17255(n17255), .n4(n4), .n26349(n26349), 
            .n4_adj_1(n4_adj_6), .n4_adj_2(n4_adj_7), .n17250(n17250), 
            .n4926(n4926), .n18467(n18467), .n20896(n20896), .n18602(n18602)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(91[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (n18758, clk32MHz, n18755, n18752, n18749, n19426, 
            r_SM_Main, n18746, n18767, n18764, n18761, n18744, n18747, 
            \r_SM_Main_2__N_3323[0] , \r_SM_Main_2__N_3320[1] , n18750, 
            tx_data, n18753, n18756, n18759, n18762, n18765, n18896, 
            VCC_net, GND_net, n18898, n18816, n18815, tx_active, 
            n18814, tx_o, n20, tx_transmit_N_3215, n26317, n45935, 
            tx_enable, n18402, n12501, n18897) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n18758;
    input clk32MHz;
    input n18755;
    input n18752;
    input n18749;
    input n19426;
    output [2:0]r_SM_Main;
    input n18746;
    input n18767;
    input n18764;
    input n18761;
    output n18744;
    output n18747;
    input \r_SM_Main_2__N_3323[0] ;
    output \r_SM_Main_2__N_3320[1] ;
    output n18750;
    input [7:0]tx_data;
    output n18753;
    output n18756;
    output n18759;
    output n18762;
    output n18765;
    output n18896;
    input VCC_net;
    input GND_net;
    input n18898;
    input n18816;
    input n18815;
    output tx_active;
    input n18814;
    output tx_o;
    input n20;
    output tx_transmit_N_3215;
    output n26317;
    output n45935;
    output tx_enable;
    output n18402;
    output n12501;
    output n18897;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n18771;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    
    wire n18774, n30354, n30353, n14689, n18473, n30352;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n30351, n30350, n30349, n30348, n30347, n1, n39583, n27403, 
        n36887, n39019, n5, n40999, n41000, n45932, n40943, n40942, 
        n7, n5_adj_3901, n10036, n42865;
    
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n18758));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n18755));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .D(n18752));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .D(n18749));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n19426));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), .D(n18746));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n18771));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n18767));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n18764));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n18761));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n18774));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_10_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[8]), 
            .I2(r_SM_Main[2]), .I3(n30354), .O(n18744)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_59_9_lut (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[7]), 
            .I2(r_SM_Main[2]), .I3(n30353), .O(n18747)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_9 (.CI(n30353), .I0(r_Clock_Count[7]), .I1(r_SM_Main[2]), 
            .CO(n30354));
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(\r_SM_Main_2__N_3323[0] ), 
            .I3(r_SM_Main[1]), .O(n14689));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3320[1] ), .O(n18473));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 add_59_8_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[6]), 
            .I2(r_SM_Main[2]), .I3(n30352), .O(n18750)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_8 (.CI(n30352), .I0(r_Clock_Count[6]), .I1(r_SM_Main[2]), 
            .CO(n30353));
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n14689), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_7_lut (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[5]), 
            .I2(r_SM_Main[2]), .I3(n30351), .O(n18753)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_7 (.CI(n30351), .I0(r_Clock_Count[5]), .I1(r_SM_Main[2]), 
            .CO(n30352));
    SB_LUT4 add_59_6_lut (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[4]), 
            .I2(r_SM_Main[2]), .I3(n30350), .O(n18756)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_6 (.CI(n30350), .I0(r_Clock_Count[4]), .I1(r_SM_Main[2]), 
            .CO(n30351));
    SB_LUT4 add_59_5_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[3]), 
            .I2(r_SM_Main[2]), .I3(n30349), .O(n18759)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_5 (.CI(n30349), .I0(r_Clock_Count[3]), .I1(r_SM_Main[2]), 
            .CO(n30350));
    SB_LUT4 add_59_4_lut (.I0(r_Clock_Count[2]), .I1(r_Clock_Count[2]), 
            .I2(r_SM_Main[2]), .I3(n30348), .O(n18762)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_4 (.CI(n30348), .I0(r_Clock_Count[2]), .I1(r_SM_Main[2]), 
            .CO(n30349));
    SB_LUT4 add_59_3_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[1]), 
            .I2(r_SM_Main[2]), .I3(n30347), .O(n18765)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_3 (.CI(n30347), .I0(r_Clock_Count[1]), .I1(r_SM_Main[2]), 
            .CO(n30348));
    SB_LUT4 add_59_2_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[0]), 
            .I2(r_SM_Main[2]), .I3(VCC_net), .O(n18896)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(r_SM_Main[2]), 
            .CO(n30347));
    SB_LUT4 i21414_2_lut (.I0(\r_SM_Main_2__N_3320[1] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n1));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i21414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut (.I0(n39583), .I1(r_Clock_Count[5]), .I2(r_Clock_Count[4]), 
            .I3(GND_net), .O(n27403));   // verilog/uart_tx.v(32[16:29])
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[1]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[0]), 
            .I3(r_Clock_Count[3]), .O(n39583));   // verilog/uart_tx.v(32[16:29])
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .D(n18898));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n36887));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n14689), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n14689), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n14689), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n14689), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n14689), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n14689), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n14689), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n18816));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n18815));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .D(n18814));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(n39019));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i38701_2_lut_3_lut (.I0(tx_active), .I1(\r_SM_Main_2__N_3323[0] ), 
            .I2(n20), .I3(GND_net), .O(tx_transmit_N_3215));
    defparam i38701_2_lut_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i21310_2_lut_3_lut (.I0(tx_active), .I1(\r_SM_Main_2__N_3323[0] ), 
            .I2(n20), .I3(GND_net), .O(n26317));
    defparam i21310_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i1_2_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(GND_net), .O(n5));   // verilog/uart_tx.v(32[16:29])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12_3_lut (.I0(n18473), .I1(r_Bit_Index[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n36887));   // verilog/uart_tx.v(31[16:25])
    defparam i12_3_lut.LUT_INIT = 16'h6464;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n40999), 
            .I2(n41000), .I3(r_Bit_Index[2]), .O(n45932));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n45932_bdd_4_lut (.I0(n45932), .I1(n40943), .I2(n40942), .I3(r_Bit_Index[2]), 
            .O(n45935));
    defparam n45932_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_868 (.I0(r_SM_Main[1]), .I1(n27403), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n7));
    defparam i2_3_lut_adj_868.LUT_INIT = 16'h3232;
    SB_LUT4 i3_3_lut_4_lut (.I0(\r_SM_Main_2__N_3320[1] ), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[2]), .I3(r_SM_Main[1]), .O(n39019));   // verilog/uart_tx.v(32[16:29])
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h0800;
    SB_LUT4 i33818_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n40942));
    defparam i33818_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33819_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n40943));
    defparam i33819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33876_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n41000));
    defparam i33876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33875_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n40999));
    defparam i33875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19664_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(tx_enable));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i19664_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24570_4_lut (.I0(n18473), .I1(r_SM_Main[1]), .I2(r_Bit_Index[1]), 
            .I3(r_Bit_Index[0]), .O(n18774));   // verilog/uart_tx.v(31[16:25])
    defparam i24570_4_lut.LUT_INIT = 16'h58d0;
    SB_LUT4 i1_2_lut_adj_869 (.I0(r_Bit_Index[0]), .I1(r_Bit_Index[1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3901));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut_adj_869.LUT_INIT = 16'h8888;
    SB_LUT4 i5260_2_lut (.I0(\r_SM_Main_2__N_3323[0] ), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n10036));   // verilog/uart_tx.v(43[7] 142[14])
    defparam i5260_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_4_lut (.I0(n10036), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(n1), .O(n18402));
    defparam i2_4_lut.LUT_INIT = 16'h3202;
    SB_LUT4 i36279_2_lut (.I0(\r_SM_Main_2__N_3320[1] ), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n42865));   // verilog/uart_tx.v(31[16:25])
    defparam i36279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i24556_4_lut (.I0(\r_SM_Main_2__N_3323[0] ), .I1(n42865), .I2(r_SM_Main[1]), 
            .I3(n5_adj_3901), .O(n12501));   // verilog/uart_tx.v(31[16:25])
    defparam i24556_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 i24564_4_lut (.I0(n18473), .I1(n5_adj_3901), .I2(r_SM_Main[1]), 
            .I3(r_Bit_Index[2]), .O(n18771));   // verilog/uart_tx.v(31[16:25])
    defparam i24564_4_lut.LUT_INIT = 16'h7580;
    SB_LUT4 i21402_4_lut (.I0(r_SM_Main[2]), .I1(n7), .I2(r_Clock_Count[6]), 
            .I3(n5), .O(n18897));
    defparam i21402_4_lut.LUT_INIT = 16'haaae;
    SB_LUT4 i3_3_lut_4_lut_adj_870 (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[7]), 
            .I2(r_Clock_Count[6]), .I3(n27403), .O(\r_SM_Main_2__N_3320[1] ));   // verilog/uart_tx.v(32[16:29])
    defparam i3_3_lut_4_lut_adj_870.LUT_INIT = 16'hfffe;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (n36985, r_Clock_Count, clk32MHz, n36987, n36989, n36919, 
            n36743, n36695, n36983, n18780, r_Bit_Index, n18777, 
            n19419, rx_data, n27445, r_SM_Main, VCC_net, rx_data_ready, 
            GND_net, n95, n16, \r_SM_Main[2] , r_Rx_Data, PIN_13_N_105, 
            n37215, n37220, n37217, n37216, n37218, n37219, n37214, 
            n18943, n18806, n18793, n18786, n18785, n18784, n18783, 
            n18782, n18781, n42920, n20874, n42919, n17255, n4, 
            n26349, n4_adj_1, n4_adj_2, n17250, n4926, n18467, n20896, 
            n18602) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n36985;
    output [7:0]r_Clock_Count;
    input clk32MHz;
    input n36987;
    input n36989;
    input n36919;
    input n36743;
    input n36695;
    input n36983;
    input n18780;
    output [2:0]r_Bit_Index;
    input n18777;
    input n19419;
    output [7:0]rx_data;
    input n27445;
    output [2:0]r_SM_Main;
    input VCC_net;
    output rx_data_ready;
    input GND_net;
    output n95;
    input n16;
    output \r_SM_Main[2] ;
    output r_Rx_Data;
    input PIN_13_N_105;
    output n37215;
    output n37220;
    output n37217;
    output n37216;
    output n37218;
    output n37219;
    output n37214;
    input n18943;
    input n18806;
    input n18793;
    input n18786;
    input n18785;
    input n18784;
    input n18783;
    input n18782;
    input n18781;
    output n42920;
    output n20874;
    output n42919;
    output n17255;
    output n4;
    output n26349;
    output n4_adj_1;
    output n4_adj_2;
    output n17250;
    output n4926;
    output n18467;
    output n20896;
    output n18602;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n36759, n117, n128;
    wire [7:0]r_Clock_Count_c;   // verilog/uart_rx.v(32[17:30])
    
    wire n130;
    wire [2:0]r_SM_Main_c;   // verilog/uart_rx.v(36[17:26])
    
    wire n93;
    wire [2:0]r_SM_Main_2__N_3249;
    
    wire n37213, n42989, n120, n37324, r_Rx_Data_R, n30346, n30345, 
        n30344, n18389, n30343, n30342, n30341, n30340;
    wire [31:0]n194;
    
    wire n24, n40, n17016, n26999;
    
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n36985));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n36987));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n36989));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n36919));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .D(n36743));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .D(n36695));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n36983));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n18780));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n18777));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n19419));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n27445));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFE r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .E(VCC_net), 
            .D(n36759));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[5]), .I1(r_Clock_Count[7]), .I2(r_Clock_Count[6]), 
            .I3(r_Clock_Count[4]), .O(n117));
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut (.I0(n117), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(GND_net), .O(n128));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i3_4_lut_adj_862 (.I0(r_Clock_Count[2]), .I1(n128), .I2(r_Clock_Count[1]), 
            .I3(r_Clock_Count_c[0]), .O(n130));
    defparam i3_4_lut_adj_862.LUT_INIT = 16'hdfff;
    SB_LUT4 i1_2_lut_adj_863 (.I0(r_SM_Main_c[0]), .I1(n130), .I2(GND_net), 
            .I3(GND_net), .O(n95));
    defparam i1_2_lut_adj_863.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_adj_864 (.I0(r_SM_Main_c[0]), .I1(n130), .I2(GND_net), 
            .I3(GND_net), .O(n93));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_adj_864.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(n93), .I1(n16), .I2(r_SM_Main_2__N_3249[2]), 
            .I3(r_SM_Main[1]), .O(n37213));
    defparam i1_4_lut.LUT_INIT = 16'h0322;
    SB_LUT4 i36524_3_lut_4_lut (.I0(r_Clock_Count_c[0]), .I1(r_Clock_Count[2]), 
            .I2(r_Clock_Count[1]), .I3(n128), .O(n42989));
    defparam i36524_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i2_2_lut_3_lut (.I0(r_Clock_Count_c[0]), .I1(r_Clock_Count[2]), 
            .I2(r_Clock_Count[1]), .I3(GND_net), .O(n120));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_DFFSR r_SM_Main_i2 (.Q(\r_SM_Main[2] ), .C(clk32MHz), .D(r_SM_Main_2__N_3249[2]), 
            .R(n37324));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(PIN_13_N_105));   // verilog/uart_rx.v(41[10] 45[8])
    SB_LUT4 add_62_9_lut (.I0(n37213), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n30346), .O(n37215)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_62_8_lut (.I0(n37213), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n30345), .O(n37220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_8 (.CI(n30345), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n30346));
    SB_LUT4 add_62_7_lut (.I0(n37213), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n30344), .O(n37217)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_7 (.CI(n30344), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n30345));
    SB_LUT4 i38707_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(\r_SM_Main[2] ), 
            .I2(r_SM_Main_c[0]), .I3(GND_net), .O(n37324));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i38707_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(\r_SM_Main[2] ), .I2(r_SM_Main_2__N_3249[2]), 
            .I3(r_SM_Main_c[0]), .O(n18389));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(\r_SM_Main[2] ), .I2(n18389), 
            .I3(rx_data_ready), .O(n36759));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    SB_LUT4 add_62_6_lut (.I0(n37213), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n30343), .O(n37216)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_6 (.CI(n30343), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n30344));
    SB_LUT4 add_62_5_lut (.I0(n37213), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n30342), .O(n37218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_5 (.CI(n30342), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n30343));
    SB_LUT4 add_62_4_lut (.I0(n37213), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n30341), .O(n37219)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_4 (.CI(n30341), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n30342));
    SB_LUT4 add_62_3_lut (.I0(n37213), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n30340), .O(n37214)) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_62_3 (.CI(n30340), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n30341));
    SB_LUT4 add_62_2_lut (.I0(GND_net), .I1(r_Clock_Count_c[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n194[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_2 (.CI(VCC_net), .I0(r_Clock_Count_c[0]), .I1(GND_net), 
            .CO(n30340));
    SB_DFFE r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .E(VCC_net), 
            .D(n18943));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count_c[0]), .C(clk32MHz), .D(n24));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main_c[0]), .C(clk32MHz), .D(n18806));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n18793));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n18786));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n18785));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n18784));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n18783));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n18782));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n18781));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i45_4_lut (.I0(n42989), .I1(r_SM_Main_2__N_3249[2]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_c[0]), .O(n40));
    defparam i45_4_lut.LUT_INIT = 16'hcacf;
    SB_LUT4 i38003_4_lut (.I0(n194[0]), .I1(r_Clock_Count_c[0]), .I2(n16), 
            .I3(n40), .O(n24));
    defparam i38003_4_lut.LUT_INIT = 16'hc0ca;
    SB_LUT4 i36278_2_lut (.I0(r_SM_Main_2__N_3249[2]), .I1(r_SM_Main_c[0]), 
            .I2(GND_net), .I3(GND_net), .O(n42920));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i36278_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15847_3_lut_3_lut (.I0(r_SM_Main_c[0]), .I1(n130), .I2(r_Rx_Data), 
            .I3(GND_net), .O(n20874));   // verilog/uart_rx.v(30[17:26])
    defparam i15847_3_lut_3_lut.LUT_INIT = 16'h8d8d;
    SB_LUT4 i36240_4_lut (.I0(r_SM_Main_c[0]), .I1(n128), .I2(r_Rx_Data), 
            .I3(n120), .O(n42919));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i36240_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i3_4_lut_adj_865 (.I0(\r_SM_Main[2] ), .I1(r_SM_Main_c[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main_2__N_3249[2]), .O(n17016));
    defparam i3_4_lut_adj_865.LUT_INIT = 16'hefff;
    SB_LUT4 i1_2_lut_adj_866 (.I0(r_Bit_Index[0]), .I1(n17016), .I2(GND_net), 
            .I3(GND_net), .O(n17255));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_866.LUT_INIT = 16'heeee;
    SB_LUT4 equal_127_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_127_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i21342_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n26349));
    defparam i21342_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_122_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_122_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_124_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_124_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_2_lut_adj_867 (.I0(n17016), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17250));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_867.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1228_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4926));   // verilog/uart_rx.v(102[36:51])
    defparam i1228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n26999));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut (.I0(n117), .I1(r_Clock_Count[3]), .I2(n120), .I3(GND_net), 
            .O(r_SM_Main_2__N_3249[2]));   // verilog/uart_rx.v(32[17:30])
    defparam i1_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main_c[0]), .I1(\r_SM_Main[2] ), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_3249[2]), .O(n18467));
    defparam i2_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i15869_3_lut (.I0(n26999), .I1(r_SM_Main_c[0]), .I2(r_SM_Main_2__N_3249[2]), 
            .I3(GND_net), .O(n20896));   // verilog/uart_rx.v(36[17:26])
    defparam i15869_3_lut.LUT_INIT = 16'h2c2c;
    SB_LUT4 i13570_3_lut (.I0(n18467), .I1(r_SM_Main[1]), .I2(n26999), 
            .I3(GND_net), .O(n18602));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13570_3_lut.LUT_INIT = 16'ha2a2;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (n19372, encoder0_position, clk32MHz, 
            n19373, n19374, n19375, n19376, n19377, n19368, n19369, 
            n19370, n19371, n19366, n19367, n19364, n19365, n19362, 
            n19363, n19360, n19361, n19358, n19359, n19355, n19356, 
            n19357, data_o, n2865, GND_net, n18802, count_enable, 
            n19406, reg_B, PIN_2_c_0, n18805, PIN_1_c_1, n39036) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n19372;
    output [23:0]encoder0_position;
    input clk32MHz;
    input n19373;
    input n19374;
    input n19375;
    input n19376;
    input n19377;
    input n19368;
    input n19369;
    input n19370;
    input n19371;
    input n19366;
    input n19367;
    input n19364;
    input n19365;
    input n19362;
    input n19363;
    input n19360;
    input n19361;
    input n19358;
    input n19359;
    input n19355;
    input n19356;
    input n19357;
    output [1:0]data_o;
    output [23:0]n2865;
    input GND_net;
    input n18802;
    output count_enable;
    input n19406;
    output [1:0]reg_B;
    input PIN_2_c_0;
    input n18805;
    input PIN_1_c_1;
    output n39036;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire B_delayed, A_delayed, n2861, n30401, n30400, n30399, n30398, 
        n30397, n30396, n30395, n30394, n30393, n30392, n30391, 
        n30390, n30389, n30388, n30387, n30386, n30385, n30384, 
        n30383, n30382, n30381, n30380, n30379, count_direction, 
        n30378;
    
    SB_DFF count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .D(n19372));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .D(n19373));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .D(n19374));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .D(n19375));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .D(n19376));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .D(n19377));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .D(n19368));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .D(n19369));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .D(n19370));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .D(n19371));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .D(n19366));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .D(n19367));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .D(n19364));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .D(n19365));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .D(n19362));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .D(n19363));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .D(n19360));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .D(n19361));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .D(n19358));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .D(n19359));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .D(n19355));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .D(n19356));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .D(n19357));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 add_617_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n2861), 
            .I3(n30401), .O(n2865[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_617_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n2861), 
            .I3(n30400), .O(n2865[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_24 (.CI(n30400), .I0(encoder0_position[22]), .I1(n2861), 
            .CO(n30401));
    SB_LUT4 add_617_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n2861), 
            .I3(n30399), .O(n2865[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_23 (.CI(n30399), .I0(encoder0_position[21]), .I1(n2861), 
            .CO(n30400));
    SB_LUT4 add_617_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n2861), 
            .I3(n30398), .O(n2865[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_22 (.CI(n30398), .I0(encoder0_position[20]), .I1(n2861), 
            .CO(n30399));
    SB_LUT4 add_617_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n2861), 
            .I3(n30397), .O(n2865[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_21 (.CI(n30397), .I0(encoder0_position[19]), .I1(n2861), 
            .CO(n30398));
    SB_LUT4 add_617_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n2861), 
            .I3(n30396), .O(n2865[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_20 (.CI(n30396), .I0(encoder0_position[18]), .I1(n2861), 
            .CO(n30397));
    SB_LUT4 add_617_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n2861), 
            .I3(n30395), .O(n2865[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_19 (.CI(n30395), .I0(encoder0_position[17]), .I1(n2861), 
            .CO(n30396));
    SB_LUT4 add_617_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n2861), 
            .I3(n30394), .O(n2865[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_18 (.CI(n30394), .I0(encoder0_position[16]), .I1(n2861), 
            .CO(n30395));
    SB_LUT4 add_617_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n2861), 
            .I3(n30393), .O(n2865[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_17 (.CI(n30393), .I0(encoder0_position[15]), .I1(n2861), 
            .CO(n30394));
    SB_LUT4 add_617_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n2861), 
            .I3(n30392), .O(n2865[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_16 (.CI(n30392), .I0(encoder0_position[14]), .I1(n2861), 
            .CO(n30393));
    SB_LUT4 add_617_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n2861), 
            .I3(n30391), .O(n2865[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_15 (.CI(n30391), .I0(encoder0_position[13]), .I1(n2861), 
            .CO(n30392));
    SB_LUT4 add_617_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n2861), 
            .I3(n30390), .O(n2865[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_14 (.CI(n30390), .I0(encoder0_position[12]), .I1(n2861), 
            .CO(n30391));
    SB_LUT4 add_617_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n2861), 
            .I3(n30389), .O(n2865[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_13 (.CI(n30389), .I0(encoder0_position[11]), .I1(n2861), 
            .CO(n30390));
    SB_LUT4 add_617_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n2861), 
            .I3(n30388), .O(n2865[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_12 (.CI(n30388), .I0(encoder0_position[10]), .I1(n2861), 
            .CO(n30389));
    SB_LUT4 add_617_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n2861), 
            .I3(n30387), .O(n2865[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_11 (.CI(n30387), .I0(encoder0_position[9]), .I1(n2861), 
            .CO(n30388));
    SB_LUT4 add_617_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n2861), 
            .I3(n30386), .O(n2865[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_10 (.CI(n30386), .I0(encoder0_position[8]), .I1(n2861), 
            .CO(n30387));
    SB_LUT4 add_617_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n2861), 
            .I3(n30385), .O(n2865[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_9 (.CI(n30385), .I0(encoder0_position[7]), .I1(n2861), 
            .CO(n30386));
    SB_LUT4 add_617_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n2861), 
            .I3(n30384), .O(n2865[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_8 (.CI(n30384), .I0(encoder0_position[6]), .I1(n2861), 
            .CO(n30385));
    SB_LUT4 add_617_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n2861), 
            .I3(n30383), .O(n2865[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_7 (.CI(n30383), .I0(encoder0_position[5]), .I1(n2861), 
            .CO(n30384));
    SB_LUT4 add_617_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n2861), 
            .I3(n30382), .O(n2865[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_6_lut.LUT_INIT = 16'hC33C;
    SB_DFF count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .D(n18802));   // quad.v(35[10] 41[6])
    SB_CARRY add_617_6 (.CI(n30382), .I0(encoder0_position[4]), .I1(n2861), 
            .CO(n30383));
    SB_LUT4 add_617_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n2861), 
            .I3(n30381), .O(n2865[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_5 (.CI(n30381), .I0(encoder0_position[3]), .I1(n2861), 
            .CO(n30382));
    SB_LUT4 add_617_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n2861), 
            .I3(n30380), .O(n2865[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_4 (.CI(n30380), .I0(encoder0_position[2]), .I1(n2861), 
            .CO(n30381));
    SB_LUT4 add_617_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n2861), 
            .I3(n30379), .O(n2865[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_3 (.CI(n30379), .I0(encoder0_position[1]), .I1(n2861), 
            .CO(n30380));
    SB_LUT4 add_617_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n30378), .O(n2865[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_617_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_617_2 (.CI(n30378), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n30379));
    SB_CARRY add_617_1 (.CI(GND_net), .I0(n2861), .I1(n2861), .CO(n30378));
    SB_LUT4 i892_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2861));   // quad.v(37[5] 40[8])
    defparam i892_1_lut_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    \grp_debouncer(2,5)_U0  debounce (.n19406(n19406), .data_o({data_o}), 
            .clk32MHz(clk32MHz), .reg_B({reg_B}), .PIN_2_c_0(PIN_2_c_0), 
            .n18805(n18805), .PIN_1_c_1(PIN_1_c_1), .GND_net(GND_net), 
            .n39036(n39036)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5)_U0 
//

module \grp_debouncer(2,5)_U0  (n19406, data_o, clk32MHz, reg_B, PIN_2_c_0, 
            n18805, PIN_1_c_1, GND_net, n39036) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n19406;
    output [1:0]data_o;
    input clk32MHz;
    output [1:0]reg_B;
    input PIN_2_c_0;
    input n18805;
    input PIN_1_c_1;
    input GND_net;
    output n39036;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    wire [2:0]n17;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire cnt_next_2__N_3559, n2;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n19406));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1150__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_2_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n18805));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1150__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1150__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_1_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n39036), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i24995_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i24995_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n39036));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i25004_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i25004_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i24997_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i24997_2_lut.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (n19395, encoder1_position, clk32MHz, 
            n19396, n19397, n19398, n19399, n19400, n19401, n19387, 
            n19388, n19389, n19390, n19391, n19392, n19393, n19394, 
            n19383, n19384, n19385, n19386, n19379, n19380, n19381, 
            n19382, data_o, GND_net, n2815, n18804, count_enable, 
            n19450, PIN_6_c_0, reg_B, PIN_7_c_1, n18830, n39886) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n19395;
    output [23:0]encoder1_position;
    input clk32MHz;
    input n19396;
    input n19397;
    input n19398;
    input n19399;
    input n19400;
    input n19401;
    input n19387;
    input n19388;
    input n19389;
    input n19390;
    input n19391;
    input n19392;
    input n19393;
    input n19394;
    input n19383;
    input n19384;
    input n19385;
    input n19386;
    input n19379;
    input n19380;
    input n19381;
    input n19382;
    output [1:0]data_o;
    input GND_net;
    output [23:0]n2815;
    input n18804;
    output count_enable;
    input n19450;
    input PIN_6_c_0;
    output [1:0]reg_B;
    input PIN_7_c_1;
    input n18830;
    output n39886;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire B_delayed, A_delayed, count_direction, n2808, n30547, n30546, 
        n30545, n30544, n30543, n30542, n30541, n30540, n30539, 
        n30538, n30537, n30536, n30535, n30534, n30533, n30532, 
        n30531, n30530, n30529, n30528, n30527, n30526, n30525, 
        n30524;
    
    SB_DFF count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .D(n19395));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .D(n19396));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .D(n19397));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .D(n19398));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .D(n19399));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .D(n19400));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .D(n19401));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .D(n19387));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .D(n19388));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .D(n19389));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .D(n19390));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .D(n19391));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .D(n19392));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .D(n19393));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .D(n19394));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .D(n19383));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .D(n19384));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .D(n19385));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .D(n19386));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .D(n19379));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .D(n19380));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .D(n19381));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .D(n19382));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_591_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2808), 
            .I3(n30547), .O(n2815[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_591_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2808), 
            .I3(n30546), .O(n2815[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_24 (.CI(n30546), .I0(encoder1_position[22]), .I1(n2808), 
            .CO(n30547));
    SB_LUT4 add_591_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2808), 
            .I3(n30545), .O(n2815[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_23 (.CI(n30545), .I0(encoder1_position[21]), .I1(n2808), 
            .CO(n30546));
    SB_LUT4 add_591_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2808), 
            .I3(n30544), .O(n2815[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_22 (.CI(n30544), .I0(encoder1_position[20]), .I1(n2808), 
            .CO(n30545));
    SB_LUT4 add_591_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2808), 
            .I3(n30543), .O(n2815[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_21 (.CI(n30543), .I0(encoder1_position[19]), .I1(n2808), 
            .CO(n30544));
    SB_LUT4 add_591_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2808), 
            .I3(n30542), .O(n2815[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_20 (.CI(n30542), .I0(encoder1_position[18]), .I1(n2808), 
            .CO(n30543));
    SB_LUT4 add_591_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2808), 
            .I3(n30541), .O(n2815[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_19 (.CI(n30541), .I0(encoder1_position[17]), .I1(n2808), 
            .CO(n30542));
    SB_LUT4 add_591_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2808), 
            .I3(n30540), .O(n2815[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_18 (.CI(n30540), .I0(encoder1_position[16]), .I1(n2808), 
            .CO(n30541));
    SB_LUT4 add_591_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2808), 
            .I3(n30539), .O(n2815[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_17 (.CI(n30539), .I0(encoder1_position[15]), .I1(n2808), 
            .CO(n30540));
    SB_LUT4 add_591_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2808), 
            .I3(n30538), .O(n2815[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_16 (.CI(n30538), .I0(encoder1_position[14]), .I1(n2808), 
            .CO(n30539));
    SB_LUT4 add_591_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2808), 
            .I3(n30537), .O(n2815[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_15 (.CI(n30537), .I0(encoder1_position[13]), .I1(n2808), 
            .CO(n30538));
    SB_LUT4 add_591_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2808), 
            .I3(n30536), .O(n2815[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_14 (.CI(n30536), .I0(encoder1_position[12]), .I1(n2808), 
            .CO(n30537));
    SB_LUT4 add_591_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2808), 
            .I3(n30535), .O(n2815[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_13 (.CI(n30535), .I0(encoder1_position[11]), .I1(n2808), 
            .CO(n30536));
    SB_LUT4 add_591_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2808), 
            .I3(n30534), .O(n2815[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_12 (.CI(n30534), .I0(encoder1_position[10]), .I1(n2808), 
            .CO(n30535));
    SB_LUT4 add_591_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2808), 
            .I3(n30533), .O(n2815[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_11 (.CI(n30533), .I0(encoder1_position[9]), .I1(n2808), 
            .CO(n30534));
    SB_LUT4 add_591_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2808), 
            .I3(n30532), .O(n2815[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_10 (.CI(n30532), .I0(encoder1_position[8]), .I1(n2808), 
            .CO(n30533));
    SB_LUT4 add_591_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2808), 
            .I3(n30531), .O(n2815[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_9 (.CI(n30531), .I0(encoder1_position[7]), .I1(n2808), 
            .CO(n30532));
    SB_LUT4 add_591_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2808), 
            .I3(n30530), .O(n2815[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_8 (.CI(n30530), .I0(encoder1_position[6]), .I1(n2808), 
            .CO(n30531));
    SB_LUT4 add_591_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2808), 
            .I3(n30529), .O(n2815[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_7 (.CI(n30529), .I0(encoder1_position[5]), .I1(n2808), 
            .CO(n30530));
    SB_LUT4 add_591_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2808), 
            .I3(n30528), .O(n2815[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_6 (.CI(n30528), .I0(encoder1_position[4]), .I1(n2808), 
            .CO(n30529));
    SB_LUT4 add_591_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2808), 
            .I3(n30527), .O(n2815[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_5 (.CI(n30527), .I0(encoder1_position[3]), .I1(n2808), 
            .CO(n30528));
    SB_LUT4 add_591_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2808), 
            .I3(n30526), .O(n2815[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_4 (.CI(n30526), .I0(encoder1_position[2]), .I1(n2808), 
            .CO(n30527));
    SB_LUT4 add_591_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2808), 
            .I3(n30525), .O(n2815[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_3 (.CI(n30525), .I0(encoder1_position[1]), .I1(n2808), 
            .CO(n30526));
    SB_LUT4 add_591_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n30524), .O(n2815[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_591_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_591_2 (.CI(n30524), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n30525));
    SB_DFF count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .D(n18804));   // quad.v(35[10] 41[6])
    SB_CARRY add_591_1 (.CI(GND_net), .I0(n2808), .I1(n2808), .CO(n30524));
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i891_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2808));   // quad.v(37[5] 40[8])
    defparam i891_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)  debounce (.n19450(n19450), .data_o({data_o}), .clk32MHz(clk32MHz), 
            .PIN_6_c_0(PIN_6_c_0), .reg_B({reg_B}), .PIN_7_c_1(PIN_7_c_1), 
            .n18830(n18830), .GND_net(GND_net), .n39886(n39886)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5) 
//

module \grp_debouncer(2,5)  (n19450, data_o, clk32MHz, PIN_6_c_0, reg_B, 
            PIN_7_c_1, n18830, GND_net, n39886) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n19450;
    output [1:0]data_o;
    input clk32MHz;
    input PIN_6_c_0;
    output [1:0]reg_B;
    input PIN_7_c_1;
    input n18830;
    input GND_net;
    output n39886;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n1;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    
    wire cnt_next_2__N_3559;
    wire [2:0]n17;
    
    wire n2;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n19450));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_6_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_7_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1151__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n1), .R(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n18830));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1151__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1151__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n39886), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3559));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i1434_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(170[42:59])
    defparam i1434_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[1]), .I2(cnt_reg[2]), 
            .I3(GND_net), .O(n39886));
    defparam i2_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i25026_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i25026_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i25019_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i25019_2_lut.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (\Kp[4] , \Kp[2] , GND_net, \Kp[3] , \Kp[0] , 
            \Kp[1] , \Kp[5] , duty, PWMLimit, \Ki[7] , IntegralLimit, 
            \Kp[6] , \Kp[7] , \Ki[1] , \Ki[0] , \Ki[2] , \Ki[3] , 
            \Ki[4] , \Ki[5] , \Ki[6] , clk32MHz, VCC_net, n25, motor_state, 
            setpoint, n45865) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input \Kp[4] ;
    input \Kp[2] ;
    input GND_net;
    input \Kp[3] ;
    input \Kp[0] ;
    input \Kp[1] ;
    input \Kp[5] ;
    output [23:0]duty;
    input [23:0]PWMLimit;
    input \Ki[7] ;
    input [23:0]IntegralLimit;
    input \Kp[6] ;
    input \Kp[7] ;
    input \Ki[1] ;
    input \Ki[0] ;
    input \Ki[2] ;
    input \Ki[3] ;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Ki[6] ;
    input clk32MHz;
    input VCC_net;
    input n25;
    input [23:0]motor_state;
    input [23:0]setpoint;
    output n45865;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n30357;
    wire [23:0]n2942;
    wire [23:0]n2967;
    
    wire n30358;
    wire [3:0]n9076;
    
    wire n6;
    wire [23:0]\PID_CONTROLLER.err ;   // verilog/motorControl.v(29[23:26])
    
    wire n8, n11, n32197;
    wire [14:0]n9241;
    
    wire n460, n32198;
    wire [23:0]duty_23__N_3478;
    
    wire n30356, n31958;
    wire [14:0]n8944;
    
    wire n31959;
    wire [15:0]n9223;
    
    wire n387, n32196;
    wire [15:0]n8926;
    
    wire n31957;
    wire [2:0]n9082;
    
    wire n4, n6_adj_3567, n314, n32195, n30099, n12, n18, n13, 
        n47;
    wire [23:0]n1;
    
    wire n30500, n4_adj_3568, n39599, n241, n32194, n31956;
    wire [23:0]n257;
    
    wire n30499, n533, n31955, n460_adj_3569, n31954, n168, n32193, 
        n387_adj_3570, n31953, n314_adj_3571, n31952, n30355, n26, 
        n95, n241_adj_3572, n31951, n30498, n30497, n30496, n168_adj_3575, 
        n31950;
    wire [16:0]n9204;
    
    wire n32192, n32191, n26_adj_3576, n95_adj_3577, n32190;
    wire [16:0]n8907;
    
    wire n31949, n31948, n32189, n31947, n32188, n32187, n31946, 
        n31945, duty_23__N_3502;
    wire [23:0]duty_23__N_3355;
    
    wire n32186, n31944, n32185, n30495, n30494;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(31[23:31])
    
    wire n524, n232, n305, n31943, n378, n32184;
    wire [23:0]n1_adj_3897;
    
    wire n30493, n451, n524_adj_3579, n89, n20_adj_3581, n162, n80, 
        n235, n308, n381, n89_adj_3582, n11_adj_3583, n20_adj_3584, 
        n341, n162_adj_3585, n454, n414, n235_adj_3586, n527, n308_adj_3587, 
        n381_adj_3588, n454_adj_3589, n527_adj_3591, n77, n153, n8_adj_3592, 
        n150, n223, n296, n226, n30492, n32183, n31942, n530, 
        n32182, n31941, n31940, n457, n32181, n299, n530_adj_3594, 
        n31939, n457_adj_3595, n31938;
    wire [23:0]\PID_CONTROLLER.err_23__N_3379 ;
    
    wire n384, n32180, n92, n384_adj_3596, n31937, n311, n31936, 
        n30491, n311_adj_3598, n32179, n238, n31935, n23, n165, 
        n238_adj_3600, n165_adj_3602, n31934, n23_adj_3603, n92_adj_3604, 
        n30490, n32178, n30489, n32177;
    wire [17:0]n8887;
    
    wire n31933, n31932, n31931;
    wire [17:0]n9184;
    
    wire n32176, n31930, n32175, n32174, n30488, n31929, n32173, 
        n31928, n32172, n32171, n31927, n32170, n30487, n31926, 
        n30486, n31925, n32169, n31924, n32168, n31923, n30485, 
        n31922, n30484, n31921, n32167, n31920, n372, n32166, 
        n31919, n32165, n31918, n32164, n31917, n32163;
    wire [18:0]n8866;
    
    wire n31916, n31915, n32162, n31914, n31913, n32161, n31912, 
        n32160, n445, n31911;
    wire [18:0]n9163;
    
    wire n32159, n32158, n31910, n32157, n31909, n30483, n31908, 
        n32156, n31907, n30482, n32155, n31906, n32154, n31905, 
        n518, n32153, n41, n31904, n39, n31903, n45, n32152, 
        n43, n37, n29, n31, n23_adj_3606, n25_c, n32151, n31902, 
        n30481, n31901, n32150, n35, n11_adj_3607, n13_adj_3608, 
        n32149, n32148, n31900, n32147, n451_adj_3610, n32146, n15_adj_3611, 
        n159, n31899, n27, n33, n17_adj_3612, n86, n30480, n9_adj_3613, 
        n378_adj_3614, n32145;
    wire [19:0]n8844;
    
    wire n31898, n31897, n17_adj_3615, n19_adj_3616, n31896, n21_adj_3618, 
        n31895, n305_adj_3619, n32144, n31894, n43517, n43469, n12_adj_3620, 
        n30, n43545, n44153, n31893, n44143, n31892, n44916, n44457, 
        n45016, n232_adj_3621, n32143, n6_adj_3622, n44674, n31891, 
        n159_adj_3623, n32142, n44675, n487, n16_adj_3624, n24, 
        n43392, n30479, n31890, n17_adj_3626, n86_adj_3627, n8_adj_3628, 
        n43388, n44611;
    wire [19:0]n9141;
    
    wire n32141, n31889, n43886, n31888, n32140, n4_adj_3629, n44669, 
        n44670, n43421, n10_adj_3630, n43416, n44958, n43888, n31887, 
        n30478, n32139, n31886, n32138, n45090, n45091, n45060, 
        n256, n26500, n32137, n521, n31885, n43394, n44830, n448, 
        n31884, n43894, n375, n31883, n42863, n44992, n32136;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3454 ;
    
    wire n30477, n80_adj_3635, n302, n31882, n32135, n229, n31881, 
        n32134, n45_adj_3636, n30476, n11_adj_3638, n156, n31880, 
        n153_adj_3639, n32133, n14_adj_3640, n83, n32132;
    wire [20:0]n8821;
    
    wire n31879, n31878, n43_adj_3641, n30475, n41_adj_3643, n30474, 
        n39_adj_3645, n30473, n37_adj_3647, n30472, n226_adj_3649, 
        n35_adj_3650, n30471, n31877, n32131, n33_adj_3652, n30470, 
        n299_adj_3654, n31_adj_3655, n30469, n372_adj_3657, n445_adj_3658, 
        n32130, n29_adj_3659, n30468, n31876, n32129, n31875, n369, 
        n27_adj_3661, n30467, n521_adj_3663, n32128, n31874, n31873, 
        n448_adj_3664, n32127, n375_adj_3665, n32126, n31872, n25_adj_3666, 
        n30466, n31871, n302_adj_3668, n32125, n31870, n229_adj_3669, 
        n32124, n31869, n31868, n156_adj_3670, n32123, n31867, n23_adj_3671, 
        n30465, n31866, n14_adj_3673, n83_adj_3674;
    wire [20:0]n9118;
    
    wire n32122, n32121, n32120, n518_adj_3675, n31865, n32119, 
        n32118, n31864, n32117, n31863, n32116, n31862, n32115, 
        n32114, n31861, n31860;
    wire [0:0]n7831;
    wire [21:0]n8797;
    
    wire n31859, n31858, n32113, n32112, n32111, n21_adj_3676, n30464, 
        n19_adj_3677, n30463, n32110, n31857, n31856, n32109, n31855, 
        n31854, n32108, n31853, n32107, n32106, n31852, n17_adj_3678, 
        n30462, n32105, n31851, n31850, n15_adj_3679, n30461, n32104, 
        n32103, n31849, n31848, n31847, n31846, n42910;
    wire [21:0]n9094;
    
    wire n32102, n31845, n13_adj_3680, n30460;
    wire [47:0]n155;
    wire [23:0]n34;
    
    wire \PID_CONTROLLER.integral_23__N_3451 , n11_adj_3681, n30459, n32101, 
        n31844, n32100, n560, n32099, n512, n31843, n9_adj_3683, 
        n30458, n442, n125_adj_3685, n56, n515, n198, n439, n31842, 
        n271_adj_3686, n32098, n32097, n366, n31841, n32096, n293, 
        n31840, n32095, n7_adj_3687, n30457, n32094, n220, n31839, 
        n147, n31838, n5_adj_3689, n74, n32093, n31837, n31836, 
        n32092, n32091, n31835, n32090, n32089, n31834, n32088, 
        n32087, n31833, n512_adj_3690, n32086, n31832, n439_adj_3691, 
        n32085, n31831, n31830, n366_adj_3693, n32084, n31829, n293_adj_3694, 
        n32083, n31828, n31827, n220_adj_3695, n32082, n147_adj_3696, 
        n32081, n31826, n5_adj_3697, n74_adj_3698, n5_adj_3699, n30456, 
        n41_adj_3701, n39_adj_3702, n45_adj_3703, n27_adj_3704, n29_adj_3705, 
        n31_adj_3706, n33_adj_3707, n35_adj_3708, n37_adj_3709, n43_adj_3710, 
        n15_adj_3711, n17_adj_3712, n19_adj_3713, n21_adj_3714, n23_adj_3715, 
        n25_adj_3716, n9_adj_3717, n43329, n13_adj_3718, n11_adj_3719, 
        n43317, n12_adj_3720, n10_adj_3721, n30_adj_3722, n43386, 
        n44061, n44053, n44896, n44423, n45012, n16_adj_3723, n6_adj_3724, 
        n44651, n44652, n8_adj_3725, n24_adj_3726, n43267, n43263, 
        n44613, n43896, n4_adj_3727, n44641, n44642, n43303, n43293, 
        n44962, n43898, n45092, n45093, n45058, n43271, n44832, 
        n43904, n44994, n31825, n32080, n32079, n31824, n32078, 
        n31823, n32077, n515_adj_3729, n31822, n32076, n442_adj_3730, 
        n31821, n32075, n369_adj_3731, n31820, n32074, n296_adj_3732, 
        n31819, n223_adj_3733, n31818, n32073, n150_adj_3734, n31817, 
        n32072, n8_adj_3735, n77_adj_3736, n32071;
    wire [5:0]n9358;
    
    wire n38956, n490, n32302, n32070;
    wire [4:0]n9366;
    
    wire n417, n32301, n32069, n344, n32300, n32068, n3_adj_3737, 
        n30455, n32299, n32067, n32066, n32298, n32065, n32064;
    wire [6:0]n9349;
    
    wire n32297, n32063, n32296, n32062, n32061, n32060, n32295, 
        n32294;
    wire [5:0]n9061;
    
    wire n490_adj_3739, n32059, n268_adj_3740, n32293, n195_adj_3741, 
        n32292;
    wire [4:0]n9069;
    
    wire n417_adj_3742, n32058, n53, n122, n344_adj_3743, n32057, 
        n271_adj_3744, n32056;
    wire [7:0]n9339;
    
    wire n32291, n557, n32290, n198_adj_3745, n32055, n484, n32289, 
        n56_adj_3746, n125_adj_3747, n411, n32288;
    wire [6:0]n9052;
    
    wire n560_adj_3748, n32054, n338, n32287, n487_adj_3749, n32053, 
        n265_adj_3750, n32286, n414_adj_3751, n32052, n341_adj_3752, 
        n32051, n192_adj_3753, n32285, n268_adj_3754, n32050, n195_adj_3755, 
        n32049, n50, n119, n53_adj_3756, n122_adj_3757;
    wire [8:0]n9328;
    
    wire n32284, n32283, n4_adj_3758;
    wire [3:0]n9373;
    
    wire n6_adj_3759, n30129, n554, n32282, n481, n32281;
    wire [7:0]n9042;
    
    wire n32048, n557_adj_3760, n32047, n484_adj_3761, n32046, n411_adj_3762, 
        n32045, n30206;
    wire [1:0]n9384;
    
    wire n4_adj_3763;
    wire [2:0]n9379;
    
    wire n62, n131, n204, n4_adj_3764, n408, n32280, n338_adj_3765, 
        n32044, n335, n32279, n265_adj_3766, n32043, n262_adj_3767, 
        n32278, n192_adj_3768, n32042, n189_adj_3769, n32277, n50_adj_3770, 
        n119_adj_3771, n47_adj_3772, n116;
    wire [8:0]n9031;
    
    wire n32041;
    wire [9:0]n9316;
    
    wire n32276, n32040, n32275, n554_adj_3773, n32039, n32274, 
        n481_adj_3774, n32038;
    wire [23:0]n1_adj_3898;
    
    wire n30523, n551, n32273, n408_adj_3776, n32037, n335_adj_3777, 
        n32036, n478, n32272, n262_adj_3778, n32035, n189_adj_3779, 
        n32034, n405, n32271, n332, n32270, n259_adj_3780, n32269, 
        n30522, n47_adj_3782, n116_adj_3783, n186_adj_3784, n32268;
    wire [9:0]n9019;
    
    wire n32033, n44, n113, n32032, n30521;
    wire [10:0]n9303;
    
    wire n32267, n32031, n32266, n32265, n551_adj_3790, n32030, 
        n32264, n548, n32263, n478_adj_3791, n32029, n475, n32262, 
        n405_adj_3792, n32028, n332_adj_3793, n32027, n402, n32261, 
        n259_adj_3794, n32026, n329, n32260, n186_adj_3795, n32025, 
        n256_adj_3796, n32259, n44_adj_3797, n113_adj_3798;
    wire [10:0]n9006;
    
    wire n32024, n32023, n32022, n32021, n183_adj_3799, n32258, 
        n548_adj_3800, n32020, n41_adj_3801, n110_adj_3802, n475_adj_3803, 
        n32019, n31207, n31206;
    wire [11:0]n9289;
    
    wire n32257, n402_adj_3804, n32018, n32256, n32255, n329_adj_3805, 
        n32017, n31205, n32254, n256_adj_3806, n32016, n31204, n30520, 
        n31203, n32253, n183_adj_3808, n32015, n41_adj_3809, n110_adj_3810, 
        n545, n32252, n31202;
    wire [11:0]n8992;
    
    wire n32014, n31201, n30519, n472, n32251, n32013, n399, n32250, 
        n32012, n31200, n31199, n31198, n32011, n326, n32249, 
        n31197, n253, n32248, n32010, n31196, n31195, n30518, 
        n180, n32247, n30377, n30376, n545_adj_3813, n32009, n38, 
        n107_adj_3814;
    wire [12:0]n9274;
    
    wire n32246, n472_adj_3815, n32008, n399_adj_3816, n32007, n31194, 
        n326_adj_3817, n32006, n31193, n32245, n253_adj_3818, n32005, 
        n31192, n32244, n180_adj_3819, n32004, n31191, n38_adj_3820, 
        n107_adj_3821, n31190, n32243;
    wire [12:0]n8977;
    
    wire n32003, n30375, n30517, n31189, n32242, n32002, n32001, 
        n31188, n32241, n30516, n31187, n30515, n542, n32240, 
        n32000, n31186, n31185, n30374, n30514, n30373, n30372, 
        n31999, n469, n32239, n31998, n396, n32238, n542_adj_3826, 
        n31997, n323, n32237, n469_adj_3827, n31996, n250, n32236, 
        n396_adj_3828, n31995, n177, n32235, n323_adj_3829, n31994, 
        n30513, n35_adj_3831, n104_adj_3832, n250_adj_3833, n31993;
    wire [13:0]n9258;
    
    wire n32234, n177_adj_3834, n31992, n32233, n35_adj_3835, n104_adj_3836, 
        n32232;
    wire [13:0]n8961;
    
    wire n31991, n31990, n32231, n31989, n32230, n31988, n32229, 
        n31987, n12_adj_3837, n31986, n32228, n31985, n8_adj_3838, 
        n30371, n539, n32227, n539_adj_3839, n31984, n11_adj_3840, 
        n6_adj_3841, n466, n32226, n466_adj_3842, n31983, n393, 
        n31982, n30512, n30231, n30511, n18_adj_3845, n13_adj_3846, 
        n393_adj_3847, n32225, n30510, n320, n31981, n30370, n320_adj_3849, 
        n32224, n247, n31980, n30509, n30369, n174, n31979, n247_adj_3851, 
        n32223, n30368, n30508, n32, n101, n174_adj_3853, n32222, 
        n31978, n32_adj_3854, n101_adj_3855, n31977, n32221, n32220, 
        n32219, n32218, n31976, n32217, n30367, n30507, n32216, 
        n32215, n30366, n31975, n30506, n30505, n31974, n32214, 
        n31973, n31972, n536, n32213, n463, n32212, n390, n32211, 
        n317, n32210, n244, n32209, n31971, n536_adj_3859, n31970, 
        n30365, n171, n32208, n463_adj_3860, n31969, n29_adj_3861, 
        n98, n30504, n390_adj_3863, n31968, n30364, n32207, n30363, 
        n32206, n32205, n317_adj_3864, n31967, n32204, n30362, n32203, 
        n32202, n244_adj_3865, n31966, n171_adj_3866, n31965, n29_adj_3867, 
        n98_adj_3868, n32201, n31964, n31963, n30361, n30503, n30360, 
        n32200, n31962, n30359, n30502, n32199, n31961, n533_adj_3871, 
        n31960, n30501, n17_adj_3874, n9_adj_3875, n11_adj_3876, n43376, 
        n43337, n46698, n44381, n43915, n46680, n43829, n43819, 
        n46673, n43593, n43618, n16_adj_3877, n43547, n8_adj_3878, 
        n24_adj_3879, n43656, n44253, n44247, n44932, n44509, n45018, 
        n43919, n46667, n43745, n46661, n12_adj_3880, n43703, n46685, 
        n10_adj_3881, n30_adj_3882, n44577, n43086, n46665, n44319, 
        n46691, n44778, n46656, n45022, n46653, n16_adj_3883, n43660, 
        n24_adj_3884, n6_adj_3885, n44720, n44721, n43666, n8_adj_3886, 
        n46651, n44607, n44604, n4_adj_3887, n44712, n44713, n12_adj_3888, 
        n43568, n10_adj_3889, n30_adj_3890, n43571, n44948, n43878, 
        n45082, n45083, n45069, n6_adj_3891, n44714, n44715, n43550, 
        n44609, n43876, n43554, n44988, n43884, n44990, n4_adj_3892, 
        n44718, n44719, n43708, n44946, n28, n45078, n45079, n45073, 
        n43668, n44984, n43874, \PID_CONTROLLER.integral_23__N_3453 , 
        n44986, n4_adj_3893, n29997, n204_adj_3894;
    wire [1:0]n9087;
    
    wire n30074, n131_adj_3895, n62_adj_3896;
    
    SB_CARRY add_628_5 (.CI(n30357), .I0(n2942[3]), .I1(n2967[3]), .CO(n30358));
    SB_LUT4 i25076_4_lut (.I0(n9076[2]), .I1(\Kp[4] ), .I2(n6), .I3(\PID_CONTROLLER.err [18]), 
            .O(n8));   // verilog/motorControl.v(42[17:23])
    defparam i25076_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(\PID_CONTROLLER.err [19]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n11));   // verilog/motorControl.v(42[17:23])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_CARRY add_4608_7 (.CI(n32197), .I0(n9241[4]), .I1(n460), .CO(n32198));
    SB_LUT4 add_628_4_lut (.I0(GND_net), .I1(n2942[2]), .I2(n2967[2]), 
            .I3(n30356), .O(duty_23__N_3478[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4586_11 (.CI(n31958), .I0(n8944[8]), .I1(GND_net), .CO(n31959));
    SB_LUT4 add_4608_6_lut (.I0(GND_net), .I1(n9241[3]), .I2(n387), .I3(n32196), 
            .O(n9223[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4586_10_lut (.I0(GND_net), .I1(n8944[7]), .I2(GND_net), 
            .I3(n31957), .O(n8926[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25107_4_lut (.I0(n9082[1]), .I1(\Kp[3] ), .I2(n4), .I3(\PID_CONTROLLER.err [19]), 
            .O(n6_adj_3567));   // verilog/motorControl.v(42[17:23])
    defparam i25107_4_lut.LUT_INIT = 16'he8a0;
    SB_CARRY add_4608_6 (.CI(n32196), .I0(n9241[3]), .I1(n387), .CO(n32197));
    SB_LUT4 add_4608_5_lut (.I0(GND_net), .I1(n9241[2]), .I2(n314), .I3(n32195), 
            .O(n9223[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4608_5 (.CI(n32195), .I0(n9241[2]), .I1(n314), .CO(n32196));
    SB_CARRY add_4586_10 (.CI(n31957), .I0(n8944[7]), .I1(GND_net), .CO(n31958));
    SB_LUT4 i25142_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n30099));   // verilog/motorControl.v(42[17:23])
    defparam i25142_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut (.I0(n6_adj_3567), .I1(n11), .I2(n8), .I3(n12), 
            .O(n18));   // verilog/motorControl.v(42[17:23])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [18]), 
            .I3(\PID_CONTROLLER.err [22]), .O(n13));   // verilog/motorControl.v(42[17:23])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(duty[23]), .I1(GND_net), .I2(n1[23]), 
            .I3(n30500), .O(n47)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n13), .I1(n18), .I2(n30099), .I3(n4_adj_3568), 
            .O(n39599));   // verilog/motorControl.v(42[17:23])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4608_4_lut (.I0(GND_net), .I1(n9241[1]), .I2(n241), .I3(n32194), 
            .O(n9223[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4586_9_lut (.I0(GND_net), .I1(n8944[6]), .I2(GND_net), 
            .I3(n31956), .O(n8926[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4586_9 (.CI(n31956), .I0(n8944[6]), .I1(GND_net), .CO(n31957));
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1[22]), 
            .I3(n30499), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4586_8_lut (.I0(GND_net), .I1(n8944[5]), .I2(n533), .I3(n31955), 
            .O(n8926[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4608_4 (.CI(n32194), .I0(n9241[1]), .I1(n241), .CO(n32195));
    SB_CARRY add_4586_8 (.CI(n31955), .I0(n8944[5]), .I1(n533), .CO(n31956));
    SB_LUT4 add_4586_7_lut (.I0(GND_net), .I1(n8944[4]), .I2(n460_adj_3569), 
            .I3(n31954), .O(n8926[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4586_7 (.CI(n31954), .I0(n8944[4]), .I1(n460_adj_3569), 
            .CO(n31955));
    SB_LUT4 add_4608_3_lut (.I0(GND_net), .I1(n9241[0]), .I2(n168), .I3(n32193), 
            .O(n9223[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4586_6_lut (.I0(GND_net), .I1(n8944[3]), .I2(n387_adj_3570), 
            .I3(n31953), .O(n8926[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4586_6 (.CI(n31953), .I0(n8944[3]), .I1(n387_adj_3570), 
            .CO(n31954));
    SB_CARRY unary_minus_16_add_3_24 (.CI(n30499), .I0(GND_net), .I1(n1[22]), 
            .CO(n30500));
    SB_CARRY add_628_4 (.CI(n30356), .I0(n2942[2]), .I1(n2967[2]), .CO(n30357));
    SB_CARRY add_4608_3 (.CI(n32193), .I0(n9241[0]), .I1(n168), .CO(n32194));
    SB_LUT4 add_4586_5_lut (.I0(GND_net), .I1(n8944[2]), .I2(n314_adj_3571), 
            .I3(n31952), .O(n8926[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_628_3_lut (.I0(GND_net), .I1(n2942[1]), .I2(n2967[1]), 
            .I3(n30355), .O(duty_23__N_3478[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4608_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n9223[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4586_5 (.CI(n31952), .I0(n8944[2]), .I1(n314_adj_3571), 
            .CO(n31953));
    SB_LUT4 add_4586_4_lut (.I0(GND_net), .I1(n8944[1]), .I2(n241_adj_3572), 
            .I3(n31951), .O(n8926[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_3 (.CI(n30355), .I0(n2942[1]), .I1(n2967[1]), .CO(n30356));
    SB_LUT4 add_628_2_lut (.I0(GND_net), .I1(n2942[0]), .I2(n2967[0]), 
            .I3(GND_net), .O(duty_23__N_3478[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1[21]), 
            .I3(n30498), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n30498), .I0(GND_net), .I1(n1[21]), 
            .CO(n30499));
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1[20]), 
            .I3(n30497), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_22 (.CI(n30497), .I0(GND_net), .I1(n1[20]), 
            .CO(n30498));
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1[19]), 
            .I3(n30496), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4608_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n32193));
    SB_CARRY add_4586_4 (.CI(n31951), .I0(n8944[1]), .I1(n241_adj_3572), 
            .CO(n31952));
    SB_LUT4 add_4586_3_lut (.I0(GND_net), .I1(n8944[0]), .I2(n168_adj_3575), 
            .I3(n31950), .O(n8926[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4607_18_lut (.I0(GND_net), .I1(n9223[15]), .I2(GND_net), 
            .I3(n32192), .O(n9204[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4607_17_lut (.I0(GND_net), .I1(n9223[14]), .I2(GND_net), 
            .I3(n32191), .O(n9204[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4586_3 (.CI(n31950), .I0(n8944[0]), .I1(n168_adj_3575), 
            .CO(n31951));
    SB_CARRY add_4607_17 (.CI(n32191), .I0(n9223[14]), .I1(GND_net), .CO(n32192));
    SB_LUT4 add_4586_2_lut (.I0(GND_net), .I1(n26_adj_3576), .I2(n95_adj_3577), 
            .I3(GND_net), .O(n8926[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4586_2 (.CI(GND_net), .I0(n26_adj_3576), .I1(n95_adj_3577), 
            .CO(n31950));
    SB_LUT4 add_4607_16_lut (.I0(GND_net), .I1(n9223[13]), .I2(GND_net), 
            .I3(n32190), .O(n9204[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4585_18_lut (.I0(GND_net), .I1(n8926[15]), .I2(GND_net), 
            .I3(n31949), .O(n8907[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4585_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4607_16 (.CI(n32190), .I0(n9223[13]), .I1(GND_net), .CO(n32191));
    SB_LUT4 add_4585_17_lut (.I0(GND_net), .I1(n8926[14]), .I2(GND_net), 
            .I3(n31948), .O(n8907[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4585_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4607_15_lut (.I0(GND_net), .I1(n9223[12]), .I2(GND_net), 
            .I3(n32189), .O(n9204[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4585_17 (.CI(n31948), .I0(n8926[14]), .I1(GND_net), .CO(n31949));
    SB_CARRY add_4607_15 (.CI(n32189), .I0(n9223[12]), .I1(GND_net), .CO(n32190));
    SB_LUT4 add_4585_16_lut (.I0(GND_net), .I1(n8926[13]), .I2(GND_net), 
            .I3(n31947), .O(n8907[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4585_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4607_14_lut (.I0(GND_net), .I1(n9223[11]), .I2(GND_net), 
            .I3(n32188), .O(n9204[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4585_16 (.CI(n31947), .I0(n8926[13]), .I1(GND_net), .CO(n31948));
    SB_CARRY unary_minus_16_add_3_21 (.CI(n30496), .I0(GND_net), .I1(n1[19]), 
            .CO(n30497));
    SB_CARRY add_4607_14 (.CI(n32188), .I0(n9223[11]), .I1(GND_net), .CO(n32189));
    SB_LUT4 add_4607_13_lut (.I0(GND_net), .I1(n9223[10]), .I2(GND_net), 
            .I3(n32187), .O(n9204[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4585_15_lut (.I0(GND_net), .I1(n8926[12]), .I2(GND_net), 
            .I3(n31946), .O(n8907[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4585_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4585_15 (.CI(n31946), .I0(n8926[12]), .I1(GND_net), .CO(n31947));
    SB_CARRY add_4607_13 (.CI(n32187), .I0(n9223[10]), .I1(GND_net), .CO(n32188));
    SB_LUT4 add_4585_14_lut (.I0(GND_net), .I1(n8926[11]), .I2(GND_net), 
            .I3(n31945), .O(n8907[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4585_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4585_14 (.CI(n31945), .I0(n8926[11]), .I1(GND_net), .CO(n31946));
    SB_LUT4 duty_23__I_0_29_i2_3_lut (.I0(duty_23__N_3478[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[1]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4607_12_lut (.I0(GND_net), .I1(n9223[9]), .I2(GND_net), 
            .I3(n32186), .O(n9204[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4585_13_lut (.I0(GND_net), .I1(n8926[10]), .I2(GND_net), 
            .I3(n31944), .O(n8907[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4585_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_2 (.CI(GND_net), .I0(n2942[0]), .I1(n2967[0]), .CO(n30355));
    SB_CARRY add_4607_12 (.CI(n32186), .I0(n9223[9]), .I1(GND_net), .CO(n32187));
    SB_CARRY add_4585_13 (.CI(n31944), .I0(n8926[10]), .I1(GND_net), .CO(n31945));
    SB_LUT4 add_4607_11_lut (.I0(GND_net), .I1(n9223[8]), .I2(GND_net), 
            .I3(n32185), .O(n9204[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1[18]), 
            .I3(n30495), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_20 (.CI(n30495), .I0(GND_net), .I1(n1[18]), 
            .CO(n30496));
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1[17]), 
            .I3(n30494), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4585_12_lut (.I0(GND_net), .I1(n8926[9]), .I2(GND_net), 
            .I3(n31943), .O(n8907[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4585_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_19 (.CI(n30494), .I0(GND_net), .I1(n1[17]), 
            .CO(n30495));
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4607_11 (.CI(n32185), .I0(n9223[8]), .I1(GND_net), .CO(n32186));
    SB_LUT4 add_4607_10_lut (.I0(GND_net), .I1(n9223[7]), .I2(GND_net), 
            .I3(n32184), .O(n9204[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[6]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1[16]), 
            .I3(n30493), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_3579));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3581));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_3582));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3583));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3584));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_3585));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_3586));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_3587));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_3588));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_3589));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_3591));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3592));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4607_10 (.CI(n32184), .I0(n9223[7]), .I1(GND_net), .CO(n32185));
    SB_CARRY add_4585_12 (.CI(n31943), .I0(n8926[9]), .I1(GND_net), .CO(n31944));
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[7]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_16_add_3_18 (.CI(n30493), .I0(GND_net), .I1(n1[16]), 
            .CO(n30494));
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1[15]), 
            .I3(n30492), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4607_9_lut (.I0(GND_net), .I1(n9223[6]), .I2(GND_net), 
            .I3(n32183), .O(n9204[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4585_11_lut (.I0(GND_net), .I1(n8926[8]), .I2(GND_net), 
            .I3(n31942), .O(n8907[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4585_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4607_9 (.CI(n32183), .I0(n9223[6]), .I1(GND_net), .CO(n32184));
    SB_CARRY add_4585_11 (.CI(n31942), .I0(n8926[8]), .I1(GND_net), .CO(n31943));
    SB_LUT4 add_4607_8_lut (.I0(GND_net), .I1(n9223[5]), .I2(n530), .I3(n32182), 
            .O(n9204[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4585_10_lut (.I0(GND_net), .I1(n8926[7]), .I2(GND_net), 
            .I3(n31941), .O(n8907[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4585_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4585_10 (.CI(n31941), .I0(n8926[7]), .I1(GND_net), .CO(n31942));
    SB_CARRY add_4607_8 (.CI(n32182), .I0(n9223[5]), .I1(n530), .CO(n32183));
    SB_LUT4 add_4585_9_lut (.I0(GND_net), .I1(n8926[6]), .I2(GND_net), 
            .I3(n31940), .O(n8907[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4585_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4607_7_lut (.I0(GND_net), .I1(n9223[4]), .I2(n457), .I3(n32181), 
            .O(n9204[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4585_9 (.CI(n31940), .I0(n8926[6]), .I1(GND_net), .CO(n31941));
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4585_8_lut (.I0(GND_net), .I1(n8926[5]), .I2(n530_adj_3594), 
            .I3(n31939), .O(n8907[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4585_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4585_8 (.CI(n31939), .I0(n8926[5]), .I1(n530_adj_3594), 
            .CO(n31940));
    SB_LUT4 add_4585_7_lut (.I0(GND_net), .I1(n8926[4]), .I2(n457_adj_3595), 
            .I3(n31938), .O(n8907[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4585_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3355[0]));   // verilog/motorControl.v(37[14] 56[8])
    SB_CARRY add_4607_7 (.CI(n32181), .I0(n9223[4]), .I1(n457), .CO(n32182));
    SB_DFF \PID_CONTROLLER.err_i0  (.Q(\PID_CONTROLLER.err [0]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [0]));   // verilog/motorControl.v(37[14] 56[8])
    SB_LUT4 add_4607_6_lut (.I0(GND_net), .I1(n9223[3]), .I2(n384), .I3(n32180), 
            .O(n9204[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4585_7 (.CI(n31938), .I0(n8926[4]), .I1(n457_adj_3595), 
            .CO(n31939));
    SB_LUT4 add_4585_6_lut (.I0(GND_net), .I1(n8926[3]), .I2(n384_adj_3596), 
            .I3(n31937), .O(n8907[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4585_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4585_6 (.CI(n31937), .I0(n8926[3]), .I1(n384_adj_3596), 
            .CO(n31938));
    SB_CARRY add_4607_6 (.CI(n32180), .I0(n9223[3]), .I1(n384), .CO(n32181));
    SB_LUT4 add_4585_5_lut (.I0(GND_net), .I1(n8926[2]), .I2(n311), .I3(n31936), 
            .O(n8907[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4585_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_17 (.CI(n30492), .I0(GND_net), .I1(n1[15]), 
            .CO(n30493));
    SB_CARRY add_4585_5 (.CI(n31936), .I0(n8926[2]), .I1(n311), .CO(n31937));
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1[14]), 
            .I3(n30491), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4607_5_lut (.I0(GND_net), .I1(n9223[2]), .I2(n311_adj_3598), 
            .I3(n32179), .O(n9204[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4585_4_lut (.I0(GND_net), .I1(n8926[1]), .I2(n238), .I3(n31935), 
            .O(n8907[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4585_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4585_4 (.CI(n31935), .I0(n8926[1]), .I1(n238), .CO(n31936));
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_3600));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4607_5 (.CI(n32179), .I0(n9223[2]), .I1(n311_adj_3598), 
            .CO(n32180));
    SB_LUT4 add_4585_3_lut (.I0(GND_net), .I1(n8926[0]), .I2(n165_adj_3602), 
            .I3(n31934), .O(n8907[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4585_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4585_3 (.CI(n31934), .I0(n8926[0]), .I1(n165_adj_3602), 
            .CO(n31935));
    SB_CARRY unary_minus_16_add_3_16 (.CI(n30491), .I0(GND_net), .I1(n1[14]), 
            .CO(n30492));
    SB_LUT4 add_4585_2_lut (.I0(GND_net), .I1(n23_adj_3603), .I2(n92_adj_3604), 
            .I3(GND_net), .O(n8907[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4585_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_3604));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1[13]), 
            .I3(n30490), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3603));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4585_2 (.CI(GND_net), .I0(n23_adj_3603), .I1(n92_adj_3604), 
            .CO(n31934));
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_3602));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n30490), .I0(GND_net), .I1(n1[13]), 
            .CO(n30491));
    SB_LUT4 add_4607_4_lut (.I0(GND_net), .I1(n9223[1]), .I2(n238_adj_3600), 
            .I3(n32178), .O(n9204[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1[12]), 
            .I3(n30489), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4607_4 (.CI(n32178), .I0(n9223[1]), .I1(n238_adj_3600), 
            .CO(n32179));
    SB_LUT4 add_4607_3_lut (.I0(GND_net), .I1(n9223[0]), .I2(n165), .I3(n32177), 
            .O(n9204[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4607_3 (.CI(n32177), .I0(n9223[0]), .I1(n165), .CO(n32178));
    SB_LUT4 add_4584_19_lut (.I0(GND_net), .I1(n8907[16]), .I2(GND_net), 
            .I3(n31933), .O(n8887[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4584_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4584_18_lut (.I0(GND_net), .I1(n8907[15]), .I2(GND_net), 
            .I3(n31932), .O(n8887[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4584_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4584_18 (.CI(n31932), .I0(n8907[15]), .I1(GND_net), .CO(n31933));
    SB_LUT4 add_4584_17_lut (.I0(GND_net), .I1(n8907[14]), .I2(GND_net), 
            .I3(n31931), .O(n8887[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4584_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4607_2_lut (.I0(GND_net), .I1(n23), .I2(n92), .I3(GND_net), 
            .O(n9204[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4607_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4607_2 (.CI(GND_net), .I0(n23), .I1(n92), .CO(n32177));
    SB_CARRY add_4584_17 (.CI(n31931), .I0(n8907[14]), .I1(GND_net), .CO(n31932));
    SB_LUT4 add_4606_19_lut (.I0(GND_net), .I1(n9204[16]), .I2(GND_net), 
            .I3(n32176), .O(n9184[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4584_16_lut (.I0(GND_net), .I1(n8907[13]), .I2(GND_net), 
            .I3(n31930), .O(n8887[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4584_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4584_16 (.CI(n31930), .I0(n8907[13]), .I1(GND_net), .CO(n31931));
    SB_LUT4 add_4606_18_lut (.I0(GND_net), .I1(n9204[15]), .I2(GND_net), 
            .I3(n32175), .O(n9184[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_18 (.CI(n32175), .I0(n9204[15]), .I1(GND_net), .CO(n32176));
    SB_LUT4 add_4606_17_lut (.I0(GND_net), .I1(n9204[14]), .I2(GND_net), 
            .I3(n32174), .O(n9184[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n30489), .I0(GND_net), .I1(n1[12]), 
            .CO(n30490));
    SB_CARRY add_4606_17 (.CI(n32174), .I0(n9204[14]), .I1(GND_net), .CO(n32175));
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1[11]), 
            .I3(n30488), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4584_15_lut (.I0(GND_net), .I1(n8907[12]), .I2(GND_net), 
            .I3(n31929), .O(n8887[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4584_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4606_16_lut (.I0(GND_net), .I1(n9204[13]), .I2(GND_net), 
            .I3(n32173), .O(n9184[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4584_15 (.CI(n31929), .I0(n8907[12]), .I1(GND_net), .CO(n31930));
    SB_CARRY add_4606_16 (.CI(n32173), .I0(n9204[13]), .I1(GND_net), .CO(n32174));
    SB_LUT4 add_4584_14_lut (.I0(GND_net), .I1(n8907[11]), .I2(GND_net), 
            .I3(n31928), .O(n8887[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4584_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4584_14 (.CI(n31928), .I0(n8907[11]), .I1(GND_net), .CO(n31929));
    SB_LUT4 add_4606_15_lut (.I0(GND_net), .I1(n9204[12]), .I2(GND_net), 
            .I3(n32172), .O(n9184[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_15 (.CI(n32172), .I0(n9204[12]), .I1(GND_net), .CO(n32173));
    SB_LUT4 add_4606_14_lut (.I0(GND_net), .I1(n9204[11]), .I2(GND_net), 
            .I3(n32171), .O(n9184[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4584_13_lut (.I0(GND_net), .I1(n8907[10]), .I2(GND_net), 
            .I3(n31927), .O(n8887[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4584_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_14 (.CI(n32171), .I0(n9204[11]), .I1(GND_net), .CO(n32172));
    SB_CARRY add_4584_13 (.CI(n31927), .I0(n8907[10]), .I1(GND_net), .CO(n31928));
    SB_LUT4 add_4606_13_lut (.I0(GND_net), .I1(n9204[10]), .I2(GND_net), 
            .I3(n32170), .O(n9184[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n30488), .I0(GND_net), .I1(n1[11]), 
            .CO(n30489));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1[10]), 
            .I3(n30487), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4584_12_lut (.I0(GND_net), .I1(n8907[9]), .I2(GND_net), 
            .I3(n31926), .O(n8887[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4584_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[8]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n30487), .I0(GND_net), .I1(n1[10]), 
            .CO(n30488));
    SB_CARRY add_4606_13 (.CI(n32170), .I0(n9204[10]), .I1(GND_net), .CO(n32171));
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1[9]), 
            .I3(n30486), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4584_12 (.CI(n31926), .I0(n8907[9]), .I1(GND_net), .CO(n31927));
    SB_LUT4 add_4584_11_lut (.I0(GND_net), .I1(n8907[8]), .I2(GND_net), 
            .I3(n31925), .O(n8887[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4584_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4606_12_lut (.I0(GND_net), .I1(n9204[9]), .I2(GND_net), 
            .I3(n32169), .O(n9184[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4584_11 (.CI(n31925), .I0(n8907[8]), .I1(GND_net), .CO(n31926));
    SB_CARRY add_4606_12 (.CI(n32169), .I0(n9204[9]), .I1(GND_net), .CO(n32170));
    SB_LUT4 add_4584_10_lut (.I0(GND_net), .I1(n8907[7]), .I2(GND_net), 
            .I3(n31924), .O(n8887[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4584_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4606_11_lut (.I0(GND_net), .I1(n9204[8]), .I2(GND_net), 
            .I3(n32168), .O(n9184[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4584_10 (.CI(n31924), .I0(n8907[7]), .I1(GND_net), .CO(n31925));
    SB_CARRY add_4606_11 (.CI(n32168), .I0(n9204[8]), .I1(GND_net), .CO(n32169));
    SB_LUT4 add_4584_9_lut (.I0(GND_net), .I1(n8907[6]), .I2(GND_net), 
            .I3(n31923), .O(n8887[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4584_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n30486), .I0(GND_net), .I1(n1[9]), 
            .CO(n30487));
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1[8]), 
            .I3(n30485), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n30485), .I0(GND_net), .I1(n1[8]), 
            .CO(n30486));
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4584_9 (.CI(n31923), .I0(n8907[6]), .I1(GND_net), .CO(n31924));
    SB_LUT4 add_4584_8_lut (.I0(GND_net), .I1(n8907[5]), .I2(n527_adj_3591), 
            .I3(n31922), .O(n8887[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4584_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4584_8 (.CI(n31922), .I0(n8907[5]), .I1(n527_adj_3591), 
            .CO(n31923));
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1[7]), 
            .I3(n30484), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4584_7_lut (.I0(GND_net), .I1(n8907[4]), .I2(n454_adj_3589), 
            .I3(n31921), .O(n8887[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4584_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4584_7 (.CI(n31921), .I0(n8907[4]), .I1(n454_adj_3589), 
            .CO(n31922));
    SB_LUT4 add_4606_10_lut (.I0(GND_net), .I1(n9204[7]), .I2(GND_net), 
            .I3(n32167), .O(n9184[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_10 (.CI(n32167), .I0(n9204[7]), .I1(GND_net), .CO(n32168));
    SB_LUT4 add_4584_6_lut (.I0(GND_net), .I1(n8907[3]), .I2(n381_adj_3588), 
            .I3(n31920), .O(n8887[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4584_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_3598));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4584_6 (.CI(n31920), .I0(n8907[3]), .I1(n381_adj_3588), 
            .CO(n31921));
    SB_LUT4 add_4606_9_lut (.I0(GND_net), .I1(n9204[6]), .I2(GND_net), 
            .I3(n32166), .O(n9184[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_9 (.CI(n32166), .I0(n9204[6]), .I1(GND_net), .CO(n32167));
    SB_LUT4 add_4584_5_lut (.I0(GND_net), .I1(n8907[2]), .I2(n308_adj_3587), 
            .I3(n31919), .O(n8887[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4584_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4584_5 (.CI(n31919), .I0(n8907[2]), .I1(n308_adj_3587), 
            .CO(n31920));
    SB_LUT4 add_4606_8_lut (.I0(GND_net), .I1(n9204[5]), .I2(n527), .I3(n32165), 
            .O(n9184[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4584_4_lut (.I0(GND_net), .I1(n8907[1]), .I2(n235_adj_3586), 
            .I3(n31918), .O(n8887[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4584_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4584_4 (.CI(n31918), .I0(n8907[1]), .I1(n235_adj_3586), 
            .CO(n31919));
    SB_CARRY add_4606_8 (.CI(n32165), .I0(n9204[5]), .I1(n527), .CO(n32166));
    SB_LUT4 add_4606_7_lut (.I0(GND_net), .I1(n9204[4]), .I2(n454), .I3(n32164), 
            .O(n9184[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4584_3_lut (.I0(GND_net), .I1(n8907[0]), .I2(n162_adj_3585), 
            .I3(n31917), .O(n8887[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4584_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4584_3 (.CI(n31917), .I0(n8907[0]), .I1(n162_adj_3585), 
            .CO(n31918));
    SB_LUT4 add_4584_2_lut (.I0(GND_net), .I1(n20_adj_3584), .I2(n89_adj_3582), 
            .I3(GND_net), .O(n8887[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4584_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4584_2 (.CI(GND_net), .I0(n20_adj_3584), .I1(n89_adj_3582), 
            .CO(n31917));
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4606_7 (.CI(n32164), .I0(n9204[4]), .I1(n454), .CO(n32165));
    SB_LUT4 add_4606_6_lut (.I0(GND_net), .I1(n9204[3]), .I2(n381), .I3(n32163), 
            .O(n9184[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_6 (.CI(n32163), .I0(n9204[3]), .I1(n381), .CO(n32164));
    SB_LUT4 add_4583_20_lut (.I0(GND_net), .I1(n8887[17]), .I2(GND_net), 
            .I3(n31916), .O(n8866[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4583_19_lut (.I0(GND_net), .I1(n8887[16]), .I2(GND_net), 
            .I3(n31915), .O(n8866[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4583_19 (.CI(n31915), .I0(n8887[16]), .I1(GND_net), .CO(n31916));
    SB_LUT4 add_4606_5_lut (.I0(GND_net), .I1(n9204[2]), .I2(n308), .I3(n32162), 
            .O(n9184[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4583_18_lut (.I0(GND_net), .I1(n8887[15]), .I2(GND_net), 
            .I3(n31914), .O(n8866[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4583_18 (.CI(n31914), .I0(n8887[15]), .I1(GND_net), .CO(n31915));
    SB_LUT4 add_4583_17_lut (.I0(GND_net), .I1(n8887[14]), .I2(GND_net), 
            .I3(n31913), .O(n8866[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_5 (.CI(n32162), .I0(n9204[2]), .I1(n308), .CO(n32163));
    SB_LUT4 add_4606_4_lut (.I0(GND_net), .I1(n9204[1]), .I2(n235), .I3(n32161), 
            .O(n9184[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4583_17 (.CI(n31913), .I0(n8887[14]), .I1(GND_net), .CO(n31914));
    SB_LUT4 add_4583_16_lut (.I0(GND_net), .I1(n8887[13]), .I2(GND_net), 
            .I3(n31912), .O(n8866[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4606_4 (.CI(n32161), .I0(n9204[1]), .I1(n235), .CO(n32162));
    SB_LUT4 add_4606_3_lut (.I0(GND_net), .I1(n9204[0]), .I2(n162), .I3(n32160), 
            .O(n9184[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4583_16 (.CI(n31912), .I0(n8887[13]), .I1(GND_net), .CO(n31913));
    SB_CARRY add_4606_3 (.CI(n32160), .I0(n9204[0]), .I1(n162), .CO(n32161));
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4606_2_lut (.I0(GND_net), .I1(n20_adj_3581), .I2(n89), 
            .I3(GND_net), .O(n9184[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4606_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4583_15_lut (.I0(GND_net), .I1(n8887[12]), .I2(GND_net), 
            .I3(n31911), .O(n8866[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4583_15 (.CI(n31911), .I0(n8887[12]), .I1(GND_net), .CO(n31912));
    SB_CARRY add_4606_2 (.CI(GND_net), .I0(n20_adj_3581), .I1(n89), .CO(n32160));
    SB_LUT4 add_4605_20_lut (.I0(GND_net), .I1(n9184[17]), .I2(GND_net), 
            .I3(n32159), .O(n9163[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4605_19_lut (.I0(GND_net), .I1(n9184[16]), .I2(GND_net), 
            .I3(n32158), .O(n9163[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_19 (.CI(n32158), .I0(n9184[16]), .I1(GND_net), .CO(n32159));
    SB_LUT4 add_4583_14_lut (.I0(GND_net), .I1(n8887[11]), .I2(GND_net), 
            .I3(n31910), .O(n8866[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4605_18_lut (.I0(GND_net), .I1(n9184[15]), .I2(GND_net), 
            .I3(n32157), .O(n9163[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n30484), .I0(GND_net), .I1(n1[7]), 
            .CO(n30485));
    SB_CARRY add_4583_14 (.CI(n31910), .I0(n8887[11]), .I1(GND_net), .CO(n31911));
    SB_LUT4 add_4583_13_lut (.I0(GND_net), .I1(n8887[10]), .I2(GND_net), 
            .I3(n31909), .O(n8866[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4583_13 (.CI(n31909), .I0(n8887[10]), .I1(GND_net), .CO(n31910));
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1[6]), 
            .I3(n30483), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_18 (.CI(n32157), .I0(n9184[15]), .I1(GND_net), .CO(n32158));
    SB_LUT4 add_4583_12_lut (.I0(GND_net), .I1(n8887[9]), .I2(GND_net), 
            .I3(n31908), .O(n8866[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4583_12 (.CI(n31908), .I0(n8887[9]), .I1(GND_net), .CO(n31909));
    SB_LUT4 add_4605_17_lut (.I0(GND_net), .I1(n9184[14]), .I2(GND_net), 
            .I3(n32156), .O(n9163[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4583_11_lut (.I0(GND_net), .I1(n8887[8]), .I2(GND_net), 
            .I3(n31907), .O(n8866[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n30483), .I0(GND_net), .I1(n1[6]), 
            .CO(n30484));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1[5]), 
            .I3(n30482), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4583_11 (.CI(n31907), .I0(n8887[8]), .I1(GND_net), .CO(n31908));
    SB_CARRY add_4605_17 (.CI(n32156), .I0(n9184[14]), .I1(GND_net), .CO(n32157));
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4605_16_lut (.I0(GND_net), .I1(n9184[13]), .I2(GND_net), 
            .I3(n32155), .O(n9163[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_16 (.CI(n32155), .I0(n9184[13]), .I1(GND_net), .CO(n32156));
    SB_LUT4 add_4583_10_lut (.I0(GND_net), .I1(n8887[7]), .I2(GND_net), 
            .I3(n31906), .O(n8866[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4583_10 (.CI(n31906), .I0(n8887[7]), .I1(GND_net), .CO(n31907));
    SB_LUT4 add_4605_15_lut (.I0(GND_net), .I1(n9184[12]), .I2(GND_net), 
            .I3(n32154), .O(n9163[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4583_9_lut (.I0(GND_net), .I1(n8887[6]), .I2(GND_net), 
            .I3(n31905), .O(n8866[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4605_15 (.CI(n32154), .I0(n9184[12]), .I1(GND_net), .CO(n32155));
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_3596));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4583_9 (.CI(n31905), .I0(n8887[6]), .I1(GND_net), .CO(n31906));
    SB_CARRY unary_minus_16_add_3_7 (.CI(n30482), .I0(GND_net), .I1(n1[5]), 
            .CO(n30483));
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4605_14_lut (.I0(GND_net), .I1(n9184[11]), .I2(GND_net), 
            .I3(n32153), .O(n9163[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(PWMLimit[20]), .I1(duty[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4583_8_lut (.I0(GND_net), .I1(n8887[5]), .I2(n524_adj_3579), 
            .I3(n31904), .O(n8866[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(PWMLimit[19]), .I1(duty[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4583_8 (.CI(n31904), .I0(n8887[5]), .I1(n524_adj_3579), 
            .CO(n31905));
    SB_LUT4 add_4583_7_lut (.I0(GND_net), .I1(n8887[4]), .I2(n451), .I3(n31903), 
            .O(n8866[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_14 (.CI(n32153), .I0(n9184[11]), .I1(GND_net), .CO(n32154));
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(PWMLimit[22]), .I1(duty[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4605_13_lut (.I0(GND_net), .I1(n9184[10]), .I2(GND_net), 
            .I3(n32152), .O(n9163[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4583_7 (.CI(n31903), .I0(n8887[4]), .I1(n451), .CO(n31904));
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(PWMLimit[18]), .I1(duty[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(PWMLimit[14]), .I1(duty[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(PWMLimit[15]), .I1(duty[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(PWMLimit[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_3606));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(PWMLimit[12]), .I1(duty[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_c));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4605_13 (.CI(n32152), .I0(n9184[10]), .I1(GND_net), .CO(n32153));
    SB_LUT4 add_4605_12_lut (.I0(GND_net), .I1(n9184[9]), .I2(GND_net), 
            .I3(n32151), .O(n9163[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4583_6_lut (.I0(GND_net), .I1(n8887[3]), .I2(n378), .I3(n31902), 
            .O(n8866[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1[4]), 
            .I3(n30481), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_12 (.CI(n32151), .I0(n9184[9]), .I1(GND_net), .CO(n32152));
    SB_CARRY add_4583_6 (.CI(n31902), .I0(n8887[3]), .I1(n378), .CO(n31903));
    SB_LUT4 add_4583_5_lut (.I0(GND_net), .I1(n8887[2]), .I2(n305), .I3(n31901), 
            .O(n8866[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4605_11_lut (.I0(GND_net), .I1(n9184[8]), .I2(GND_net), 
            .I3(n32150), .O(n9163[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4583_5 (.CI(n31901), .I0(n8887[2]), .I1(n305), .CO(n31902));
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(PWMLimit[17]), .I1(duty[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n30481), .I0(GND_net), .I1(n1[4]), 
            .CO(n30482));
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(PWMLimit[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_3607));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4605_11 (.CI(n32150), .I0(n9184[8]), .I1(GND_net), .CO(n32151));
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(PWMLimit[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_3608));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4605_10_lut (.I0(GND_net), .I1(n9184[7]), .I2(GND_net), 
            .I3(n32149), .O(n9163[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_10 (.CI(n32149), .I0(n9184[7]), .I1(GND_net), .CO(n32150));
    SB_LUT4 add_4605_9_lut (.I0(GND_net), .I1(n9184[6]), .I2(GND_net), 
            .I3(n32148), .O(n9163[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_9 (.CI(n32148), .I0(n9184[6]), .I1(GND_net), .CO(n32149));
    SB_LUT4 add_4583_4_lut (.I0(GND_net), .I1(n8887[1]), .I2(n232), .I3(n31900), 
            .O(n8866[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4605_8_lut (.I0(GND_net), .I1(n9184[5]), .I2(n524), .I3(n32147), 
            .O(n9163[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_8 (.CI(n32147), .I0(n9184[5]), .I1(n524), .CO(n32148));
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[9]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4605_7_lut (.I0(GND_net), .I1(n9184[4]), .I2(n451_adj_3610), 
            .I3(n32146), .O(n9163[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(PWMLimit[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_3611));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4583_4 (.CI(n31900), .I0(n8887[1]), .I1(n232), .CO(n31901));
    SB_LUT4 add_4583_3_lut (.I0(GND_net), .I1(n8887[0]), .I2(n159), .I3(n31899), 
            .O(n8866[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4583_3 (.CI(n31899), .I0(n8887[0]), .I1(n159), .CO(n31900));
    SB_CARRY add_4605_7 (.CI(n32146), .I0(n9184[4]), .I1(n451_adj_3610), 
            .CO(n32147));
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(PWMLimit[13]), .I1(duty[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4583_2_lut (.I0(GND_net), .I1(n17_adj_3612), .I2(n86), 
            .I3(GND_net), .O(n8866[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4583_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4583_2 (.CI(GND_net), .I0(n17_adj_3612), .I1(n86), .CO(n31899));
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1[3]), 
            .I3(n30480), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(PWMLimit[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_3613));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4605_6_lut (.I0(GND_net), .I1(n9184[3]), .I2(n378_adj_3614), 
            .I3(n32145), .O(n9163[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4582_21_lut (.I0(GND_net), .I1(n8866[18]), .I2(GND_net), 
            .I3(n31898), .O(n8844[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4582_20_lut (.I0(GND_net), .I1(n8866[17]), .I2(GND_net), 
            .I3(n31897), .O(n8844[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(PWMLimit[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_3615));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_4582_20 (.CI(n31897), .I0(n8866[17]), .I1(GND_net), .CO(n31898));
    SB_CARRY add_4605_6 (.CI(n32145), .I0(n9184[3]), .I1(n378_adj_3614), 
            .CO(n32146));
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(PWMLimit[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_3616));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[10]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4582_19_lut (.I0(GND_net), .I1(n8866[16]), .I2(GND_net), 
            .I3(n31896), .O(n8844[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4582_19 (.CI(n31896), .I0(n8866[16]), .I1(GND_net), .CO(n31897));
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(PWMLimit[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_3618));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_4582_18_lut (.I0(GND_net), .I1(n8866[15]), .I2(GND_net), 
            .I3(n31895), .O(n8844[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4582_18 (.CI(n31895), .I0(n8866[15]), .I1(GND_net), .CO(n31896));
    SB_LUT4 add_4605_5_lut (.I0(GND_net), .I1(n9184[2]), .I2(n305_adj_3619), 
            .I3(n32144), .O(n9163[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4582_17_lut (.I0(GND_net), .I1(n8866[14]), .I2(GND_net), 
            .I3(n31894), .O(n8844[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4582_17 (.CI(n31894), .I0(n8866[14]), .I1(GND_net), .CO(n31895));
    SB_LUT4 i36392_4_lut (.I0(n21_adj_3618), .I1(n19_adj_3616), .I2(n17_adj_3615), 
            .I3(n9_adj_3613), .O(n43517));
    defparam i36392_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36344_4_lut (.I0(n27), .I1(n15_adj_3611), .I2(n13_adj_3608), 
            .I3(n11_adj_3607), .O(n43469));
    defparam i36344_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12_adj_3620), .I1(duty[17]), .I2(n35), 
            .I3(GND_net), .O(n30));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37028_4_lut (.I0(n13_adj_3608), .I1(n11_adj_3607), .I2(n9_adj_3613), 
            .I3(n43545), .O(n44153));
    defparam i37028_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_4582_16_lut (.I0(GND_net), .I1(n8866[13]), .I2(GND_net), 
            .I3(n31893), .O(n8844[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37018_4_lut (.I0(n19_adj_3616), .I1(n17_adj_3615), .I2(n15_adj_3611), 
            .I3(n44153), .O(n44143));
    defparam i37018_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_4605_5 (.CI(n32144), .I0(n9184[2]), .I1(n305_adj_3619), 
            .CO(n32145));
    SB_CARRY add_4582_16 (.CI(n31893), .I0(n8866[13]), .I1(GND_net), .CO(n31894));
    SB_LUT4 add_4582_15_lut (.I0(GND_net), .I1(n8866[12]), .I2(GND_net), 
            .I3(n31892), .O(n8844[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37791_4_lut (.I0(n25_c), .I1(n23_adj_3606), .I2(n21_adj_3618), 
            .I3(n44143), .O(n44916));
    defparam i37791_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i37332_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n44916), 
            .O(n44457));
    defparam i37332_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i37891_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n44457), 
            .O(n45016));
    defparam i37891_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_4605_4_lut (.I0(GND_net), .I1(n9184[1]), .I2(n232_adj_3621), 
            .I3(n32143), .O(n9163[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_4 (.CI(n32143), .I0(n9184[1]), .I1(n232_adj_3621), 
            .CO(n32144));
    SB_CARRY add_4582_15 (.CI(n31892), .I0(n8866[12]), .I1(GND_net), .CO(n31893));
    SB_LUT4 i37549_3_lut (.I0(n6_adj_3622), .I1(duty[10]), .I2(n21_adj_3618), 
            .I3(GND_net), .O(n44674));   // verilog/motorControl.v(44[10:25])
    defparam i37549_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_4582_14_lut (.I0(GND_net), .I1(n8866[11]), .I2(GND_net), 
            .I3(n31891), .O(n8844[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n30480), .I0(GND_net), .I1(n1[3]), 
            .CO(n30481));
    SB_LUT4 add_4605_3_lut (.I0(GND_net), .I1(n9184[0]), .I2(n159_adj_3623), 
            .I3(n32142), .O(n9163[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4582_14 (.CI(n31891), .I0(n8866[11]), .I1(GND_net), .CO(n31892));
    SB_LUT4 i37550_3_lut (.I0(n44674), .I1(duty[11]), .I2(n23_adj_3606), 
            .I3(GND_net), .O(n44675));   // verilog/motorControl.v(44[10:25])
    defparam i37550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16_adj_3624), .I1(duty[22]), .I2(n45), 
            .I3(GND_net), .O(n24));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36267_4_lut (.I0(n43), .I1(n25_c), .I2(n23_adj_3606), .I3(n43517), 
            .O(n43392));
    defparam i36267_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1[2]), 
            .I3(n30479), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4605_3 (.CI(n32142), .I0(n9184[0]), .I1(n159_adj_3623), 
            .CO(n32143));
    SB_LUT4 add_4582_13_lut (.I0(GND_net), .I1(n8866[10]), .I2(GND_net), 
            .I3(n31890), .O(n8844[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4582_13 (.CI(n31890), .I0(n8866[10]), .I1(GND_net), .CO(n31891));
    SB_LUT4 add_4605_2_lut (.I0(GND_net), .I1(n17_adj_3626), .I2(n86_adj_3627), 
            .I3(GND_net), .O(n9163[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4605_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37486_4_lut (.I0(n24), .I1(n8_adj_3628), .I2(n45), .I3(n43388), 
            .O(n44611));   // verilog/motorControl.v(44[10:25])
    defparam i37486_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_4605_2 (.CI(GND_net), .I0(n17_adj_3626), .I1(n86_adj_3627), 
            .CO(n32142));
    SB_LUT4 add_4604_21_lut (.I0(GND_net), .I1(n9163[18]), .I2(GND_net), 
            .I3(n32141), .O(n9141[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4582_12_lut (.I0(GND_net), .I1(n8866[9]), .I2(GND_net), 
            .I3(n31889), .O(n8844[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36761_3_lut (.I0(n44675), .I1(duty[12]), .I2(n25_c), .I3(GND_net), 
            .O(n43886));   // verilog/motorControl.v(44[10:25])
    defparam i36761_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4582_12 (.CI(n31889), .I0(n8866[9]), .I1(GND_net), .CO(n31890));
    SB_LUT4 add_4582_11_lut (.I0(GND_net), .I1(n8866[8]), .I2(GND_net), 
            .I3(n31888), .O(n8844[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4604_20_lut (.I0(GND_net), .I1(n9163[17]), .I2(GND_net), 
            .I3(n32140), .O(n9141[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_20 (.CI(n32140), .I0(n9163[17]), .I1(GND_net), .CO(n32141));
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(PWMLimit[1]), 
            .I3(PWMLimit[0]), .O(n4_adj_3629));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_CARRY add_4582_11 (.CI(n31888), .I0(n8866[8]), .I1(GND_net), .CO(n31889));
    SB_LUT4 i37544_3_lut (.I0(n4_adj_3629), .I1(duty[13]), .I2(n27), .I3(GND_net), 
            .O(n44669));   // verilog/motorControl.v(44[10:25])
    defparam i37544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37545_3_lut (.I0(n44669), .I1(duty[14]), .I2(n29), .I3(GND_net), 
            .O(n44670));   // verilog/motorControl.v(44[10:25])
    defparam i37545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36296_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n43469), 
            .O(n43421));
    defparam i36296_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37833_4_lut (.I0(n30), .I1(n10_adj_3630), .I2(n35), .I3(n43416), 
            .O(n44958));   // verilog/motorControl.v(44[10:25])
    defparam i37833_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36763_3_lut (.I0(n44670), .I1(duty[15]), .I2(n31), .I3(GND_net), 
            .O(n43888));   // verilog/motorControl.v(44[10:25])
    defparam i36763_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n30479), .I0(GND_net), .I1(n1[2]), 
            .CO(n30480));
    SB_LUT4 add_4582_10_lut (.I0(GND_net), .I1(n8866[7]), .I2(GND_net), 
            .I3(n31887), .O(n8844[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1[1]), 
            .I3(n30478), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4604_19_lut (.I0(GND_net), .I1(n9163[16]), .I2(GND_net), 
            .I3(n32139), .O(n9141[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_19 (.CI(n32139), .I0(n9163[16]), .I1(GND_net), .CO(n32140));
    SB_CARRY add_4582_10 (.CI(n31887), .I0(n8866[7]), .I1(GND_net), .CO(n31888));
    SB_LUT4 add_4582_9_lut (.I0(GND_net), .I1(n8866[6]), .I2(GND_net), 
            .I3(n31886), .O(n8844[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4582_9 (.CI(n31886), .I0(n8866[6]), .I1(GND_net), .CO(n31887));
    SB_LUT4 add_4604_18_lut (.I0(GND_net), .I1(n9163[15]), .I2(GND_net), 
            .I3(n32138), .O(n9141[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i37965_4_lut (.I0(n43888), .I1(n44958), .I2(n35), .I3(n43421), 
            .O(n45090));   // verilog/motorControl.v(44[10:25])
    defparam i37965_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_4604_18 (.CI(n32138), .I0(n9163[15]), .I1(GND_net), .CO(n32139));
    SB_LUT4 i37966_3_lut (.I0(n45090), .I1(duty[18]), .I2(n37), .I3(GND_net), 
            .O(n45091));   // verilog/motorControl.v(44[10:25])
    defparam i37966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37935_3_lut (.I0(n45091), .I1(duty[19]), .I2(n39), .I3(GND_net), 
            .O(n45060));   // verilog/motorControl.v(44[10:25])
    defparam i37935_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21493_1_lut (.I0(n256), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n26500));   // verilog/motorControl.v(46[19:35])
    defparam i21493_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4604_17_lut (.I0(GND_net), .I1(n9163[14]), .I2(GND_net), 
            .I3(n32137), .O(n9141[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4582_8_lut (.I0(GND_net), .I1(n8866[5]), .I2(n521), .I3(n31885), 
            .O(n8844[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36269_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n45016), 
            .O(n43394));
    defparam i36269_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_4604_17 (.CI(n32137), .I0(n9163[14]), .I1(GND_net), .CO(n32138));
    SB_LUT4 i37705_4_lut (.I0(n43886), .I1(n44611), .I2(n45), .I3(n43392), 
            .O(n44830));   // verilog/motorControl.v(44[10:25])
    defparam i37705_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_4582_8 (.CI(n31885), .I0(n8866[5]), .I1(n521), .CO(n31886));
    SB_LUT4 add_4582_7_lut (.I0(GND_net), .I1(n8866[4]), .I2(n448), .I3(n31884), 
            .O(n8844[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n30478), .I0(GND_net), .I1(n1[1]), 
            .CO(n30479));
    SB_LUT4 i36769_3_lut (.I0(n45060), .I1(duty[20]), .I2(n41), .I3(GND_net), 
            .O(n43894));   // verilog/motorControl.v(44[10:25])
    defparam i36769_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4582_7 (.CI(n31884), .I0(n8866[4]), .I1(n448), .CO(n31885));
    SB_LUT4 add_4582_6_lut (.I0(GND_net), .I1(n8866[3]), .I2(n375), .I3(n31883), 
            .O(n8844[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n25), .I1(GND_net), .I2(n1[0]), 
            .I3(VCC_net), .O(n42863)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i37867_4_lut (.I0(n43894), .I1(n44830), .I2(n45), .I3(n43394), 
            .O(n44992));   // verilog/motorControl.v(44[10:25])
    defparam i37867_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1[0]), 
            .CO(n30478));
    SB_LUT4 i37868_3_lut (.I0(n44992), .I1(PWMLimit[23]), .I2(duty[23]), 
            .I3(GND_net), .O(duty_23__N_3502));   // verilog/motorControl.v(44[10:25])
    defparam i37868_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_4604_16_lut (.I0(GND_net), .I1(n9163[13]), .I2(GND_net), 
            .I3(n32136), .O(n9141[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3897[23]), 
            .I3(n30477), .O(\PID_CONTROLLER.integral_23__N_3454 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_3635));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4582_6 (.CI(n31883), .I0(n8866[3]), .I1(n375), .CO(n31884));
    SB_CARRY add_4604_16 (.CI(n32136), .I0(n9163[13]), .I1(GND_net), .CO(n32137));
    SB_LUT4 add_4582_5_lut (.I0(GND_net), .I1(n8866[2]), .I2(n302), .I3(n31882), 
            .O(n8844[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4604_15_lut (.I0(GND_net), .I1(n9163[12]), .I2(GND_net), 
            .I3(n32135), .O(n9141[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4582_5 (.CI(n31882), .I0(n8866[2]), .I1(n302), .CO(n31883));
    SB_LUT4 add_4582_4_lut (.I0(GND_net), .I1(n8866[1]), .I2(n229), .I3(n31881), 
            .O(n8844[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_15 (.CI(n32135), .I0(n9163[12]), .I1(GND_net), .CO(n32136));
    SB_LUT4 add_4604_14_lut (.I0(GND_net), .I1(n9163[11]), .I2(GND_net), 
            .I3(n32134), .O(n9141[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1_adj_3897[22]), .I3(n30476), .O(n45_adj_3636)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3638));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i1_3_lut (.I0(duty_23__N_3478[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[0]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_4604_14 (.CI(n32134), .I0(n9163[11]), .I1(GND_net), .CO(n32135));
    SB_CARRY add_4582_4 (.CI(n31881), .I0(n8866[1]), .I1(n229), .CO(n31882));
    SB_LUT4 add_4582_3_lut (.I0(GND_net), .I1(n8866[0]), .I2(n156), .I3(n31880), 
            .O(n8844[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_3595));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_3639));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4582_3 (.CI(n31880), .I0(n8866[0]), .I1(n156), .CO(n31881));
    SB_LUT4 add_4604_13_lut (.I0(GND_net), .I1(n9163[10]), .I2(GND_net), 
            .I3(n32133), .O(n9141[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_3594));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n30476), .I0(GND_net), .I1(n1_adj_3897[22]), 
            .CO(n30477));
    SB_LUT4 add_4582_2_lut (.I0(GND_net), .I1(n14_adj_3640), .I2(n83), 
            .I3(GND_net), .O(n8844[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4582_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_13 (.CI(n32133), .I0(n9163[10]), .I1(GND_net), .CO(n32134));
    SB_LUT4 add_4604_12_lut (.I0(GND_net), .I1(n9163[9]), .I2(GND_net), 
            .I3(n32132), .O(n9141[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_12 (.CI(n32132), .I0(n9163[9]), .I1(GND_net), .CO(n32133));
    SB_CARRY add_4582_2 (.CI(GND_net), .I0(n14_adj_3640), .I1(n83), .CO(n31880));
    SB_LUT4 add_4581_22_lut (.I0(GND_net), .I1(n8844[19]), .I2(GND_net), 
            .I3(n31879), .O(n8821[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4581_21_lut (.I0(GND_net), .I1(n8844[18]), .I2(GND_net), 
            .I3(n31878), .O(n8821[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1_adj_3897[21]), .I3(n30475), .O(n43_adj_3641)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4581_21 (.CI(n31878), .I0(n8844[18]), .I1(GND_net), .CO(n31879));
    SB_CARRY unary_minus_5_add_3_23 (.CI(n30475), .I0(GND_net), .I1(n1_adj_3897[21]), 
            .CO(n30476));
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1_adj_3897[20]), .I3(n30474), .O(n41_adj_3643)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n30474), .I0(GND_net), .I1(n1_adj_3897[20]), 
            .CO(n30475));
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1_adj_3897[19]), .I3(n30473), .O(n39_adj_3645)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n30473), .I0(GND_net), .I1(n1_adj_3897[19]), 
            .CO(n30474));
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1_adj_3897[18]), .I3(n30472), .O(n37_adj_3647)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_3649));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n30472), .I0(GND_net), .I1(n1_adj_3897[18]), 
            .CO(n30473));
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1_adj_3897[17]), .I3(n30471), .O(n35_adj_3650)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n30471), .I0(GND_net), .I1(n1_adj_3897[17]), 
            .CO(n30472));
    SB_LUT4 add_4581_20_lut (.I0(GND_net), .I1(n8844[17]), .I2(GND_net), 
            .I3(n31877), .O(n8821[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4604_11_lut (.I0(GND_net), .I1(n9163[8]), .I2(GND_net), 
            .I3(n32131), .O(n9141[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4581_20 (.CI(n31877), .I0(n8844[17]), .I1(GND_net), .CO(n31878));
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1_adj_3897[16]), .I3(n30470), .O(n33_adj_3652)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n30470), .I0(GND_net), .I1(n1_adj_3897[16]), 
            .CO(n30471));
    SB_CARRY add_4604_11 (.CI(n32131), .I0(n9163[8]), .I1(GND_net), .CO(n32132));
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_3654));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1_adj_3897[15]), .I3(n30469), .O(n31_adj_3655)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_3657));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_3658));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4604_10_lut (.I0(GND_net), .I1(n9163[7]), .I2(GND_net), 
            .I3(n32130), .O(n9141[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_17 (.CI(n30469), .I0(GND_net), .I1(n1_adj_3897[15]), 
            .CO(n30470));
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1_adj_3897[14]), .I3(n30468), .O(n29_adj_3659)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4581_19_lut (.I0(GND_net), .I1(n8844[16]), .I2(GND_net), 
            .I3(n31876), .O(n8821[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_10 (.CI(n32130), .I0(n9163[7]), .I1(GND_net), .CO(n32131));
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4604_9_lut (.I0(GND_net), .I1(n9163[6]), .I2(GND_net), 
            .I3(n32129), .O(n9141[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4581_19 (.CI(n31876), .I0(n8844[16]), .I1(GND_net), .CO(n31877));
    SB_LUT4 add_4581_18_lut (.I0(GND_net), .I1(n8844[15]), .I2(GND_net), 
            .I3(n31875), .O(n8821[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4604_9 (.CI(n32129), .I0(n9163[6]), .I1(GND_net), .CO(n32130));
    SB_CARRY add_4581_18 (.CI(n31875), .I0(n8844[15]), .I1(GND_net), .CO(n31876));
    SB_CARRY unary_minus_5_add_3_16 (.CI(n30468), .I0(GND_net), .I1(n1_adj_3897[14]), 
            .CO(n30469));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1_adj_3897[13]), .I3(n30467), .O(n27_adj_3661)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4604_8_lut (.I0(GND_net), .I1(n9163[5]), .I2(n521_adj_3663), 
            .I3(n32128), .O(n9141[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4581_17_lut (.I0(GND_net), .I1(n8844[14]), .I2(GND_net), 
            .I3(n31874), .O(n8821[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_8 (.CI(n32128), .I0(n9163[5]), .I1(n521_adj_3663), 
            .CO(n32129));
    SB_CARRY add_4581_17 (.CI(n31874), .I0(n8844[14]), .I1(GND_net), .CO(n31875));
    SB_LUT4 add_4581_16_lut (.I0(GND_net), .I1(n8844[13]), .I2(GND_net), 
            .I3(n31873), .O(n8821[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n30467), .I0(GND_net), .I1(n1_adj_3897[13]), 
            .CO(n30468));
    SB_LUT4 add_4604_7_lut (.I0(GND_net), .I1(n9163[4]), .I2(n448_adj_3664), 
            .I3(n32127), .O(n9141[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4581_16 (.CI(n31873), .I0(n8844[13]), .I1(GND_net), .CO(n31874));
    SB_CARRY add_4604_7 (.CI(n32127), .I0(n9163[4]), .I1(n448_adj_3664), 
            .CO(n32128));
    SB_LUT4 add_4604_6_lut (.I0(GND_net), .I1(n9163[3]), .I2(n375_adj_3665), 
            .I3(n32126), .O(n9141[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4581_15_lut (.I0(GND_net), .I1(n8844[12]), .I2(GND_net), 
            .I3(n31872), .O(n8821[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1_adj_3897[12]), .I3(n30466), .O(n25_adj_3666)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4581_15 (.CI(n31872), .I0(n8844[12]), .I1(GND_net), .CO(n31873));
    SB_CARRY add_4604_6 (.CI(n32126), .I0(n9163[3]), .I1(n375_adj_3665), 
            .CO(n32127));
    SB_LUT4 add_4581_14_lut (.I0(GND_net), .I1(n8844[11]), .I2(GND_net), 
            .I3(n31871), .O(n8821[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4604_5_lut (.I0(GND_net), .I1(n9163[2]), .I2(n302_adj_3668), 
            .I3(n32125), .O(n9141[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_5 (.CI(n32125), .I0(n9163[2]), .I1(n302_adj_3668), 
            .CO(n32126));
    SB_CARRY add_4581_14 (.CI(n31871), .I0(n8844[11]), .I1(GND_net), .CO(n31872));
    SB_LUT4 add_4581_13_lut (.I0(GND_net), .I1(n8844[10]), .I2(GND_net), 
            .I3(n31870), .O(n8821[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4581_13 (.CI(n31870), .I0(n8844[10]), .I1(GND_net), .CO(n31871));
    SB_LUT4 add_4604_4_lut (.I0(GND_net), .I1(n9163[1]), .I2(n229_adj_3669), 
            .I3(n32124), .O(n9141[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_4 (.CI(n32124), .I0(n9163[1]), .I1(n229_adj_3669), 
            .CO(n32125));
    SB_LUT4 add_4581_12_lut (.I0(GND_net), .I1(n8844[9]), .I2(GND_net), 
            .I3(n31869), .O(n8821[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n30466), .I0(GND_net), .I1(n1_adj_3897[12]), 
            .CO(n30467));
    SB_CARRY add_4581_12 (.CI(n31869), .I0(n8844[9]), .I1(GND_net), .CO(n31870));
    SB_LUT4 add_4581_11_lut (.I0(GND_net), .I1(n8844[8]), .I2(GND_net), 
            .I3(n31868), .O(n8821[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4604_3_lut (.I0(GND_net), .I1(n9163[0]), .I2(n156_adj_3670), 
            .I3(n32123), .O(n9141[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4581_11 (.CI(n31868), .I0(n8844[8]), .I1(GND_net), .CO(n31869));
    SB_LUT4 add_4581_10_lut (.I0(GND_net), .I1(n8844[7]), .I2(GND_net), 
            .I3(n31867), .O(n8821[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1_adj_3897[11]), .I3(n30465), .O(n23_adj_3671)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4604_3 (.CI(n32123), .I0(n9163[0]), .I1(n156_adj_3670), 
            .CO(n32124));
    SB_CARRY add_4581_10 (.CI(n31867), .I0(n8844[7]), .I1(GND_net), .CO(n31868));
    SB_LUT4 add_4581_9_lut (.I0(GND_net), .I1(n8844[6]), .I2(GND_net), 
            .I3(n31866), .O(n8821[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n30465), .I0(GND_net), .I1(n1_adj_3897[11]), 
            .CO(n30466));
    SB_LUT4 add_4604_2_lut (.I0(GND_net), .I1(n14_adj_3673), .I2(n83_adj_3674), 
            .I3(GND_net), .O(n9141[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4604_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4604_2 (.CI(GND_net), .I0(n14_adj_3673), .I1(n83_adj_3674), 
            .CO(n32123));
    SB_LUT4 add_4603_22_lut (.I0(GND_net), .I1(n9141[19]), .I2(GND_net), 
            .I3(n32122), .O(n9118[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4581_9 (.CI(n31866), .I0(n8844[6]), .I1(GND_net), .CO(n31867));
    SB_LUT4 add_4603_21_lut (.I0(GND_net), .I1(n9141[18]), .I2(GND_net), 
            .I3(n32121), .O(n9118[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_21 (.CI(n32121), .I0(n9141[18]), .I1(GND_net), .CO(n32122));
    SB_LUT4 add_4603_20_lut (.I0(GND_net), .I1(n9141[17]), .I2(GND_net), 
            .I3(n32120), .O(n9118[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4581_8_lut (.I0(GND_net), .I1(n8844[5]), .I2(n518_adj_3675), 
            .I3(n31865), .O(n8821[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_20 (.CI(n32120), .I0(n9141[17]), .I1(GND_net), .CO(n32121));
    SB_LUT4 add_4603_19_lut (.I0(GND_net), .I1(n9141[16]), .I2(GND_net), 
            .I3(n32119), .O(n9118[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4581_8 (.CI(n31865), .I0(n8844[5]), .I1(n518_adj_3675), 
            .CO(n31866));
    SB_CARRY add_4603_19 (.CI(n32119), .I0(n9141[16]), .I1(GND_net), .CO(n32120));
    SB_LUT4 add_4603_18_lut (.I0(GND_net), .I1(n9141[15]), .I2(GND_net), 
            .I3(n32118), .O(n9118[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4581_7_lut (.I0(GND_net), .I1(n8844[4]), .I2(n445_adj_3658), 
            .I3(n31864), .O(n8821[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4581_7 (.CI(n31864), .I0(n8844[4]), .I1(n445_adj_3658), 
            .CO(n31865));
    SB_CARRY add_4603_18 (.CI(n32118), .I0(n9141[15]), .I1(GND_net), .CO(n32119));
    SB_LUT4 add_4603_17_lut (.I0(GND_net), .I1(n9141[14]), .I2(GND_net), 
            .I3(n32117), .O(n9118[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_17 (.CI(n32117), .I0(n9141[14]), .I1(GND_net), .CO(n32118));
    SB_LUT4 add_4581_6_lut (.I0(GND_net), .I1(n8844[3]), .I2(n372_adj_3657), 
            .I3(n31863), .O(n8821[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4581_6 (.CI(n31863), .I0(n8844[3]), .I1(n372_adj_3657), 
            .CO(n31864));
    SB_LUT4 add_4603_16_lut (.I0(GND_net), .I1(n9141[13]), .I2(GND_net), 
            .I3(n32116), .O(n9118[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4581_5_lut (.I0(GND_net), .I1(n8844[2]), .I2(n299_adj_3654), 
            .I3(n31862), .O(n8821[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4581_5 (.CI(n31862), .I0(n8844[2]), .I1(n299_adj_3654), 
            .CO(n31863));
    SB_CARRY add_4603_16 (.CI(n32116), .I0(n9141[13]), .I1(GND_net), .CO(n32117));
    SB_LUT4 add_4603_15_lut (.I0(GND_net), .I1(n9141[12]), .I2(GND_net), 
            .I3(n32115), .O(n9118[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_15 (.CI(n32115), .I0(n9141[12]), .I1(GND_net), .CO(n32116));
    SB_LUT4 add_4603_14_lut (.I0(GND_net), .I1(n9141[11]), .I2(GND_net), 
            .I3(n32114), .O(n9118[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4581_4_lut (.I0(GND_net), .I1(n8844[1]), .I2(n226_adj_3649), 
            .I3(n31861), .O(n8821[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4581_4 (.CI(n31861), .I0(n8844[1]), .I1(n226_adj_3649), 
            .CO(n31862));
    SB_LUT4 add_4581_3_lut (.I0(GND_net), .I1(n8844[0]), .I2(n153_adj_3639), 
            .I3(n31860), .O(n8821[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4581_3 (.CI(n31860), .I0(n8844[0]), .I1(n153_adj_3639), 
            .CO(n31861));
    SB_LUT4 add_4581_2_lut (.I0(GND_net), .I1(n11_adj_3638), .I2(n80_adj_3635), 
            .I3(GND_net), .O(n8821[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4581_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4581_2 (.CI(GND_net), .I0(n11_adj_3638), .I1(n80_adj_3635), 
            .CO(n31860));
    SB_CARRY add_4603_14 (.CI(n32114), .I0(n9141[11]), .I1(GND_net), .CO(n32115));
    SB_LUT4 mult_10_add_1225_24_lut (.I0(\PID_CONTROLLER.err [23]), .I1(n8797[21]), 
            .I2(GND_net), .I3(n31859), .O(n7831[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(n26500), .I1(n8797[20]), .I2(GND_net), 
            .I3(n31858), .O(n2942[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_4603_13_lut (.I0(GND_net), .I1(n9141[10]), .I2(GND_net), 
            .I3(n32113), .O(n9118[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_13 (.CI(n32113), .I0(n9141[10]), .I1(GND_net), .CO(n32114));
    SB_LUT4 add_4603_12_lut (.I0(GND_net), .I1(n9141[9]), .I2(GND_net), 
            .I3(n32112), .O(n9118[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_12 (.CI(n32112), .I0(n9141[9]), .I1(GND_net), .CO(n32113));
    SB_LUT4 add_4603_11_lut (.I0(GND_net), .I1(n9141[8]), .I2(GND_net), 
            .I3(n32111), .O(n9118[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4603_11 (.CI(n32111), .I0(n9141[8]), .I1(GND_net), .CO(n32112));
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1_adj_3897[10]), .I3(n30464), .O(n21_adj_3676)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_3577));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_3576));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_3575));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_626_i1_4_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(PWMLimit[0]), 
            .I2(n256), .I3(\Ki[0] ), .O(n2967[0]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i1_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 i21299_3_lut (.I0(\Kp[0] ), .I1(n256), .I2(\PID_CONTROLLER.err [0]), 
            .I3(GND_net), .O(n2942[0]));   // verilog/motorControl.v(46[16] 48[10])
    defparam i21299_3_lut.LUT_INIT = 16'hecec;
    SB_CARRY unary_minus_5_add_3_12 (.CI(n30464), .I0(GND_net), .I1(n1_adj_3897[10]), 
            .CO(n30465));
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1_adj_3897[9]), .I3(n30463), .O(n19_adj_3677)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_4603_10_lut (.I0(GND_net), .I1(n9141[7]), .I2(GND_net), 
            .I3(n32110), .O(n9118[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_23 (.CI(n31858), .I0(n8797[20]), .I1(GND_net), 
            .CO(n31859));
    SB_CARRY add_4603_10 (.CI(n32110), .I0(n9141[7]), .I1(GND_net), .CO(n32111));
    SB_LUT4 mult_10_add_1225_22_lut (.I0(n26500), .I1(n8797[19]), .I2(GND_net), 
            .I3(n31857), .O(n2942[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_22 (.CI(n31857), .I0(n8797[19]), .I1(GND_net), 
            .CO(n31858));
    SB_LUT4 mult_10_add_1225_21_lut (.I0(n26500), .I1(n8797[18]), .I2(GND_net), 
            .I3(n31856), .O(n2942[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_21 (.CI(n31856), .I0(n8797[18]), .I1(GND_net), 
            .CO(n31857));
    SB_LUT4 add_4603_9_lut (.I0(GND_net), .I1(n9141[6]), .I2(GND_net), 
            .I3(n32109), .O(n9118[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_20_lut (.I0(n26500), .I1(n8797[17]), .I2(GND_net), 
            .I3(n31855), .O(n2942[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_20 (.CI(n31855), .I0(n8797[17]), .I1(GND_net), 
            .CO(n31856));
    SB_CARRY add_4603_9 (.CI(n32109), .I0(n9141[6]), .I1(GND_net), .CO(n32110));
    SB_LUT4 mult_10_add_1225_19_lut (.I0(n26500), .I1(n8797[16]), .I2(GND_net), 
            .I3(n31854), .O(n2942[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_4603_8_lut (.I0(GND_net), .I1(n9141[5]), .I2(n518), .I3(n32108), 
            .O(n9118[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_19 (.CI(n31854), .I0(n8797[16]), .I1(GND_net), 
            .CO(n31855));
    SB_LUT4 mult_10_add_1225_18_lut (.I0(n26500), .I1(n8797[15]), .I2(GND_net), 
            .I3(n31853), .O(n2942[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4603_8 (.CI(n32108), .I0(n9141[5]), .I1(n518), .CO(n32109));
    SB_LUT4 add_4603_7_lut (.I0(GND_net), .I1(n9141[4]), .I2(n445), .I3(n32107), 
            .O(n9118[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_18 (.CI(n31853), .I0(n8797[15]), .I1(GND_net), 
            .CO(n31854));
    SB_CARRY add_4603_7 (.CI(n32107), .I0(n9141[4]), .I1(n445), .CO(n32108));
    SB_CARRY unary_minus_5_add_3_11 (.CI(n30463), .I0(GND_net), .I1(n1_adj_3897[9]), 
            .CO(n30464));
    SB_LUT4 add_4603_6_lut (.I0(GND_net), .I1(n9141[3]), .I2(n372), .I3(n32106), 
            .O(n9118[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_17_lut (.I0(n26500), .I1(n8797[14]), .I2(GND_net), 
            .I3(n31852), .O(n2942[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4603_6 (.CI(n32106), .I0(n9141[3]), .I1(n372), .CO(n32107));
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1_adj_3897[8]), .I3(n30462), .O(n17_adj_3678)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_CARRY mult_10_add_1225_17 (.CI(n31852), .I0(n8797[14]), .I1(GND_net), 
            .CO(n31853));
    SB_LUT4 add_4603_5_lut (.I0(GND_net), .I1(n9141[2]), .I2(n299), .I3(n32105), 
            .O(n9118[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_16_lut (.I0(n26500), .I1(n8797[13]), .I2(GND_net), 
            .I3(n31851), .O(n2942[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_16 (.CI(n31851), .I0(n8797[13]), .I1(GND_net), 
            .CO(n31852));
    SB_LUT4 mult_10_add_1225_15_lut (.I0(n26500), .I1(n8797[12]), .I2(GND_net), 
            .I3(n31850), .O(n2942[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_3675));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n30462), .I0(GND_net), .I1(n1_adj_3897[8]), 
            .CO(n30463));
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83_adj_3674));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1_adj_3897[7]), .I3(n30461), .O(n15_adj_3679)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_4603_5 (.CI(n32105), .I0(n9141[2]), .I1(n299), .CO(n32106));
    SB_LUT4 add_4603_4_lut (.I0(GND_net), .I1(n9141[1]), .I2(n226), .I3(n32104), 
            .O(n9118[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_15 (.CI(n31850), .I0(n8797[12]), .I1(GND_net), 
            .CO(n31851));
    SB_CARRY add_4603_4 (.CI(n32104), .I0(n9141[1]), .I1(n226), .CO(n32105));
    SB_LUT4 add_4603_3_lut (.I0(GND_net), .I1(n9141[0]), .I2(n153), .I3(n32103), 
            .O(n9118[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_14_lut (.I0(n26500), .I1(n8797[11]), .I2(GND_net), 
            .I3(n31849), .O(n2942[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_4603_3 (.CI(n32103), .I0(n9141[0]), .I1(n153), .CO(n32104));
    SB_CARRY mult_10_add_1225_14 (.CI(n31849), .I0(n8797[11]), .I1(GND_net), 
            .CO(n31850));
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3673));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_add_1225_13_lut (.I0(n26500), .I1(n8797[10]), .I2(GND_net), 
            .I3(n31848), .O(n2942[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_13 (.CI(n31848), .I0(n8797[10]), .I1(GND_net), 
            .CO(n31849));
    SB_LUT4 mult_10_add_1225_12_lut (.I0(n26500), .I1(n8797[9]), .I2(GND_net), 
            .I3(n31847), .O(n2942[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_4603_2_lut (.I0(GND_net), .I1(n11_adj_3583), .I2(n80), 
            .I3(GND_net), .O(n9118[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4603_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_12 (.CI(n31847), .I0(n8797[9]), .I1(GND_net), 
            .CO(n31848));
    SB_LUT4 mult_10_add_1225_11_lut (.I0(n26500), .I1(n8797[8]), .I2(GND_net), 
            .I3(n31846), .O(n2942[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_11 (.CI(n31846), .I0(n8797[8]), .I1(GND_net), 
            .CO(n31847));
    SB_CARRY add_4603_2 (.CI(GND_net), .I0(n11_adj_3583), .I1(n80), .CO(n32103));
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(n9094[21]), 
            .I2(GND_net), .I3(n32102), .O(n42910)) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_1225_10_lut (.I0(n26500), .I1(n8797[7]), .I2(GND_net), 
            .I3(n31845), .O(n2942[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[11]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n30461), .I0(GND_net), .I1(n1_adj_3897[7]), 
            .CO(n30462));
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1_adj_3897[6]), .I3(n30460), .O(n13_adj_3680)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n30460), .I0(GND_net), .I1(n1_adj_3897[6]), 
            .CO(n30461));
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_3572));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_3670));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_626_i2_3_lut (.I0(n155[1]), .I1(PWMLimit[1]), .I2(n256), 
            .I3(GND_net), .O(n2967[1]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i2_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFFE \PID_CONTROLLER.integral_1149__i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[0]));   // verilog/motorControl.v(40[21:33])
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1_adj_3897[5]), .I3(n30459), .O(n11_adj_3681)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n9094[20]), .I2(GND_net), 
            .I3(n32101), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n30459), .I0(GND_net), .I1(n1_adj_3897[5]), 
            .CO(n30460));
    SB_CARRY mult_10_add_1225_10 (.CI(n31845), .I0(n8797[7]), .I1(GND_net), 
            .CO(n31846));
    SB_CARRY mult_11_add_1225_23 (.CI(n32101), .I0(n9094[20]), .I1(GND_net), 
            .CO(n32102));
    SB_LUT4 mult_10_add_1225_9_lut (.I0(n26500), .I1(n8797[6]), .I2(GND_net), 
            .I3(n31844), .O(n2942[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n9094[19]), .I2(GND_net), 
            .I3(n32100), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_9 (.CI(n31844), .I0(n8797[6]), .I1(GND_net), 
            .CO(n31845));
    SB_CARRY mult_11_add_1225_22 (.CI(n32100), .I0(n9094[19]), .I1(GND_net), 
            .CO(n32101));
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n9094[18]), .I2(GND_net), 
            .I3(n32099), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_8_lut (.I0(n26500), .I1(n8797[5]), .I2(n512), 
            .I3(n31843), .O(n2942[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1_adj_3897[4]), .I3(n30458), .O(n9_adj_3683)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_3685));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_8 (.CI(n31843), .I0(n8797[5]), .I1(n512), 
            .CO(n31844));
    SB_LUT4 mult_10_add_1225_7_lut (.I0(n26500), .I1(n8797[4]), .I2(n439), 
            .I3(n31842), .O(n2942[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n30458), .I0(GND_net), .I1(n1_adj_3897[4]), 
            .CO(n30459));
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_3686));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_21 (.CI(n32099), .I0(n9094[18]), .I1(GND_net), 
            .CO(n32100));
    SB_CARRY mult_10_add_1225_7 (.CI(n31842), .I0(n8797[4]), .I1(n439), 
            .CO(n31843));
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n9094[17]), .I2(GND_net), 
            .I3(n32098), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_20 (.CI(n32098), .I0(n9094[17]), .I1(GND_net), 
            .CO(n32099));
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n9094[16]), .I2(GND_net), 
            .I3(n32097), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_19 (.CI(n32097), .I0(n9094[16]), .I1(GND_net), 
            .CO(n32098));
    SB_LUT4 mult_10_add_1225_6_lut (.I0(n26500), .I1(n8797[3]), .I2(n366), 
            .I3(n31841), .O(n2942[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n9094[15]), .I2(GND_net), 
            .I3(n32096), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_3669));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_3668));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_6 (.CI(n31841), .I0(n8797[3]), .I1(n366), 
            .CO(n31842));
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_3571));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[12]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_3665));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_18 (.CI(n32096), .I0(n9094[15]), .I1(GND_net), 
            .CO(n32097));
    SB_LUT4 mult_10_add_1225_5_lut (.I0(n26500), .I1(n8797[2]), .I2(n293), 
            .I3(n31840), .O(n2942[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n9094[14]), .I2(GND_net), 
            .I3(n32095), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_5 (.CI(n31840), .I0(n8797[2]), .I1(n293), 
            .CO(n31841));
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1_adj_3897[3]), .I3(n30457), .O(n7_adj_3687)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY mult_11_add_1225_17 (.CI(n32095), .I0(n9094[14]), .I1(GND_net), 
            .CO(n32096));
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n9094[13]), .I2(GND_net), 
            .I3(n32094), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_4_lut (.I0(n26500), .I1(n8797[1]), .I2(n220), 
            .I3(n31839), .O(n2942[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_4 (.CI(n31839), .I0(n8797[1]), .I1(n220), 
            .CO(n31840));
    SB_LUT4 mult_10_add_1225_3_lut (.I0(n26500), .I1(n8797[0]), .I2(n147), 
            .I3(n31838), .O(n2942[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_11_add_1225_16 (.CI(n32094), .I0(n9094[13]), .I1(GND_net), 
            .CO(n32095));
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_3664));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_3 (.CI(n31838), .I0(n8797[0]), .I1(n147), 
            .CO(n31839));
    SB_LUT4 mult_10_add_1225_2_lut (.I0(n26500), .I1(n5_adj_3689), .I2(n74), 
            .I3(GND_net), .O(n2942[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n9094[12]), .I2(GND_net), 
            .I3(n32093), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5_adj_3689), .I1(n74), 
            .CO(n31838));
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_11_add_1225_15 (.CI(n32093), .I0(n9094[12]), .I1(GND_net), 
            .CO(n32094));
    SB_LUT4 add_4580_23_lut (.I0(GND_net), .I1(n8821[20]), .I2(GND_net), 
            .I3(n31837), .O(n8797[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4580_22_lut (.I0(GND_net), .I1(n8821[19]), .I2(GND_net), 
            .I3(n31836), .O(n8797[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n9094[11]), .I2(GND_net), 
            .I3(n32092), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_3663));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_11_add_1225_14 (.CI(n32092), .I0(n9094[11]), .I1(GND_net), 
            .CO(n32093));
    SB_CARRY add_4580_22 (.CI(n31836), .I0(n8821[19]), .I1(GND_net), .CO(n31837));
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n9094[10]), .I2(GND_net), 
            .I3(n32091), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4580_21_lut (.I0(GND_net), .I1(n8821[18]), .I2(GND_net), 
            .I3(n31835), .O(n8797[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_13 (.CI(n32091), .I0(n9094[10]), .I1(GND_net), 
            .CO(n32092));
    SB_CARRY add_4580_21 (.CI(n31835), .I0(n8821[18]), .I1(GND_net), .CO(n31836));
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n9094[9]), .I2(GND_net), 
            .I3(n32090), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_12 (.CI(n32090), .I0(n9094[9]), .I1(GND_net), 
            .CO(n32091));
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[13]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[14]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n9094[8]), .I2(GND_net), 
            .I3(n32089), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4580_20_lut (.I0(GND_net), .I1(n8821[17]), .I2(GND_net), 
            .I3(n31834), .O(n8797[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4580_20 (.CI(n31834), .I0(n8821[17]), .I1(GND_net), .CO(n31835));
    SB_CARRY mult_11_add_1225_11 (.CI(n32089), .I0(n9094[8]), .I1(GND_net), 
            .CO(n32090));
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n9094[7]), .I2(GND_net), 
            .I3(n32088), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n32088), .I0(n9094[7]), .I1(GND_net), 
            .CO(n32089));
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n9094[6]), .I2(GND_net), 
            .I3(n32087), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4580_19_lut (.I0(GND_net), .I1(n8821[16]), .I2(GND_net), 
            .I3(n31833), .O(n8797[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_9 (.CI(n32087), .I0(n9094[6]), .I1(GND_net), 
            .CO(n32088));
    SB_CARRY add_4580_19 (.CI(n31833), .I0(n8821[16]), .I1(GND_net), .CO(n31834));
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n9094[5]), .I2(n512_adj_3690), 
            .I3(n32086), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4580_18_lut (.I0(GND_net), .I1(n8821[15]), .I2(GND_net), 
            .I3(n31832), .O(n8797[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_8 (.CI(n32086), .I0(n9094[5]), .I1(n512_adj_3690), 
            .CO(n32087));
    SB_CARRY add_4580_18 (.CI(n31832), .I0(n8821[15]), .I1(GND_net), .CO(n31833));
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n9094[4]), .I2(n439_adj_3691), 
            .I3(n32085), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4580_17_lut (.I0(GND_net), .I1(n8821[14]), .I2(GND_net), 
            .I3(n31831), .O(n8797[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4580_17 (.CI(n31831), .I0(n8821[14]), .I1(GND_net), .CO(n31832));
    SB_CARRY mult_11_add_1225_7 (.CI(n32085), .I0(n9094[4]), .I1(n439_adj_3691), 
            .CO(n32086));
    SB_LUT4 add_4580_16_lut (.I0(GND_net), .I1(n8821[13]), .I2(GND_net), 
            .I3(n31830), .O(n8797[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n9094[3]), .I2(n366_adj_3693), 
            .I3(n32084), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4580_16 (.CI(n31830), .I0(n8821[13]), .I1(GND_net), .CO(n31831));
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[15]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mult_11_add_1225_6 (.CI(n32084), .I0(n9094[3]), .I1(n366_adj_3693), 
            .CO(n32085));
    SB_LUT4 add_4580_15_lut (.I0(GND_net), .I1(n8821[12]), .I2(GND_net), 
            .I3(n31829), .O(n8797[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n9094[2]), .I2(n293_adj_3694), 
            .I3(n32083), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4580_15 (.CI(n31829), .I0(n8821[12]), .I1(GND_net), .CO(n31830));
    SB_CARRY unary_minus_5_add_3_5 (.CI(n30457), .I0(GND_net), .I1(n1_adj_3897[3]), 
            .CO(n30458));
    SB_LUT4 add_4580_14_lut (.I0(GND_net), .I1(n8821[11]), .I2(GND_net), 
            .I3(n31828), .O(n8797[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_5 (.CI(n32083), .I0(n9094[2]), .I1(n293_adj_3694), 
            .CO(n32084));
    SB_CARRY add_4580_14 (.CI(n31828), .I0(n8821[11]), .I1(GND_net), .CO(n31829));
    SB_LUT4 add_4580_13_lut (.I0(GND_net), .I1(n8821[10]), .I2(GND_net), 
            .I3(n31827), .O(n8797[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n9094[1]), .I2(n220_adj_3695), 
            .I3(n32082), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_4 (.CI(n32082), .I0(n9094[1]), .I1(n220_adj_3695), 
            .CO(n32083));
    SB_CARRY add_4580_13 (.CI(n31827), .I0(n8821[10]), .I1(GND_net), .CO(n31828));
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n9094[0]), .I2(n147_adj_3696), 
            .I3(n32081), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n32081), .I0(n9094[0]), .I1(n147_adj_3696), 
            .CO(n32082));
    SB_LUT4 add_4580_12_lut (.I0(GND_net), .I1(n8821[9]), .I2(GND_net), 
            .I3(n31826), .O(n8797[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[16]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_3697), .I2(n74_adj_3698), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[17]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[18]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[19]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[20]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[21]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_3570));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_3569));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_3640));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1_adj_3897[2]), .I3(n30456), .O(n5_adj_3699)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[22]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[23]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty[20]), .I1(n257[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_3701));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty[19]), .I1(n257[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_3702));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty[22]), .I1(n257[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_3703));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty[13]), .I1(n257[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_3704));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty[14]), .I1(n257[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_3705));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty[15]), .I1(n257[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_3706));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty[16]), .I1(n257[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_3707));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty[17]), .I1(n257[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_3708));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty[18]), .I1(n257[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_3709));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty[21]), .I1(n257[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_3710));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty[7]), .I1(n257[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_3711));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty[8]), .I1(n257[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_3712));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty[9]), .I1(n257[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_3713));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty[10]), .I1(n257[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_3714));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty[11]), .I1(n257[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_3715));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty[12]), .I1(n257[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_3716));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36205_4_lut (.I0(n21_adj_3714), .I1(n19_adj_3713), .I2(n17_adj_3712), 
            .I3(n9_adj_3717), .O(n43329));
    defparam i36205_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36193_4_lut (.I0(n27_adj_3704), .I1(n15_adj_3711), .I2(n13_adj_3718), 
            .I3(n11_adj_3719), .O(n43317));
    defparam i36193_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_3707), 
            .I3(GND_net), .O(n12_adj_3720));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_3718), 
            .I3(GND_net), .O(n10_adj_3721));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_3720), .I1(n257[17]), .I2(n35_adj_3708), 
            .I3(GND_net), .O(n30_adj_3722));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36936_4_lut (.I0(n13_adj_3718), .I1(n11_adj_3719), .I2(n9_adj_3717), 
            .I3(n43386), .O(n44061));
    defparam i36936_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i36928_4_lut (.I0(n19_adj_3713), .I1(n17_adj_3712), .I2(n15_adj_3711), 
            .I3(n44061), .O(n44053));
    defparam i36928_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i37771_4_lut (.I0(n25_adj_3716), .I1(n23_adj_3715), .I2(n21_adj_3714), 
            .I3(n44053), .O(n44896));
    defparam i37771_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i37298_4_lut (.I0(n31_adj_3706), .I1(n29_adj_3705), .I2(n27_adj_3704), 
            .I3(n44896), .O(n44423));
    defparam i37298_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i37887_4_lut (.I0(n37_adj_3709), .I1(n35_adj_3708), .I2(n33_adj_3707), 
            .I3(n44423), .O(n45012));
    defparam i37887_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_3710), 
            .I3(GND_net), .O(n16_adj_3723));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37526_3_lut (.I0(n6_adj_3724), .I1(n257[10]), .I2(n21_adj_3714), 
            .I3(GND_net), .O(n44651));   // verilog/motorControl.v(46[19:35])
    defparam i37526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37527_3_lut (.I0(n44651), .I1(n257[11]), .I2(n23_adj_3715), 
            .I3(GND_net), .O(n44652));   // verilog/motorControl.v(46[19:35])
    defparam i37527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_3712), 
            .I3(GND_net), .O(n8_adj_3725));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_3723), .I1(n257[22]), .I2(n45_adj_3703), 
            .I3(GND_net), .O(n24_adj_3726));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36143_4_lut (.I0(n43_adj_3710), .I1(n25_adj_3716), .I2(n23_adj_3715), 
            .I3(n43329), .O(n43267));
    defparam i36143_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37488_4_lut (.I0(n24_adj_3726), .I1(n8_adj_3725), .I2(n45_adj_3703), 
            .I3(n43263), .O(n44613));   // verilog/motorControl.v(46[19:35])
    defparam i37488_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36771_3_lut (.I0(n44652), .I1(n257[12]), .I2(n25_adj_3716), 
            .I3(GND_net), .O(n43896));   // verilog/motorControl.v(46[19:35])
    defparam i36771_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_3_lut (.I0(n42863), .I1(n257[1]), .I2(duty[1]), 
            .I3(GND_net), .O(n4_adj_3727));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i37516_3_lut (.I0(n4_adj_3727), .I1(n257[13]), .I2(n27_adj_3704), 
            .I3(GND_net), .O(n44641));   // verilog/motorControl.v(46[19:35])
    defparam i37516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37517_3_lut (.I0(n44641), .I1(n257[14]), .I2(n29_adj_3705), 
            .I3(GND_net), .O(n44642));   // verilog/motorControl.v(46[19:35])
    defparam i37517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36179_4_lut (.I0(n33_adj_3707), .I1(n31_adj_3706), .I2(n29_adj_3705), 
            .I3(n43317), .O(n43303));
    defparam i36179_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37837_4_lut (.I0(n30_adj_3722), .I1(n10_adj_3721), .I2(n35_adj_3708), 
            .I3(n43293), .O(n44962));   // verilog/motorControl.v(46[19:35])
    defparam i37837_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36773_3_lut (.I0(n44642), .I1(n257[15]), .I2(n31_adj_3706), 
            .I3(GND_net), .O(n43898));   // verilog/motorControl.v(46[19:35])
    defparam i36773_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37967_4_lut (.I0(n43898), .I1(n44962), .I2(n35_adj_3708), 
            .I3(n43303), .O(n45092));   // verilog/motorControl.v(46[19:35])
    defparam i37967_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i37968_3_lut (.I0(n45092), .I1(n257[18]), .I2(n37_adj_3709), 
            .I3(GND_net), .O(n45093));   // verilog/motorControl.v(46[19:35])
    defparam i37968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37933_3_lut (.I0(n45093), .I1(n257[19]), .I2(n39_adj_3702), 
            .I3(GND_net), .O(n45058));   // verilog/motorControl.v(46[19:35])
    defparam i37933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36147_4_lut (.I0(n43_adj_3710), .I1(n41_adj_3701), .I2(n39_adj_3702), 
            .I3(n45012), .O(n43271));
    defparam i36147_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37707_4_lut (.I0(n43896), .I1(n44613), .I2(n45_adj_3703), 
            .I3(n43267), .O(n44832));   // verilog/motorControl.v(46[19:35])
    defparam i37707_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36779_3_lut (.I0(n45058), .I1(n257[20]), .I2(n41_adj_3701), 
            .I3(GND_net), .O(n43904));   // verilog/motorControl.v(46[19:35])
    defparam i36779_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37869_4_lut (.I0(n43904), .I1(n44832), .I2(n45_adj_3703), 
            .I3(n43271), .O(n44994));   // verilog/motorControl.v(46[19:35])
    defparam i37869_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i37870_3_lut (.I0(n44994), .I1(duty[23]), .I2(n47), .I3(GND_net), 
            .O(n256));   // verilog/motorControl.v(46[19:35])
    defparam i37870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_626_i3_3_lut (.I0(n155[2]), .I1(PWMLimit[2]), .I2(n256), 
            .I3(GND_net), .O(n2967[2]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21516_2_lut_2_lut (.I0(n256), .I1(n7831[0]), .I2(GND_net), 
            .I3(GND_net), .O(n2942[23]));   // verilog/motorControl.v(46[19:35])
    defparam i21516_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[0]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4580_12 (.CI(n31826), .I0(n8821[9]), .I1(GND_net), .CO(n31827));
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_3697), .I1(n74_adj_3698), 
            .CO(n32081));
    SB_LUT4 add_4580_11_lut (.I0(GND_net), .I1(n8821[8]), .I2(GND_net), 
            .I3(n31825), .O(n8797[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36420_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty[3]), .I2(duty[2]), 
            .I3(PWMLimit[2]), .O(n43545));   // verilog/motorControl.v(44[10:25])
    defparam i36420_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_4602_23_lut (.I0(GND_net), .I1(n9118[20]), .I2(GND_net), 
            .I3(n32080), .O(n9094[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4580_11 (.CI(n31825), .I0(n8821[8]), .I1(GND_net), .CO(n31826));
    SB_LUT4 add_4602_22_lut (.I0(GND_net), .I1(n9118[19]), .I2(GND_net), 
            .I3(n32079), .O(n9094[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4580_10_lut (.I0(GND_net), .I1(n8821[7]), .I2(GND_net), 
            .I3(n31824), .O(n8797[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_22 (.CI(n32079), .I0(n9118[19]), .I1(GND_net), .CO(n32080));
    SB_CARRY add_4580_10 (.CI(n31824), .I0(n8821[7]), .I1(GND_net), .CO(n31825));
    SB_LUT4 add_4602_21_lut (.I0(GND_net), .I1(n9118[18]), .I2(GND_net), 
            .I3(n32078), .O(n9094[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4580_9_lut (.I0(GND_net), .I1(n8821[6]), .I2(GND_net), 
            .I3(n31823), .O(n8797[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_21 (.CI(n32078), .I0(n9118[18]), .I1(GND_net), .CO(n32079));
    SB_CARRY add_4580_9 (.CI(n31823), .I0(n8821[6]), .I1(GND_net), .CO(n31824));
    SB_LUT4 add_4602_20_lut (.I0(GND_net), .I1(n9118[17]), .I2(GND_net), 
            .I3(n32077), .O(n9094[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty[3]), 
            .I2(duty[2]), .I3(GND_net), .O(n6_adj_3622));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 add_4580_8_lut (.I0(GND_net), .I1(n8821[5]), .I2(n515_adj_3729), 
            .I3(n31822), .O(n8797[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_20 (.CI(n32077), .I0(n9118[17]), .I1(GND_net), .CO(n32078));
    SB_CARRY add_4580_8 (.CI(n31822), .I0(n8821[5]), .I1(n515_adj_3729), 
            .CO(n31823));
    SB_LUT4 add_4602_19_lut (.I0(GND_net), .I1(n9118[16]), .I2(GND_net), 
            .I3(n32076), .O(n9094[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4580_7_lut (.I0(GND_net), .I1(n8821[4]), .I2(n442_adj_3730), 
            .I3(n31821), .O(n8797[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_19 (.CI(n32076), .I0(n9118[16]), .I1(GND_net), .CO(n32077));
    SB_CARRY add_4580_7 (.CI(n31821), .I0(n8821[4]), .I1(n442_adj_3730), 
            .CO(n31822));
    SB_LUT4 add_4602_18_lut (.I0(GND_net), .I1(n9118[15]), .I2(GND_net), 
            .I3(n32075), .O(n9094[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4580_6_lut (.I0(GND_net), .I1(n8821[3]), .I2(n369_adj_3731), 
            .I3(n31820), .O(n8797[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_18 (.CI(n32075), .I0(n9118[15]), .I1(GND_net), .CO(n32076));
    SB_CARRY add_4580_6 (.CI(n31820), .I0(n8821[3]), .I1(n369_adj_3731), 
            .CO(n31821));
    SB_LUT4 add_4602_17_lut (.I0(GND_net), .I1(n9118[14]), .I2(GND_net), 
            .I3(n32074), .O(n9094[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_17 (.CI(n32074), .I0(n9118[14]), .I1(GND_net), .CO(n32075));
    SB_LUT4 add_4580_5_lut (.I0(GND_net), .I1(n8821[2]), .I2(n296_adj_3732), 
            .I3(n31819), .O(n8797[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4580_5 (.CI(n31819), .I0(n8821[2]), .I1(n296_adj_3732), 
            .CO(n31820));
    SB_LUT4 add_4580_4_lut (.I0(GND_net), .I1(n8821[1]), .I2(n223_adj_3733), 
            .I3(n31818), .O(n8797[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4602_16_lut (.I0(GND_net), .I1(n9118[13]), .I2(GND_net), 
            .I3(n32073), .O(n9094[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4580_4 (.CI(n31818), .I0(n8821[1]), .I1(n223_adj_3733), 
            .CO(n31819));
    SB_CARRY add_4602_16 (.CI(n32073), .I0(n9118[13]), .I1(GND_net), .CO(n32074));
    SB_CARRY unary_minus_5_add_3_4 (.CI(n30456), .I0(GND_net), .I1(n1_adj_3897[2]), 
            .CO(n30457));
    SB_LUT4 add_4580_3_lut (.I0(GND_net), .I1(n8821[0]), .I2(n150_adj_3734), 
            .I3(n31817), .O(n8797[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4580_3 (.CI(n31817), .I0(n8821[0]), .I1(n150_adj_3734), 
            .CO(n31818));
    SB_LUT4 add_4602_15_lut (.I0(GND_net), .I1(n9118[12]), .I2(GND_net), 
            .I3(n32072), .O(n9094[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4580_2_lut (.I0(GND_net), .I1(n8_adj_3735), .I2(n77_adj_3736), 
            .I3(GND_net), .O(n8797[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4580_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_15 (.CI(n32072), .I0(n9118[12]), .I1(GND_net), .CO(n32073));
    SB_LUT4 add_4602_14_lut (.I0(GND_net), .I1(n9118[11]), .I2(GND_net), 
            .I3(n32071), .O(n9094[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_14 (.CI(n32071), .I0(n9118[11]), .I1(GND_net), .CO(n32072));
    SB_CARRY add_4580_2 (.CI(GND_net), .I0(n8_adj_3735), .I1(n77_adj_3736), 
            .CO(n31817));
    SB_LUT4 add_4618_7_lut (.I0(GND_net), .I1(n38956), .I2(n490), .I3(n32302), 
            .O(n9358[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4618_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4602_13_lut (.I0(GND_net), .I1(n9118[10]), .I2(GND_net), 
            .I3(n32070), .O(n9094[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_13 (.CI(n32070), .I0(n9118[10]), .I1(GND_net), .CO(n32071));
    SB_LUT4 add_4618_6_lut (.I0(GND_net), .I1(n9366[3]), .I2(n417), .I3(n32301), 
            .O(n9358[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4618_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4602_12_lut (.I0(GND_net), .I1(n9118[9]), .I2(GND_net), 
            .I3(n32069), .O(n9094[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4618_6 (.CI(n32301), .I0(n9366[3]), .I1(n417), .CO(n32302));
    SB_CARRY add_4602_12 (.CI(n32069), .I0(n9118[9]), .I1(GND_net), .CO(n32070));
    SB_LUT4 add_4618_5_lut (.I0(GND_net), .I1(n9366[2]), .I2(n344), .I3(n32300), 
            .O(n9358[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4618_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4602_11_lut (.I0(GND_net), .I1(n9118[8]), .I2(GND_net), 
            .I3(n32068), .O(n9094[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4618_5 (.CI(n32300), .I0(n9366[2]), .I1(n344), .CO(n32301));
    SB_CARRY add_4602_11 (.CI(n32068), .I0(n9118[8]), .I1(GND_net), .CO(n32069));
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1_adj_3897[1]), .I3(n30455), .O(n3_adj_3737)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_3 (.CI(n30455), .I0(GND_net), .I1(n1_adj_3897[1]), 
            .CO(n30456));
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_3897[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3454 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_3897[0]), 
            .CO(n30455));
    SB_LUT4 add_4618_4_lut (.I0(GND_net), .I1(n9366[1]), .I2(n271_adj_3686), 
            .I3(n32299), .O(n9358[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4618_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4602_10_lut (.I0(GND_net), .I1(n9118[7]), .I2(GND_net), 
            .I3(n32067), .O(n9094[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_10 (.CI(n32067), .I0(n9118[7]), .I1(GND_net), .CO(n32068));
    SB_CARRY add_4618_4 (.CI(n32299), .I0(n9366[1]), .I1(n271_adj_3686), 
            .CO(n32300));
    SB_LUT4 add_4602_9_lut (.I0(GND_net), .I1(n9118[6]), .I2(GND_net), 
            .I3(n32066), .O(n9094[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4618_3_lut (.I0(GND_net), .I1(n9366[0]), .I2(n198), .I3(n32298), 
            .O(n9358[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4618_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_9 (.CI(n32066), .I0(n9118[6]), .I1(GND_net), .CO(n32067));
    SB_CARRY add_4618_3 (.CI(n32298), .I0(n9366[0]), .I1(n198), .CO(n32299));
    SB_LUT4 add_4602_8_lut (.I0(GND_net), .I1(n9118[5]), .I2(n515), .I3(n32065), 
            .O(n9094[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4618_2_lut (.I0(GND_net), .I1(n56), .I2(n125_adj_3685), 
            .I3(GND_net), .O(n9358[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4618_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_8 (.CI(n32065), .I0(n9118[5]), .I1(n515), .CO(n32066));
    SB_CARRY add_4618_2 (.CI(GND_net), .I0(n56), .I1(n125_adj_3685), .CO(n32298));
    SB_LUT4 add_4602_7_lut (.I0(GND_net), .I1(n9118[4]), .I2(n442), .I3(n32064), 
            .O(n9094[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4617_8_lut (.I0(GND_net), .I1(n9358[5]), .I2(n560), .I3(n32297), 
            .O(n9349[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4617_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_7 (.CI(n32064), .I0(n9118[4]), .I1(n442), .CO(n32065));
    SB_LUT4 add_4602_6_lut (.I0(GND_net), .I1(n9118[3]), .I2(n369), .I3(n32063), 
            .O(n9094[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4617_7_lut (.I0(GND_net), .I1(n9358[4]), .I2(n487), .I3(n32296), 
            .O(n9349[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4617_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4617_7 (.CI(n32296), .I0(n9358[4]), .I1(n487), .CO(n32297));
    SB_CARRY add_4602_6 (.CI(n32063), .I0(n9118[3]), .I1(n369), .CO(n32064));
    SB_LUT4 add_4602_5_lut (.I0(GND_net), .I1(n9118[2]), .I2(n296), .I3(n32062), 
            .O(n9094[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_5 (.CI(n32062), .I0(n9118[2]), .I1(n296), .CO(n32063));
    SB_LUT4 add_4602_4_lut (.I0(GND_net), .I1(n9118[1]), .I2(n223), .I3(n32061), 
            .O(n9094[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_4 (.CI(n32061), .I0(n9118[1]), .I1(n223), .CO(n32062));
    SB_LUT4 add_4602_3_lut (.I0(GND_net), .I1(n9118[0]), .I2(n150), .I3(n32060), 
            .O(n9094[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4602_3 (.CI(n32060), .I0(n9118[0]), .I1(n150), .CO(n32061));
    SB_LUT4 add_4602_2_lut (.I0(GND_net), .I1(n8_adj_3592), .I2(n77), 
            .I3(GND_net), .O(n9094[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4602_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4617_6_lut (.I0(GND_net), .I1(n9358[3]), .I2(n414), .I3(n32295), 
            .O(n9349[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4617_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4617_6 (.CI(n32295), .I0(n9358[3]), .I1(n414), .CO(n32296));
    SB_LUT4 add_4617_5_lut (.I0(GND_net), .I1(n9358[2]), .I2(n341), .I3(n32294), 
            .O(n9349[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4617_5_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3355[1]));   // verilog/motorControl.v(37[14] 56[8])
    SB_CARRY add_4602_2 (.CI(GND_net), .I0(n8_adj_3592), .I1(n77), .CO(n32060));
    SB_CARRY add_4617_5 (.CI(n32294), .I0(n9358[2]), .I1(n341), .CO(n32295));
    SB_LUT4 add_4596_7_lut (.I0(GND_net), .I1(n39599), .I2(n490_adj_3739), 
            .I3(n32059), .O(n9061[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4596_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4617_4_lut (.I0(GND_net), .I1(n9358[1]), .I2(n268_adj_3740), 
            .I3(n32293), .O(n9349[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4617_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4617_4 (.CI(n32293), .I0(n9358[1]), .I1(n268_adj_3740), 
            .CO(n32294));
    SB_LUT4 add_4617_3_lut (.I0(GND_net), .I1(n9358[0]), .I2(n195_adj_3741), 
            .I3(n32292), .O(n9349[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4617_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4617_3 (.CI(n32292), .I0(n9358[0]), .I1(n195_adj_3741), 
            .CO(n32293));
    SB_LUT4 add_4596_6_lut (.I0(GND_net), .I1(n9069[3]), .I2(n417_adj_3742), 
            .I3(n32058), .O(n9061[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4596_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4596_6 (.CI(n32058), .I0(n9069[3]), .I1(n417_adj_3742), 
            .CO(n32059));
    SB_LUT4 add_4617_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n9349[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4617_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4596_5_lut (.I0(GND_net), .I1(n9069[2]), .I2(n344_adj_3743), 
            .I3(n32057), .O(n9061[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4596_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4617_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n32292));
    SB_CARRY add_4596_5 (.CI(n32057), .I0(n9069[2]), .I1(n344_adj_3743), 
            .CO(n32058));
    SB_LUT4 add_4596_4_lut (.I0(GND_net), .I1(n9069[1]), .I2(n271_adj_3744), 
            .I3(n32056), .O(n9061[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4596_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4616_9_lut (.I0(GND_net), .I1(n9349[6]), .I2(GND_net), 
            .I3(n32291), .O(n9339[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4616_8_lut (.I0(GND_net), .I1(n9349[5]), .I2(n557), .I3(n32290), 
            .O(n9339[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4596_4 (.CI(n32056), .I0(n9069[1]), .I1(n271_adj_3744), 
            .CO(n32057));
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[1]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_4616_8 (.CI(n32290), .I0(n9349[5]), .I1(n557), .CO(n32291));
    SB_LUT4 add_4596_3_lut (.I0(GND_net), .I1(n9069[0]), .I2(n198_adj_3745), 
            .I3(n32055), .O(n9061[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4596_3_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3355[2]));   // verilog/motorControl.v(37[14] 56[8])
    SB_LUT4 add_4616_7_lut (.I0(GND_net), .I1(n9349[4]), .I2(n484), .I3(n32289), 
            .O(n9339[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3355[3]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3355[4]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3355[5]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3355[6]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3355[7]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3355[8]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3355[9]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3355[10]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3355[11]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3355[12]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3355[13]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3355[14]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3355[15]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3355[16]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3355[17]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3355[18]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3355[19]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3355[20]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3355[21]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3355[22]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3355[23]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i1  (.Q(\PID_CONTROLLER.err [1]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [1]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i2  (.Q(\PID_CONTROLLER.err [2]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [2]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i3  (.Q(\PID_CONTROLLER.err [3]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [3]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i4  (.Q(\PID_CONTROLLER.err [4]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [4]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i5  (.Q(\PID_CONTROLLER.err [5]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [5]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i6  (.Q(\PID_CONTROLLER.err [6]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [6]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i7  (.Q(\PID_CONTROLLER.err [7]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [7]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i8  (.Q(\PID_CONTROLLER.err [8]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [8]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i9  (.Q(\PID_CONTROLLER.err [9]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [9]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i10  (.Q(\PID_CONTROLLER.err [10]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [10]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i11  (.Q(\PID_CONTROLLER.err [11]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [11]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i12  (.Q(\PID_CONTROLLER.err [12]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [12]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i13  (.Q(\PID_CONTROLLER.err [13]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [13]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i14  (.Q(\PID_CONTROLLER.err [14]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [14]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i15  (.Q(\PID_CONTROLLER.err [15]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [15]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i16  (.Q(\PID_CONTROLLER.err [16]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [16]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i17  (.Q(\PID_CONTROLLER.err [17]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [17]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i18  (.Q(\PID_CONTROLLER.err [18]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [18]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i19  (.Q(\PID_CONTROLLER.err [19]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [19]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i20  (.Q(\PID_CONTROLLER.err [20]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [20]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i21  (.Q(\PID_CONTROLLER.err [21]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [21]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i22  (.Q(\PID_CONTROLLER.err [22]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [22]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i23  (.Q(\PID_CONTROLLER.err [23]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3379 [23]));   // verilog/motorControl.v(37[14] 56[8])
    SB_CARRY add_4596_3 (.CI(n32055), .I0(n9069[0]), .I1(n198_adj_3745), 
            .CO(n32056));
    SB_CARRY add_4616_7 (.CI(n32289), .I0(n9349[4]), .I1(n484), .CO(n32290));
    SB_LUT4 add_4596_2_lut (.I0(GND_net), .I1(n56_adj_3746), .I2(n125_adj_3747), 
            .I3(GND_net), .O(n9061[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4596_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4616_6_lut (.I0(GND_net), .I1(n9349[3]), .I2(n411), .I3(n32288), 
            .O(n9339[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4596_2 (.CI(GND_net), .I0(n56_adj_3746), .I1(n125_adj_3747), 
            .CO(n32055));
    SB_CARRY add_4616_6 (.CI(n32288), .I0(n9349[3]), .I1(n411), .CO(n32289));
    SB_LUT4 add_4595_8_lut (.I0(GND_net), .I1(n9061[5]), .I2(n560_adj_3748), 
            .I3(n32054), .O(n9052[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4616_5_lut (.I0(GND_net), .I1(n9349[2]), .I2(n338), .I3(n32287), 
            .O(n9339[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4595_7_lut (.I0(GND_net), .I1(n9061[4]), .I2(n487_adj_3749), 
            .I3(n32053), .O(n9052[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4616_5 (.CI(n32287), .I0(n9349[2]), .I1(n338), .CO(n32288));
    SB_CARRY add_4595_7 (.CI(n32053), .I0(n9061[4]), .I1(n487_adj_3749), 
            .CO(n32054));
    SB_LUT4 add_4616_4_lut (.I0(GND_net), .I1(n9349[1]), .I2(n265_adj_3750), 
            .I3(n32286), .O(n9339[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4595_6_lut (.I0(GND_net), .I1(n9061[3]), .I2(n414_adj_3751), 
            .I3(n32052), .O(n9052[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4595_6 (.CI(n32052), .I0(n9061[3]), .I1(n414_adj_3751), 
            .CO(n32053));
    SB_LUT4 add_4595_5_lut (.I0(GND_net), .I1(n9061[2]), .I2(n341_adj_3752), 
            .I3(n32051), .O(n9052[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4616_4 (.CI(n32286), .I0(n9349[1]), .I1(n265_adj_3750), 
            .CO(n32287));
    SB_CARRY add_4595_5 (.CI(n32051), .I0(n9061[2]), .I1(n341_adj_3752), 
            .CO(n32052));
    SB_LUT4 add_4616_3_lut (.I0(GND_net), .I1(n9349[0]), .I2(n192_adj_3753), 
            .I3(n32285), .O(n9339[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4595_4_lut (.I0(GND_net), .I1(n9061[1]), .I2(n268_adj_3754), 
            .I3(n32050), .O(n9052[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4595_4 (.CI(n32050), .I0(n9061[1]), .I1(n268_adj_3754), 
            .CO(n32051));
    SB_CARRY add_4616_3 (.CI(n32285), .I0(n9349[0]), .I1(n192_adj_3753), 
            .CO(n32286));
    SB_LUT4 add_4595_3_lut (.I0(GND_net), .I1(n9061[0]), .I2(n195_adj_3755), 
            .I3(n32049), .O(n9052[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4595_3 (.CI(n32049), .I0(n9061[0]), .I1(n195_adj_3755), 
            .CO(n32050));
    SB_LUT4 add_4616_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n9339[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4616_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4595_2_lut (.I0(GND_net), .I1(n53_adj_3756), .I2(n122_adj_3757), 
            .I3(GND_net), .O(n9052[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4595_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4616_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n32285));
    SB_CARRY add_4595_2 (.CI(GND_net), .I0(n53_adj_3756), .I1(n122_adj_3757), 
            .CO(n32049));
    SB_LUT4 add_4615_10_lut (.I0(GND_net), .I1(n9339[7]), .I2(GND_net), 
            .I3(n32284), .O(n9328[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4615_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4615_9_lut (.I0(GND_net), .I1(n9339[6]), .I2(GND_net), 
            .I3(n32283), .O(n9328[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4615_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4615_9 (.CI(n32283), .I0(n9339[6]), .I1(GND_net), .CO(n32284));
    SB_LUT4 i25190_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n4_adj_3758), .I3(n9373[1]), .O(n6_adj_3759));   // verilog/motorControl.v(42[26:37])
    defparam i25190_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n9373[1]), .I3(n4_adj_3758), .O(n9366[2]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_846 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n9373[0]), .I3(n30129), .O(n9366[1]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut_adj_846.LUT_INIT = 16'h8778;
    SB_LUT4 i25182_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n30129), .I3(n9373[0]), .O(n4_adj_3758));   // verilog/motorControl.v(42[26:37])
    defparam i25182_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i25171_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(\Ki[1] ), .O(n30129));   // verilog/motorControl.v(42[26:37])
    defparam i25171_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i25169_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(\Ki[1] ), .O(n9366[0]));   // verilog/motorControl.v(42[26:37])
    defparam i25169_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_4615_8_lut (.I0(GND_net), .I1(n9339[5]), .I2(n554), .I3(n32282), 
            .O(n9328[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4615_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4615_8 (.CI(n32282), .I0(n9339[5]), .I1(n554), .CO(n32283));
    SB_LUT4 add_4615_7_lut (.I0(GND_net), .I1(n9339[4]), .I2(n481), .I3(n32281), 
            .O(n9328[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4615_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4594_9_lut (.I0(GND_net), .I1(n9052[6]), .I2(GND_net), 
            .I3(n32048), .O(n9042[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4594_8_lut (.I0(GND_net), .I1(n9052[5]), .I2(n557_adj_3760), 
            .I3(n32047), .O(n9042[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_8 (.CI(n32047), .I0(n9052[5]), .I1(n557_adj_3760), 
            .CO(n32048));
    SB_LUT4 add_4594_7_lut (.I0(GND_net), .I1(n9052[4]), .I2(n484_adj_3761), 
            .I3(n32046), .O(n9042[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4615_7 (.CI(n32281), .I0(n9339[4]), .I1(n481), .CO(n32282));
    SB_CARRY add_4594_7 (.CI(n32046), .I0(n9052[4]), .I1(n484_adj_3761), 
            .CO(n32047));
    SB_LUT4 add_4594_6_lut (.I0(GND_net), .I1(n9052[3]), .I2(n411_adj_3762), 
            .I3(n32045), .O(n9042[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25252_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n30206), .I3(n9384[0]), .O(n4_adj_3763));   // verilog/motorControl.v(42[26:37])
    defparam i25252_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_847 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n9384[0]), .I3(n30206), .O(n9379[1]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut_adj_847.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_848 (.I0(n62), .I1(n131), .I2(n9379[0]), 
            .I3(n204), .O(n9373[1]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut_adj_848.LUT_INIT = 16'h8778;
    SB_LUT4 i25221_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n9379[0]), 
            .O(n4_adj_3764));   // verilog/motorControl.v(42[26:37])
    defparam i25221_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i25241_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(\Ki[1] ), .O(n30206));   // verilog/motorControl.v(42[26:37])
    defparam i25241_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i25239_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(\Ki[1] ), .O(n9379[0]));   // verilog/motorControl.v(42[26:37])
    defparam i25239_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_4615_6_lut (.I0(GND_net), .I1(n9339[3]), .I2(n408), .I3(n32280), 
            .O(n9328[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4615_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_6 (.CI(n32045), .I0(n9052[3]), .I1(n411_adj_3762), 
            .CO(n32046));
    SB_CARRY add_4615_6 (.CI(n32280), .I0(n9339[3]), .I1(n408), .CO(n32281));
    SB_LUT4 add_4594_5_lut (.I0(GND_net), .I1(n9052[2]), .I2(n338_adj_3765), 
            .I3(n32044), .O(n9042[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4615_5_lut (.I0(GND_net), .I1(n9339[2]), .I2(n335), .I3(n32279), 
            .O(n9328[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4615_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_5 (.CI(n32044), .I0(n9052[2]), .I1(n338_adj_3765), 
            .CO(n32045));
    SB_CARRY add_4615_5 (.CI(n32279), .I0(n9339[2]), .I1(n335), .CO(n32280));
    SB_LUT4 add_4594_4_lut (.I0(GND_net), .I1(n9052[1]), .I2(n265_adj_3766), 
            .I3(n32043), .O(n9042[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4615_4_lut (.I0(GND_net), .I1(n9339[1]), .I2(n262_adj_3767), 
            .I3(n32278), .O(n9328[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4615_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_4 (.CI(n32043), .I0(n9052[1]), .I1(n265_adj_3766), 
            .CO(n32044));
    SB_CARRY add_4615_4 (.CI(n32278), .I0(n9339[1]), .I1(n262_adj_3767), 
            .CO(n32279));
    SB_LUT4 add_4594_3_lut (.I0(GND_net), .I1(n9052[0]), .I2(n192_adj_3768), 
            .I3(n32042), .O(n9042[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4615_3_lut (.I0(GND_net), .I1(n9339[0]), .I2(n189_adj_3769), 
            .I3(n32277), .O(n9328[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4615_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_3 (.CI(n32042), .I0(n9052[0]), .I1(n192_adj_3768), 
            .CO(n32043));
    SB_LUT4 add_4594_2_lut (.I0(GND_net), .I1(n50_adj_3770), .I2(n119_adj_3771), 
            .I3(GND_net), .O(n9042[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4594_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4615_3 (.CI(n32277), .I0(n9339[0]), .I1(n189_adj_3769), 
            .CO(n32278));
    SB_LUT4 add_4615_2_lut (.I0(GND_net), .I1(n47_adj_3772), .I2(n116), 
            .I3(GND_net), .O(n9328[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4615_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4594_2 (.CI(GND_net), .I0(n50_adj_3770), .I1(n119_adj_3771), 
            .CO(n32042));
    SB_CARRY add_4615_2 (.CI(GND_net), .I0(n47_adj_3772), .I1(n116), .CO(n32277));
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4593_10_lut (.I0(GND_net), .I1(n9042[7]), .I2(GND_net), 
            .I3(n32041), .O(n9031[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4593_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4614_11_lut (.I0(GND_net), .I1(n9328[8]), .I2(GND_net), 
            .I3(n32276), .O(n9316[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4614_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4593_9_lut (.I0(GND_net), .I1(n9042[6]), .I2(GND_net), 
            .I3(n32040), .O(n9031[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4593_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4593_9 (.CI(n32040), .I0(n9042[6]), .I1(GND_net), .CO(n32041));
    SB_LUT4 add_4614_10_lut (.I0(GND_net), .I1(n9328[7]), .I2(GND_net), 
            .I3(n32275), .O(n9316[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4614_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4593_8_lut (.I0(GND_net), .I1(n9042[5]), .I2(n554_adj_3773), 
            .I3(n32039), .O(n9031[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4593_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4614_10 (.CI(n32275), .I0(n9328[7]), .I1(GND_net), .CO(n32276));
    SB_CARRY add_4593_8 (.CI(n32039), .I0(n9042[5]), .I1(n554_adj_3773), 
            .CO(n32040));
    SB_LUT4 add_4614_9_lut (.I0(GND_net), .I1(n9328[6]), .I2(GND_net), 
            .I3(n32274), .O(n9316[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4614_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4593_7_lut (.I0(GND_net), .I1(n9042[4]), .I2(n481_adj_3774), 
            .I3(n32038), .O(n9031[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4593_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4614_9 (.CI(n32274), .I0(n9328[6]), .I1(GND_net), .CO(n32275));
    SB_CARRY add_4593_7 (.CI(n32038), .I0(n9042[4]), .I1(n481_adj_3774), 
            .CO(n32039));
    SB_LUT4 state_23__I_0_add_2_25_lut (.I0(GND_net), .I1(motor_state[23]), 
            .I2(n1_adj_3898[23]), .I3(n30523), .O(\PID_CONTROLLER.err_23__N_3379 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4614_8_lut (.I0(GND_net), .I1(n9328[5]), .I2(n551), .I3(n32273), 
            .O(n9316[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4614_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4593_6_lut (.I0(GND_net), .I1(n9042[3]), .I2(n408_adj_3776), 
            .I3(n32037), .O(n9031[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4593_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4593_6 (.CI(n32037), .I0(n9042[3]), .I1(n408_adj_3776), 
            .CO(n32038));
    SB_CARRY add_4614_8 (.CI(n32273), .I0(n9328[5]), .I1(n551), .CO(n32274));
    SB_LUT4 add_4593_5_lut (.I0(GND_net), .I1(n9042[2]), .I2(n335_adj_3777), 
            .I3(n32036), .O(n9031[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4593_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4593_5 (.CI(n32036), .I0(n9042[2]), .I1(n335_adj_3777), 
            .CO(n32037));
    SB_LUT4 add_4614_7_lut (.I0(GND_net), .I1(n9328[4]), .I2(n478), .I3(n32272), 
            .O(n9316[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4614_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4593_4_lut (.I0(GND_net), .I1(n9042[1]), .I2(n262_adj_3778), 
            .I3(n32035), .O(n9031[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4593_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4593_4 (.CI(n32035), .I0(n9042[1]), .I1(n262_adj_3778), 
            .CO(n32036));
    SB_CARRY add_4614_7 (.CI(n32272), .I0(n9328[4]), .I1(n478), .CO(n32273));
    SB_LUT4 add_4593_3_lut (.I0(GND_net), .I1(n9042[0]), .I2(n189_adj_3779), 
            .I3(n32034), .O(n9031[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4593_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4614_6_lut (.I0(GND_net), .I1(n9328[3]), .I2(n405), .I3(n32271), 
            .O(n9316[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4614_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4614_6 (.CI(n32271), .I0(n9328[3]), .I1(n405), .CO(n32272));
    SB_LUT4 add_4614_5_lut (.I0(GND_net), .I1(n9328[2]), .I2(n332), .I3(n32270), 
            .O(n9316[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4614_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4614_5 (.CI(n32270), .I0(n9328[2]), .I1(n332), .CO(n32271));
    SB_LUT4 add_4614_4_lut (.I0(GND_net), .I1(n9328[1]), .I2(n259_adj_3780), 
            .I3(n32269), .O(n9316[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4614_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4614_4 (.CI(n32269), .I0(n9328[1]), .I1(n259_adj_3780), 
            .CO(n32270));
    SB_CARRY add_4593_3 (.CI(n32034), .I0(n9042[0]), .I1(n189_adj_3779), 
            .CO(n32035));
    SB_LUT4 state_23__I_0_add_2_24_lut (.I0(GND_net), .I1(motor_state[22]), 
            .I2(n1_adj_3898[22]), .I3(n30522), .O(\PID_CONTROLLER.err_23__N_3379 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4593_2_lut (.I0(GND_net), .I1(n47_adj_3782), .I2(n116_adj_3783), 
            .I3(GND_net), .O(n9031[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4593_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4614_3_lut (.I0(GND_net), .I1(n9328[0]), .I2(n186_adj_3784), 
            .I3(n32268), .O(n9316[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4614_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4614_3 (.CI(n32268), .I0(n9328[0]), .I1(n186_adj_3784), 
            .CO(n32269));
    SB_CARRY add_4593_2 (.CI(GND_net), .I0(n47_adj_3782), .I1(n116_adj_3783), 
            .CO(n32034));
    SB_LUT4 add_4592_11_lut (.I0(GND_net), .I1(n9031[8]), .I2(GND_net), 
            .I3(n32033), .O(n9019[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4592_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4614_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n9316[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4614_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_24 (.CI(n30522), .I0(motor_state[22]), 
            .I1(n1_adj_3898[22]), .CO(n30523));
    SB_LUT4 add_4592_10_lut (.I0(GND_net), .I1(n9031[7]), .I2(GND_net), 
            .I3(n32032), .O(n9019[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4592_10_lut.LUT_INIT = 16'hC33C;
    SB_DFFE \PID_CONTROLLER.integral_1149__i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[1]));   // verilog/motorControl.v(40[21:33])
    SB_LUT4 state_23__I_0_add_2_23_lut (.I0(GND_net), .I1(motor_state[21]), 
            .I2(n1_adj_3898[21]), .I3(n30521), .O(\PID_CONTROLLER.err_23__N_3379 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_23 (.CI(n30521), .I0(motor_state[21]), 
            .I1(n1_adj_3898[21]), .CO(n30522));
    SB_DFFE \PID_CONTROLLER.integral_1149__i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[2]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[3]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[4]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[5]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[6]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[7]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[8]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[9]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[10]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[11]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[12]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[13]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[14]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[15]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[16]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[17]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[18]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[19]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[20]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[21]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[22]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1149__i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3451 ), .D(n34[23]));   // verilog/motorControl.v(40[21:33])
    SB_CARRY add_4614_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n32268));
    SB_CARRY add_4592_10 (.CI(n32032), .I0(n9031[7]), .I1(GND_net), .CO(n32033));
    SB_LUT4 add_4613_12_lut (.I0(GND_net), .I1(n9316[9]), .I2(GND_net), 
            .I3(n32267), .O(n9303[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4613_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4592_9_lut (.I0(GND_net), .I1(n9031[6]), .I2(GND_net), 
            .I3(n32031), .O(n9019[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4592_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4613_11_lut (.I0(GND_net), .I1(n9316[8]), .I2(GND_net), 
            .I3(n32266), .O(n9303[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4613_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4592_9 (.CI(n32031), .I0(n9031[6]), .I1(GND_net), .CO(n32032));
    SB_CARRY add_4613_11 (.CI(n32266), .I0(n9316[8]), .I1(GND_net), .CO(n32267));
    SB_LUT4 add_4613_10_lut (.I0(GND_net), .I1(n9316[7]), .I2(GND_net), 
            .I3(n32265), .O(n9303[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4613_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4592_8_lut (.I0(GND_net), .I1(n9031[5]), .I2(n551_adj_3790), 
            .I3(n32030), .O(n9019[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4592_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4613_10 (.CI(n32265), .I0(n9316[7]), .I1(GND_net), .CO(n32266));
    SB_LUT4 add_4613_9_lut (.I0(GND_net), .I1(n9316[6]), .I2(GND_net), 
            .I3(n32264), .O(n9303[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4613_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4592_8 (.CI(n32030), .I0(n9031[5]), .I1(n551_adj_3790), 
            .CO(n32031));
    SB_CARRY add_4613_9 (.CI(n32264), .I0(n9316[6]), .I1(GND_net), .CO(n32265));
    SB_LUT4 add_4613_8_lut (.I0(GND_net), .I1(n9316[5]), .I2(n548), .I3(n32263), 
            .O(n9303[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4613_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4592_7_lut (.I0(GND_net), .I1(n9031[4]), .I2(n478_adj_3791), 
            .I3(n32029), .O(n9019[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4592_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4613_8 (.CI(n32263), .I0(n9316[5]), .I1(n548), .CO(n32264));
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4613_7_lut (.I0(GND_net), .I1(n9316[4]), .I2(n475), .I3(n32262), 
            .O(n9303[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4613_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4592_7 (.CI(n32029), .I0(n9031[4]), .I1(n478_adj_3791), 
            .CO(n32030));
    SB_LUT4 i2_4_lut (.I0(n6_adj_3759), .I1(\Ki[4] ), .I2(n9373[2]), .I3(\PID_CONTROLLER.integral [18]), 
            .O(n9366[3]));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 add_4592_6_lut (.I0(GND_net), .I1(n9031[3]), .I2(n405_adj_3792), 
            .I3(n32028), .O(n9019[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4592_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4613_7 (.CI(n32262), .I0(n9316[4]), .I1(n475), .CO(n32263));
    SB_CARRY add_4592_6 (.CI(n32028), .I0(n9031[3]), .I1(n405_adj_3792), 
            .CO(n32029));
    SB_LUT4 add_4592_5_lut (.I0(GND_net), .I1(n9031[2]), .I2(n332_adj_3793), 
            .I3(n32027), .O(n9019[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4592_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4613_6_lut (.I0(GND_net), .I1(n9316[3]), .I2(n402), .I3(n32261), 
            .O(n9303[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4613_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4592_5 (.CI(n32027), .I0(n9031[2]), .I1(n332_adj_3793), 
            .CO(n32028));
    SB_CARRY add_4613_6 (.CI(n32261), .I0(n9316[3]), .I1(n402), .CO(n32262));
    SB_LUT4 add_4592_4_lut (.I0(GND_net), .I1(n9031[1]), .I2(n259_adj_3794), 
            .I3(n32026), .O(n9019[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4592_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4592_4 (.CI(n32026), .I0(n9031[1]), .I1(n259_adj_3794), 
            .CO(n32027));
    SB_LUT4 add_4613_5_lut (.I0(GND_net), .I1(n9316[2]), .I2(n329), .I3(n32260), 
            .O(n9303[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4613_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4592_3_lut (.I0(GND_net), .I1(n9031[0]), .I2(n186_adj_3795), 
            .I3(n32025), .O(n9019[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4592_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4613_5 (.CI(n32260), .I0(n9316[2]), .I1(n329), .CO(n32261));
    SB_CARRY add_4592_3 (.CI(n32025), .I0(n9031[0]), .I1(n186_adj_3795), 
            .CO(n32026));
    SB_LUT4 add_4613_4_lut (.I0(GND_net), .I1(n9316[1]), .I2(n256_adj_3796), 
            .I3(n32259), .O(n9303[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4613_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4592_2_lut (.I0(GND_net), .I1(n44_adj_3797), .I2(n113_adj_3798), 
            .I3(GND_net), .O(n9019[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4592_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4592_2 (.CI(GND_net), .I0(n44_adj_3797), .I1(n113_adj_3798), 
            .CO(n32025));
    SB_CARRY add_4613_4 (.CI(n32259), .I0(n9316[1]), .I1(n256_adj_3796), 
            .CO(n32260));
    SB_LUT4 add_4591_12_lut (.I0(GND_net), .I1(n9019[9]), .I2(GND_net), 
            .I3(n32024), .O(n9006[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4591_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4591_11_lut (.I0(GND_net), .I1(n9019[8]), .I2(GND_net), 
            .I3(n32023), .O(n9006[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4591_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4591_11 (.CI(n32023), .I0(n9019[8]), .I1(GND_net), .CO(n32024));
    SB_LUT4 add_4591_10_lut (.I0(GND_net), .I1(n9019[7]), .I2(GND_net), 
            .I3(n32022), .O(n9006[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4591_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4591_10 (.CI(n32022), .I0(n9019[7]), .I1(GND_net), .CO(n32023));
    SB_LUT4 add_4591_9_lut (.I0(GND_net), .I1(n9019[6]), .I2(GND_net), 
            .I3(n32021), .O(n9006[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4591_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4591_9 (.CI(n32021), .I0(n9019[6]), .I1(GND_net), .CO(n32022));
    SB_LUT4 add_4613_3_lut (.I0(GND_net), .I1(n9316[0]), .I2(n183_adj_3799), 
            .I3(n32258), .O(n9303[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4613_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4591_8_lut (.I0(GND_net), .I1(n9019[5]), .I2(n548_adj_3800), 
            .I3(n32020), .O(n9006[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4591_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4613_3 (.CI(n32258), .I0(n9316[0]), .I1(n183_adj_3799), 
            .CO(n32259));
    SB_LUT4 add_4613_2_lut (.I0(GND_net), .I1(n41_adj_3801), .I2(n110_adj_3802), 
            .I3(GND_net), .O(n9303[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4613_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4591_8 (.CI(n32020), .I0(n9019[5]), .I1(n548_adj_3800), 
            .CO(n32021));
    SB_LUT4 add_4591_7_lut (.I0(GND_net), .I1(n9019[4]), .I2(n475_adj_3803), 
            .I3(n32019), .O(n9006[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4591_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4613_2 (.CI(GND_net), .I0(n41_adj_3801), .I1(n110_adj_3802), 
            .CO(n32258));
    SB_CARRY add_4591_7 (.CI(n32019), .I0(n9019[4]), .I1(n475_adj_3803), 
            .CO(n32020));
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_25_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(n31207), .O(n34[23])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_25_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_24_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(n31206), .O(n34[22])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_24_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_4612_13_lut (.I0(GND_net), .I1(n9303[10]), .I2(GND_net), 
            .I3(n32257), .O(n9289[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4591_6_lut (.I0(GND_net), .I1(n9019[3]), .I2(n402_adj_3804), 
            .I3(n32018), .O(n9006[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4591_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4612_12_lut (.I0(GND_net), .I1(n9303[9]), .I2(GND_net), 
            .I3(n32256), .O(n9289[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4591_6 (.CI(n32018), .I0(n9019[3]), .I1(n402_adj_3804), 
            .CO(n32019));
    SB_CARRY add_4612_12 (.CI(n32256), .I0(n9303[9]), .I1(GND_net), .CO(n32257));
    SB_LUT4 add_4612_11_lut (.I0(GND_net), .I1(n9303[8]), .I2(GND_net), 
            .I3(n32255), .O(n9289[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4591_5_lut (.I0(GND_net), .I1(n9019[2]), .I2(n329_adj_3805), 
            .I3(n32017), .O(n9006[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4591_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_24  (.CI(n31206), .I0(\PID_CONTROLLER.err [22]), 
            .I1(\PID_CONTROLLER.integral [22]), .CO(n31207));
    SB_CARRY add_4612_11 (.CI(n32255), .I0(n9303[8]), .I1(GND_net), .CO(n32256));
    SB_CARRY add_4591_5 (.CI(n32017), .I0(n9019[2]), .I1(n329_adj_3805), 
            .CO(n32018));
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_23_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(n31205), .O(n34[21])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_23_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_4612_10_lut (.I0(GND_net), .I1(n9303[7]), .I2(GND_net), 
            .I3(n32254), .O(n9289[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4591_4_lut (.I0(GND_net), .I1(n9019[1]), .I2(n256_adj_3806), 
            .I3(n32016), .O(n9006[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4591_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_23  (.CI(n31205), .I0(\PID_CONTROLLER.err [21]), 
            .I1(\PID_CONTROLLER.integral [21]), .CO(n31206));
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_22_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(n31204), .O(n34[20])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_22_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_4591_4 (.CI(n32016), .I0(n9019[1]), .I1(n256_adj_3806), 
            .CO(n32017));
    SB_LUT4 state_23__I_0_add_2_22_lut (.I0(GND_net), .I1(motor_state[20]), 
            .I2(n1_adj_3898[20]), .I3(n30520), .O(\PID_CONTROLLER.err_23__N_3379 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_22 (.CI(n30520), .I0(motor_state[20]), 
            .I1(n1_adj_3898[20]), .CO(n30521));
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_22  (.CI(n31204), .I0(\PID_CONTROLLER.err [20]), 
            .I1(\PID_CONTROLLER.integral [20]), .CO(n31205));
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_21_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.integral [19]), .I3(n31203), .O(n34[19])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_21_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_4612_10 (.CI(n32254), .I0(n9303[7]), .I1(GND_net), .CO(n32255));
    SB_LUT4 add_4612_9_lut (.I0(GND_net), .I1(n9303[6]), .I2(GND_net), 
            .I3(n32253), .O(n9289[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4591_3_lut (.I0(GND_net), .I1(n9019[0]), .I2(n183_adj_3808), 
            .I3(n32015), .O(n9006[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4591_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4612_9 (.CI(n32253), .I0(n9303[6]), .I1(GND_net), .CO(n32254));
    SB_CARRY add_4591_3 (.CI(n32015), .I0(n9019[0]), .I1(n183_adj_3808), 
            .CO(n32016));
    SB_LUT4 add_4591_2_lut (.I0(GND_net), .I1(n41_adj_3809), .I2(n110_adj_3810), 
            .I3(GND_net), .O(n9006[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4591_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_21  (.CI(n31203), .I0(\PID_CONTROLLER.err [19]), 
            .I1(\PID_CONTROLLER.integral [19]), .CO(n31204));
    SB_LUT4 add_4612_8_lut (.I0(GND_net), .I1(n9303[5]), .I2(n545), .I3(n32252), 
            .O(n9289[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4591_2 (.CI(GND_net), .I0(n41_adj_3809), .I1(n110_adj_3810), 
            .CO(n32015));
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_20_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [18]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(n31202), .O(n34[18])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_20_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_20  (.CI(n31202), .I0(\PID_CONTROLLER.err [18]), 
            .I1(\PID_CONTROLLER.integral [18]), .CO(n31203));
    SB_CARRY add_4612_8 (.CI(n32252), .I0(n9303[5]), .I1(n545), .CO(n32253));
    SB_LUT4 add_4590_13_lut (.I0(GND_net), .I1(n9006[10]), .I2(GND_net), 
            .I3(n32014), .O(n8992[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4590_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_19_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(n31201), .O(n34[17])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_19_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_21_lut (.I0(GND_net), .I1(motor_state[19]), 
            .I2(n1_adj_3898[19]), .I3(n30519), .O(\PID_CONTROLLER.err_23__N_3379 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4612_7_lut (.I0(GND_net), .I1(n9303[4]), .I2(n472), .I3(n32251), 
            .O(n9289[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4590_12_lut (.I0(GND_net), .I1(n9006[9]), .I2(GND_net), 
            .I3(n32013), .O(n8992[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4590_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4612_7 (.CI(n32251), .I0(n9303[4]), .I1(n472), .CO(n32252));
    SB_CARRY add_4590_12 (.CI(n32013), .I0(n9006[9]), .I1(GND_net), .CO(n32014));
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_19  (.CI(n31201), .I0(\PID_CONTROLLER.err [17]), 
            .I1(\PID_CONTROLLER.integral [17]), .CO(n31202));
    SB_LUT4 add_4612_6_lut (.I0(GND_net), .I1(n9303[3]), .I2(n399), .I3(n32250), 
            .O(n9289[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4590_11_lut (.I0(GND_net), .I1(n9006[8]), .I2(GND_net), 
            .I3(n32012), .O(n8992[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4590_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_18_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(n31200), .O(n34[16])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_18_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_4590_11 (.CI(n32012), .I0(n9006[8]), .I1(GND_net), .CO(n32013));
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_18  (.CI(n31200), .I0(\PID_CONTROLLER.err [16]), 
            .I1(\PID_CONTROLLER.integral [16]), .CO(n31201));
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_17_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [15]), 
            .I2(\PID_CONTROLLER.integral [15]), .I3(n31199), .O(n34[15])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_17_lut .LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_21 (.CI(n30519), .I0(motor_state[19]), 
            .I1(n1_adj_3898[19]), .CO(n30520));
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_17  (.CI(n31199), .I0(\PID_CONTROLLER.err [15]), 
            .I1(\PID_CONTROLLER.integral [15]), .CO(n31200));
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_16_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [14]), 
            .I2(\PID_CONTROLLER.integral [14]), .I3(n31198), .O(n34[14])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_16_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_16  (.CI(n31198), .I0(\PID_CONTROLLER.err [14]), 
            .I1(\PID_CONTROLLER.integral [14]), .CO(n31199));
    SB_CARRY add_4612_6 (.CI(n32250), .I0(n9303[3]), .I1(n399), .CO(n32251));
    SB_LUT4 add_4590_10_lut (.I0(GND_net), .I1(n9006[7]), .I2(GND_net), 
            .I3(n32011), .O(n8992[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4590_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4612_5_lut (.I0(GND_net), .I1(n9303[2]), .I2(n326), .I3(n32249), 
            .O(n9289[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4612_5 (.CI(n32249), .I0(n9303[2]), .I1(n326), .CO(n32250));
    SB_CARRY add_4590_10 (.CI(n32011), .I0(n9006[7]), .I1(GND_net), .CO(n32012));
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_15_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [13]), 
            .I2(\PID_CONTROLLER.integral [13]), .I3(n31197), .O(n34[13])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_15_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_15  (.CI(n31197), .I0(\PID_CONTROLLER.err [13]), 
            .I1(\PID_CONTROLLER.integral [13]), .CO(n31198));
    SB_LUT4 add_4612_4_lut (.I0(GND_net), .I1(n9303[1]), .I2(n253), .I3(n32248), 
            .O(n9289[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4590_9_lut (.I0(GND_net), .I1(n9006[6]), .I2(GND_net), 
            .I3(n32010), .O(n8992[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4590_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_14_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [12]), 
            .I2(\PID_CONTROLLER.integral [12]), .I3(n31196), .O(n34[12])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_14_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_4612_4 (.CI(n32248), .I0(n9303[1]), .I1(n253), .CO(n32249));
    SB_CARRY add_4590_9 (.CI(n32010), .I0(n9006[6]), .I1(GND_net), .CO(n32011));
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_14  (.CI(n31196), .I0(\PID_CONTROLLER.err [12]), 
            .I1(\PID_CONTROLLER.integral [12]), .CO(n31197));
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_13_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [11]), 
            .I2(\PID_CONTROLLER.integral [11]), .I3(n31195), .O(n34[11])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_13_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_20_lut (.I0(GND_net), .I1(motor_state[18]), 
            .I2(n1_adj_3898[18]), .I3(n30518), .O(\PID_CONTROLLER.err_23__N_3379 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4612_3_lut (.I0(GND_net), .I1(n9303[0]), .I2(n180), .I3(n32247), 
            .O(n9289[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_628_25_lut (.I0(GND_net), .I1(n2942[23]), .I2(n2967[23]), 
            .I3(n30377), .O(duty_23__N_3478[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_628_24_lut (.I0(GND_net), .I1(n2942[22]), .I2(n2967[22]), 
            .I3(n30376), .O(duty_23__N_3478[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4612_3 (.CI(n32247), .I0(n9303[0]), .I1(n180), .CO(n32248));
    SB_LUT4 add_4590_8_lut (.I0(GND_net), .I1(n9006[5]), .I2(n545_adj_3813), 
            .I3(n32009), .O(n8992[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4590_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4612_2_lut (.I0(GND_net), .I1(n38), .I2(n107_adj_3814), 
            .I3(GND_net), .O(n9289[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4612_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4590_8 (.CI(n32009), .I0(n9006[5]), .I1(n545_adj_3813), 
            .CO(n32010));
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_13  (.CI(n31195), .I0(\PID_CONTROLLER.err [11]), 
            .I1(\PID_CONTROLLER.integral [11]), .CO(n31196));
    SB_CARRY add_4612_2 (.CI(GND_net), .I0(n38), .I1(n107_adj_3814), .CO(n32247));
    SB_LUT4 add_4611_14_lut (.I0(GND_net), .I1(n9289[11]), .I2(GND_net), 
            .I3(n32246), .O(n9274[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4590_7_lut (.I0(GND_net), .I1(n9006[4]), .I2(n472_adj_3815), 
            .I3(n32008), .O(n8992[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4590_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4590_7 (.CI(n32008), .I0(n9006[4]), .I1(n472_adj_3815), 
            .CO(n32009));
    SB_LUT4 add_4590_6_lut (.I0(GND_net), .I1(n9006[3]), .I2(n399_adj_3816), 
            .I3(n32007), .O(n8992[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4590_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_12_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [10]), 
            .I2(\PID_CONTROLLER.integral [10]), .I3(n31194), .O(n34[10])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_12_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_12  (.CI(n31194), .I0(\PID_CONTROLLER.err [10]), 
            .I1(\PID_CONTROLLER.integral [10]), .CO(n31195));
    SB_CARRY add_4590_6 (.CI(n32007), .I0(n9006[3]), .I1(n399_adj_3816), 
            .CO(n32008));
    SB_LUT4 add_4590_5_lut (.I0(GND_net), .I1(n9006[2]), .I2(n326_adj_3817), 
            .I3(n32006), .O(n8992[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4590_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_11_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [9]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(n31193), .O(n34[9])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_11_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_4611_13_lut (.I0(GND_net), .I1(n9289[10]), .I2(GND_net), 
            .I3(n32245), .O(n9274[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4590_5 (.CI(n32006), .I0(n9006[2]), .I1(n326_adj_3817), 
            .CO(n32007));
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_11  (.CI(n31193), .I0(\PID_CONTROLLER.err [9]), 
            .I1(\PID_CONTROLLER.integral [9]), .CO(n31194));
    SB_LUT4 add_4590_4_lut (.I0(GND_net), .I1(n9006[1]), .I2(n253_adj_3818), 
            .I3(n32005), .O(n8992[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4590_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_10_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(n31192), .O(n34[8])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_10_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_628_24 (.CI(n30376), .I0(n2942[22]), .I1(n2967[22]), 
            .CO(n30377));
    SB_CARRY add_4611_13 (.CI(n32245), .I0(n9289[10]), .I1(GND_net), .CO(n32246));
    SB_CARRY add_4590_4 (.CI(n32005), .I0(n9006[1]), .I1(n253_adj_3818), 
            .CO(n32006));
    SB_LUT4 add_4611_12_lut (.I0(GND_net), .I1(n9289[9]), .I2(GND_net), 
            .I3(n32244), .O(n9274[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_10  (.CI(n31192), .I0(\PID_CONTROLLER.err [8]), 
            .I1(\PID_CONTROLLER.integral [8]), .CO(n31193));
    SB_LUT4 add_4590_3_lut (.I0(GND_net), .I1(n9006[0]), .I2(n180_adj_3819), 
            .I3(n32004), .O(n8992[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4590_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_9_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [7]), 
            .I2(\PID_CONTROLLER.integral [7]), .I3(n31191), .O(n34[7])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_9_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_4611_12 (.CI(n32244), .I0(n9289[9]), .I1(GND_net), .CO(n32245));
    SB_CARRY add_4590_3 (.CI(n32004), .I0(n9006[0]), .I1(n180_adj_3819), 
            .CO(n32005));
    SB_LUT4 add_4590_2_lut (.I0(GND_net), .I1(n38_adj_3820), .I2(n107_adj_3821), 
            .I3(GND_net), .O(n8992[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4590_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_9  (.CI(n31191), .I0(\PID_CONTROLLER.err [7]), 
            .I1(\PID_CONTROLLER.integral [7]), .CO(n31192));
    SB_CARRY state_23__I_0_add_2_20 (.CI(n30518), .I0(motor_state[18]), 
            .I1(n1_adj_3898[18]), .CO(n30519));
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_8_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(n31190), .O(n34[6])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_8_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_4611_11_lut (.I0(GND_net), .I1(n9289[8]), .I2(GND_net), 
            .I3(n32243), .O(n9274[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4590_2 (.CI(GND_net), .I0(n38_adj_3820), .I1(n107_adj_3821), 
            .CO(n32004));
    SB_LUT4 add_4589_14_lut (.I0(GND_net), .I1(n8992[11]), .I2(GND_net), 
            .I3(n32003), .O(n8977[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4589_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_8  (.CI(n31190), .I0(\PID_CONTROLLER.err [6]), 
            .I1(\PID_CONTROLLER.integral [6]), .CO(n31191));
    SB_LUT4 add_628_23_lut (.I0(GND_net), .I1(n2942[21]), .I2(n2967[21]), 
            .I3(n30375), .O(duty_23__N_3478[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4611_11 (.CI(n32243), .I0(n9289[8]), .I1(GND_net), .CO(n32244));
    SB_LUT4 state_23__I_0_add_2_19_lut (.I0(GND_net), .I1(motor_state[17]), 
            .I2(n1_adj_3898[17]), .I3(n30517), .O(\PID_CONTROLLER.err_23__N_3379 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_7_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [5]), 
            .I2(\PID_CONTROLLER.integral [5]), .I3(n31189), .O(n34[5])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_7_lut .LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_19 (.CI(n30517), .I0(motor_state[17]), 
            .I1(n1_adj_3898[17]), .CO(n30518));
    SB_LUT4 add_4611_10_lut (.I0(GND_net), .I1(n9289[7]), .I2(GND_net), 
            .I3(n32242), .O(n9274[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4589_13_lut (.I0(GND_net), .I1(n8992[10]), .I2(GND_net), 
            .I3(n32002), .O(n8977[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4589_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_7  (.CI(n31189), .I0(\PID_CONTROLLER.err [5]), 
            .I1(\PID_CONTROLLER.integral [5]), .CO(n31190));
    SB_CARRY add_4611_10 (.CI(n32242), .I0(n9289[7]), .I1(GND_net), .CO(n32243));
    SB_CARRY add_4589_13 (.CI(n32002), .I0(n8992[10]), .I1(GND_net), .CO(n32003));
    SB_LUT4 add_4589_12_lut (.I0(GND_net), .I1(n8992[9]), .I2(GND_net), 
            .I3(n32001), .O(n8977[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4589_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_6_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [4]), 
            .I2(\PID_CONTROLLER.integral [4]), .I3(n31188), .O(n34[4])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_6_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_4611_9_lut (.I0(GND_net), .I1(n9289[6]), .I2(GND_net), 
            .I3(n32241), .O(n9274[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_18_lut (.I0(GND_net), .I1(motor_state[16]), 
            .I2(n1_adj_3898[16]), .I3(n30516), .O(\PID_CONTROLLER.err_23__N_3379 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_18 (.CI(n30516), .I0(motor_state[16]), 
            .I1(n1_adj_3898[16]), .CO(n30517));
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_6  (.CI(n31188), .I0(\PID_CONTROLLER.err [4]), 
            .I1(\PID_CONTROLLER.integral [4]), .CO(n31189));
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_5_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(n31187), .O(n34[3])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_5_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_17_lut (.I0(GND_net), .I1(motor_state[15]), 
            .I2(n1_adj_3898[15]), .I3(n30515), .O(\PID_CONTROLLER.err_23__N_3379 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4611_9 (.CI(n32241), .I0(n9289[6]), .I1(GND_net), .CO(n32242));
    SB_CARRY add_4589_12 (.CI(n32001), .I0(n8992[9]), .I1(GND_net), .CO(n32002));
    SB_LUT4 add_4611_8_lut (.I0(GND_net), .I1(n9289[5]), .I2(n542), .I3(n32240), 
            .O(n9274[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4589_11_lut (.I0(GND_net), .I1(n8992[8]), .I2(GND_net), 
            .I3(n32000), .O(n8977[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4589_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_5  (.CI(n31187), .I0(\PID_CONTROLLER.err [3]), 
            .I1(\PID_CONTROLLER.integral [3]), .CO(n31188));
    SB_CARRY state_23__I_0_add_2_17 (.CI(n30515), .I0(motor_state[15]), 
            .I1(n1_adj_3898[15]), .CO(n30516));
    SB_CARRY add_628_23 (.CI(n30375), .I0(n2942[21]), .I1(n2967[21]), 
            .CO(n30376));
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_4_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [2]), 
            .I2(\PID_CONTROLLER.integral [2]), .I3(n31186), .O(n34[2])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_4_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_4611_8 (.CI(n32240), .I0(n9289[5]), .I1(n542), .CO(n32241));
    SB_CARRY add_4589_11 (.CI(n32000), .I0(n8992[8]), .I1(GND_net), .CO(n32001));
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_4  (.CI(n31186), .I0(\PID_CONTROLLER.err [2]), 
            .I1(\PID_CONTROLLER.integral [2]), .CO(n31187));
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_3_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [1]), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(n31185), .O(n34[1])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_3_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_3  (.CI(n31185), .I0(\PID_CONTROLLER.err [1]), 
            .I1(\PID_CONTROLLER.integral [1]), .CO(n31186));
    SB_LUT4 mult_11_i138_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_628_22_lut (.I0(GND_net), .I1(n2942[20]), .I2(n2967[20]), 
            .I3(n30374), .O(duty_23__N_3478[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_16_lut (.I0(GND_net), .I1(motor_state[14]), 
            .I2(n1_adj_3898[14]), .I3(n30514), .O(\PID_CONTROLLER.err_23__N_3379 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_22 (.CI(n30374), .I0(n2942[20]), .I1(n2967[20]), 
            .CO(n30375));
    SB_LUT4 i25262_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [22]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n9384[0]));   // verilog/motorControl.v(42[26:37])
    defparam i25262_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_628_21_lut (.I0(GND_net), .I1(n2942[19]), .I2(n2967[19]), 
            .I3(n30373), .O(duty_23__N_3478[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_21 (.CI(n30373), .I0(n2942[19]), .I1(n2967[19]), 
            .CO(n30374));
    SB_LUT4 add_628_20_lut (.I0(GND_net), .I1(n2942[18]), .I2(n2967[18]), 
            .I3(n30372), .O(duty_23__N_3478[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4589_10_lut (.I0(GND_net), .I1(n8992[7]), .I2(GND_net), 
            .I3(n31999), .O(n8977[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4589_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4611_7_lut (.I0(GND_net), .I1(n9289[4]), .I2(n469), .I3(n32239), 
            .O(n9274[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4611_7 (.CI(n32239), .I0(n9289[4]), .I1(n469), .CO(n32240));
    SB_CARRY add_4589_10 (.CI(n31999), .I0(n8992[7]), .I1(GND_net), .CO(n32000));
    SB_LUT4 \PID_CONTROLLER.integral_1149_add_4_2_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [0]), 
            .I2(\PID_CONTROLLER.integral [0]), .I3(GND_net), .O(n34[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1149_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_4589_9_lut (.I0(GND_net), .I1(n8992[6]), .I2(GND_net), 
            .I3(n31998), .O(n8977[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4589_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4611_6_lut (.I0(GND_net), .I1(n9289[3]), .I2(n396), .I3(n32238), 
            .O(n9274[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4589_9 (.CI(n31998), .I0(n8992[6]), .I1(GND_net), .CO(n31999));
    SB_CARRY \PID_CONTROLLER.integral_1149_add_4_2  (.CI(GND_net), .I0(\PID_CONTROLLER.err [0]), 
            .I1(\PID_CONTROLLER.integral [0]), .CO(n31185));
    SB_CARRY state_23__I_0_add_2_16 (.CI(n30514), .I0(motor_state[14]), 
            .I1(n1_adj_3898[14]), .CO(n30515));
    SB_LUT4 mult_11_i89_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i89_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4611_6 (.CI(n32238), .I0(n9289[3]), .I1(n396), .CO(n32239));
    SB_LUT4 add_4589_8_lut (.I0(GND_net), .I1(n8992[5]), .I2(n542_adj_3826), 
            .I3(n31997), .O(n8977[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4589_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4611_5_lut (.I0(GND_net), .I1(n9289[2]), .I2(n323), .I3(n32237), 
            .O(n9274[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4589_8 (.CI(n31997), .I0(n8992[5]), .I1(n542_adj_3826), 
            .CO(n31998));
    SB_LUT4 mult_11_i42_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i42_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4611_5 (.CI(n32237), .I0(n9289[2]), .I1(n323), .CO(n32238));
    SB_LUT4 add_4589_7_lut (.I0(GND_net), .I1(n8992[4]), .I2(n469_adj_3827), 
            .I3(n31996), .O(n8977[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4589_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4611_4_lut (.I0(GND_net), .I1(n9289[1]), .I2(n250), .I3(n32236), 
            .O(n9274[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4589_7 (.CI(n31996), .I0(n8992[4]), .I1(n469_adj_3827), 
            .CO(n31997));
    SB_CARRY add_4611_4 (.CI(n32236), .I0(n9289[1]), .I1(n250), .CO(n32237));
    SB_LUT4 add_4589_6_lut (.I0(GND_net), .I1(n8992[3]), .I2(n396_adj_3828), 
            .I3(n31995), .O(n8977[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4589_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4611_3_lut (.I0(GND_net), .I1(n9289[0]), .I2(n177), .I3(n32235), 
            .O(n9274[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4589_6 (.CI(n31995), .I0(n8992[3]), .I1(n396_adj_3828), 
            .CO(n31996));
    SB_LUT4 add_4589_5_lut (.I0(GND_net), .I1(n8992[2]), .I2(n323_adj_3829), 
            .I3(n31994), .O(n8977[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4589_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_15_lut (.I0(GND_net), .I1(motor_state[13]), 
            .I2(n1_adj_3898[13]), .I3(n30513), .O(\PID_CONTROLLER.err_23__N_3379 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4611_3 (.CI(n32235), .I0(n9289[0]), .I1(n177), .CO(n32236));
    SB_CARRY add_4589_5 (.CI(n31994), .I0(n8992[2]), .I1(n323_adj_3829), 
            .CO(n31995));
    SB_LUT4 add_4611_2_lut (.I0(GND_net), .I1(n35_adj_3831), .I2(n104_adj_3832), 
            .I3(GND_net), .O(n9274[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4611_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4589_4_lut (.I0(GND_net), .I1(n8992[1]), .I2(n250_adj_3833), 
            .I3(n31993), .O(n8977[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4589_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4611_2 (.CI(GND_net), .I0(n35_adj_3831), .I1(n104_adj_3832), 
            .CO(n32235));
    SB_CARRY add_4589_4 (.CI(n31993), .I0(n8992[1]), .I1(n250_adj_3833), 
            .CO(n31994));
    SB_LUT4 add_4610_15_lut (.I0(GND_net), .I1(n9274[12]), .I2(GND_net), 
            .I3(n32234), .O(n9258[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4589_3_lut (.I0(GND_net), .I1(n8992[0]), .I2(n177_adj_3834), 
            .I3(n31992), .O(n8977[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4589_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4610_14_lut (.I0(GND_net), .I1(n9274[11]), .I2(GND_net), 
            .I3(n32233), .O(n9258[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4589_3 (.CI(n31992), .I0(n8992[0]), .I1(n177_adj_3834), 
            .CO(n31993));
    SB_CARRY add_4610_14 (.CI(n32233), .I0(n9274[11]), .I1(GND_net), .CO(n32234));
    SB_LUT4 add_4589_2_lut (.I0(GND_net), .I1(n35_adj_3835), .I2(n104_adj_3836), 
            .I3(GND_net), .O(n8977[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4589_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4589_2 (.CI(GND_net), .I0(n35_adj_3835), .I1(n104_adj_3836), 
            .CO(n31992));
    SB_CARRY state_23__I_0_add_2_15 (.CI(n30513), .I0(motor_state[13]), 
            .I1(n1_adj_3898[13]), .CO(n30514));
    SB_LUT4 add_4610_13_lut (.I0(GND_net), .I1(n9274[10]), .I2(GND_net), 
            .I3(n32232), .O(n9258[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4610_13 (.CI(n32232), .I0(n9274[10]), .I1(GND_net), .CO(n32233));
    SB_LUT4 add_4588_15_lut (.I0(GND_net), .I1(n8977[12]), .I2(GND_net), 
            .I3(n31991), .O(n8961[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4588_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4588_14_lut (.I0(GND_net), .I1(n8977[11]), .I2(GND_net), 
            .I3(n31990), .O(n8961[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4588_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_20 (.CI(n30372), .I0(n2942[18]), .I1(n2967[18]), 
            .CO(n30373));
    SB_LUT4 add_4610_12_lut (.I0(GND_net), .I1(n9274[9]), .I2(GND_net), 
            .I3(n32231), .O(n9258[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4588_14 (.CI(n31990), .I0(n8977[11]), .I1(GND_net), .CO(n31991));
    SB_CARRY add_4610_12 (.CI(n32231), .I0(n9274[9]), .I1(GND_net), .CO(n32232));
    SB_LUT4 add_4588_13_lut (.I0(GND_net), .I1(n8977[10]), .I2(GND_net), 
            .I3(n31989), .O(n8961[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4588_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4610_11_lut (.I0(GND_net), .I1(n9274[8]), .I2(GND_net), 
            .I3(n32230), .O(n9258[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4588_13 (.CI(n31989), .I0(n8977[10]), .I1(GND_net), .CO(n31990));
    SB_LUT4 add_4588_12_lut (.I0(GND_net), .I1(n8977[9]), .I2(GND_net), 
            .I3(n31988), .O(n8961[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4588_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_849 (.I0(n4_adj_3764), .I1(\Ki[3] ), .I2(n9379[1]), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n9373[2]));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut_adj_849.LUT_INIT = 16'h965a;
    SB_CARRY add_4610_11 (.CI(n32230), .I0(n9274[8]), .I1(GND_net), .CO(n32231));
    SB_CARRY add_4588_12 (.CI(n31988), .I0(n8977[9]), .I1(GND_net), .CO(n31989));
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4610_10_lut (.I0(GND_net), .I1(n9274[7]), .I2(GND_net), 
            .I3(n32229), .O(n9258[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4588_11_lut (.I0(GND_net), .I1(n8977[8]), .I2(GND_net), 
            .I3(n31987), .O(n8961[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4588_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_850 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral [23]), 
            .I3(\PID_CONTROLLER.integral [20]), .O(n12_adj_3837));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut_adj_850.LUT_INIT = 16'h9c50;
    SB_CARRY add_4610_10 (.CI(n32229), .I0(n9274[7]), .I1(GND_net), .CO(n32230));
    SB_CARRY add_4588_11 (.CI(n31987), .I0(n8977[8]), .I1(GND_net), .CO(n31988));
    SB_LUT4 add_4588_10_lut (.I0(GND_net), .I1(n8977[7]), .I2(GND_net), 
            .I3(n31986), .O(n8961[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4588_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4610_9_lut (.I0(GND_net), .I1(n9274[6]), .I2(GND_net), 
            .I3(n32228), .O(n9258[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4588_10 (.CI(n31986), .I0(n8977[7]), .I1(GND_net), .CO(n31987));
    SB_CARRY add_4610_9 (.CI(n32228), .I0(n9274[6]), .I1(GND_net), .CO(n32229));
    SB_LUT4 add_4588_9_lut (.I0(GND_net), .I1(n8977[6]), .I2(GND_net), 
            .I3(n31985), .O(n8961[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4588_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4588_9 (.CI(n31985), .I0(n8977[6]), .I1(GND_net), .CO(n31986));
    SB_LUT4 i25198_4_lut (.I0(n9373[2]), .I1(\Ki[4] ), .I2(n6_adj_3759), 
            .I3(\PID_CONTROLLER.integral [18]), .O(n8_adj_3838));   // verilog/motorControl.v(42[26:37])
    defparam i25198_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 add_628_19_lut (.I0(GND_net), .I1(n2942[17]), .I2(n2967[17]), 
            .I3(n30371), .O(duty_23__N_3478[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4610_8_lut (.I0(GND_net), .I1(n9274[5]), .I2(n539), .I3(n32227), 
            .O(n9258[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4588_8_lut (.I0(GND_net), .I1(n8977[5]), .I2(n539_adj_3839), 
            .I3(n31984), .O(n8961[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4588_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_851 (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n11_adj_3840));   // verilog/motorControl.v(42[26:37])
    defparam i1_4_lut_adj_851.LUT_INIT = 16'h6ca0;
    SB_CARRY add_4610_8 (.CI(n32227), .I0(n9274[5]), .I1(n539), .CO(n32228));
    SB_CARRY add_4588_8 (.CI(n31984), .I0(n8977[5]), .I1(n539_adj_3839), 
            .CO(n31985));
    SB_LUT4 i25229_4_lut (.I0(n9379[1]), .I1(\Ki[3] ), .I2(n4_adj_3764), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n6_adj_3841));   // verilog/motorControl.v(42[26:37])
    defparam i25229_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 add_4610_7_lut (.I0(GND_net), .I1(n9274[4]), .I2(n466), .I3(n32226), 
            .O(n9258[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4588_7_lut (.I0(GND_net), .I1(n8977[4]), .I2(n466_adj_3842), 
            .I3(n31983), .O(n8961[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4588_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4588_7 (.CI(n31983), .I0(n8977[4]), .I1(n466_adj_3842), 
            .CO(n31984));
    SB_CARRY add_4610_7 (.CI(n32226), .I0(n9274[4]), .I1(n466), .CO(n32227));
    SB_LUT4 add_4588_6_lut (.I0(GND_net), .I1(n8977[3]), .I2(n393), .I3(n31982), 
            .O(n8961[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4588_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4588_6 (.CI(n31982), .I0(n8977[3]), .I1(n393), .CO(n31983));
    SB_LUT4 state_23__I_0_add_2_14_lut (.I0(GND_net), .I1(motor_state[12]), 
            .I2(n1_adj_3898[12]), .I3(n30512), .O(\PID_CONTROLLER.err_23__N_3379 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_14 (.CI(n30512), .I0(motor_state[12]), 
            .I1(n1_adj_3898[12]), .CO(n30513));
    SB_LUT4 i25264_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [22]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n30231));   // verilog/motorControl.v(42[26:37])
    defparam i25264_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 state_23__I_0_add_2_13_lut (.I0(GND_net), .I1(motor_state[11]), 
            .I2(n1_adj_3898[11]), .I3(n30511), .O(\PID_CONTROLLER.err_23__N_3379 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8_4_lut_adj_852 (.I0(n6_adj_3841), .I1(n11_adj_3840), .I2(n8_adj_3838), 
            .I3(n12_adj_3837), .O(n18_adj_3845));   // verilog/motorControl.v(42[26:37])
    defparam i8_4_lut_adj_852.LUT_INIT = 16'h6996;
    SB_CARRY state_23__I_0_add_2_13 (.CI(n30511), .I0(motor_state[11]), 
            .I1(n1_adj_3898[11]), .CO(n30512));
    SB_LUT4 i3_4_lut_adj_853 (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(\PID_CONTROLLER.integral [22]), .O(n13_adj_3846));   // verilog/motorControl.v(42[26:37])
    defparam i3_4_lut_adj_853.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_4610_6_lut (.I0(GND_net), .I1(n9274[3]), .I2(n393_adj_3847), 
            .I3(n32225), .O(n9258[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_12_lut (.I0(GND_net), .I1(motor_state[10]), 
            .I2(n1_adj_3898[10]), .I3(n30510), .O(\PID_CONTROLLER.err_23__N_3379 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4588_5_lut (.I0(GND_net), .I1(n8977[2]), .I2(n320), .I3(n31981), 
            .O(n8961[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4588_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4610_6 (.CI(n32225), .I0(n9274[3]), .I1(n393_adj_3847), 
            .CO(n32226));
    SB_CARRY add_4588_5 (.CI(n31981), .I0(n8977[2]), .I1(n320), .CO(n31982));
    SB_CARRY add_628_19 (.CI(n30371), .I0(n2942[17]), .I1(n2967[17]), 
            .CO(n30372));
    SB_LUT4 add_628_18_lut (.I0(GND_net), .I1(n2942[16]), .I2(n2967[16]), 
            .I3(n30370), .O(duty_23__N_3478[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4610_5_lut (.I0(GND_net), .I1(n9274[2]), .I2(n320_adj_3849), 
            .I3(n32224), .O(n9258[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_12 (.CI(n30510), .I0(motor_state[10]), 
            .I1(n1_adj_3898[10]), .CO(n30511));
    SB_CARRY add_4610_5 (.CI(n32224), .I0(n9274[2]), .I1(n320_adj_3849), 
            .CO(n32225));
    SB_LUT4 add_4588_4_lut (.I0(GND_net), .I1(n8977[1]), .I2(n247), .I3(n31980), 
            .O(n8961[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4588_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4588_4 (.CI(n31980), .I0(n8977[1]), .I1(n247), .CO(n31981));
    SB_CARRY add_628_18 (.CI(n30370), .I0(n2942[16]), .I1(n2967[16]), 
            .CO(n30371));
    SB_LUT4 state_23__I_0_add_2_11_lut (.I0(GND_net), .I1(motor_state[9]), 
            .I2(n1_adj_3898[9]), .I3(n30509), .O(\PID_CONTROLLER.err_23__N_3379 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_628_17_lut (.I0(GND_net), .I1(n2942[15]), .I2(n2967[15]), 
            .I3(n30369), .O(duty_23__N_3478[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9_4_lut_adj_854 (.I0(n13_adj_3846), .I1(n18_adj_3845), .I2(n30231), 
            .I3(n4_adj_3763), .O(n38956));   // verilog/motorControl.v(42[26:37])
    defparam i9_4_lut_adj_854.LUT_INIT = 16'h6996;
    SB_CARRY add_628_17 (.CI(n30369), .I0(n2942[15]), .I1(n2967[15]), 
            .CO(n30370));
    SB_LUT4 add_4588_3_lut (.I0(GND_net), .I1(n8977[0]), .I2(n174), .I3(n31979), 
            .O(n8961[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4588_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4610_4_lut (.I0(GND_net), .I1(n9274[1]), .I2(n247_adj_3851), 
            .I3(n32223), .O(n9258[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4588_3 (.CI(n31979), .I0(n8977[0]), .I1(n174), .CO(n31980));
    SB_LUT4 add_628_16_lut (.I0(GND_net), .I1(n2942[14]), .I2(n2967[14]), 
            .I3(n30368), .O(duty_23__N_3478[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_11 (.CI(n30509), .I0(motor_state[9]), .I1(n1_adj_3898[9]), 
            .CO(n30510));
    SB_LUT4 state_23__I_0_add_2_10_lut (.I0(GND_net), .I1(motor_state[8]), 
            .I2(n1_adj_3898[8]), .I3(n30508), .O(\PID_CONTROLLER.err_23__N_3379 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_10 (.CI(n30508), .I0(motor_state[8]), .I1(n1_adj_3898[8]), 
            .CO(n30509));
    SB_LUT4 add_4588_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n8961[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4588_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_16 (.CI(n30368), .I0(n2942[14]), .I1(n2967[14]), 
            .CO(n30369));
    SB_CARRY add_4610_4 (.CI(n32223), .I0(n9274[1]), .I1(n247_adj_3851), 
            .CO(n32224));
    SB_CARRY add_4588_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n31979));
    SB_LUT4 add_4610_3_lut (.I0(GND_net), .I1(n9274[0]), .I2(n174_adj_3853), 
            .I3(n32222), .O(n9258[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4610_3 (.CI(n32222), .I0(n9274[0]), .I1(n174_adj_3853), 
            .CO(n32223));
    SB_LUT4 add_4587_16_lut (.I0(GND_net), .I1(n8961[13]), .I2(GND_net), 
            .I3(n31978), .O(n8944[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4587_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4610_2_lut (.I0(GND_net), .I1(n32_adj_3854), .I2(n101_adj_3855), 
            .I3(GND_net), .O(n9258[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4610_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4587_15_lut (.I0(GND_net), .I1(n8961[12]), .I2(GND_net), 
            .I3(n31977), .O(n8944[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4587_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4610_2 (.CI(GND_net), .I0(n32_adj_3854), .I1(n101_adj_3855), 
            .CO(n32222));
    SB_LUT4 add_4609_16_lut (.I0(GND_net), .I1(n9258[13]), .I2(GND_net), 
            .I3(n32221), .O(n9241[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4609_15_lut (.I0(GND_net), .I1(n9258[12]), .I2(GND_net), 
            .I3(n32220), .O(n9241[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_15 (.CI(n32220), .I0(n9258[12]), .I1(GND_net), .CO(n32221));
    SB_LUT4 add_4609_14_lut (.I0(GND_net), .I1(n9258[11]), .I2(GND_net), 
            .I3(n32219), .O(n9241[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4587_15 (.CI(n31977), .I0(n8961[12]), .I1(GND_net), .CO(n31978));
    SB_CARRY add_4609_14 (.CI(n32219), .I0(n9258[11]), .I1(GND_net), .CO(n32220));
    SB_LUT4 add_4609_13_lut (.I0(GND_net), .I1(n9258[10]), .I2(GND_net), 
            .I3(n32218), .O(n9241[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4587_14_lut (.I0(GND_net), .I1(n8961[11]), .I2(GND_net), 
            .I3(n31976), .O(n8944[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4587_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_13 (.CI(n32218), .I0(n9258[10]), .I1(GND_net), .CO(n32219));
    SB_LUT4 add_4609_12_lut (.I0(GND_net), .I1(n9258[9]), .I2(GND_net), 
            .I3(n32217), .O(n9241[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_628_15_lut (.I0(GND_net), .I1(n2942[13]), .I2(n2967[13]), 
            .I3(n30367), .O(duty_23__N_3478[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_9_lut (.I0(GND_net), .I1(motor_state[7]), 
            .I2(n1_adj_3898[7]), .I3(n30507), .O(\PID_CONTROLLER.err_23__N_3379 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_12 (.CI(n32217), .I0(n9258[9]), .I1(GND_net), .CO(n32218));
    SB_LUT4 add_4609_11_lut (.I0(GND_net), .I1(n9258[8]), .I2(GND_net), 
            .I3(n32216), .O(n9241[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_11 (.CI(n32216), .I0(n9258[8]), .I1(GND_net), .CO(n32217));
    SB_LUT4 add_4609_10_lut (.I0(GND_net), .I1(n9258[7]), .I2(GND_net), 
            .I3(n32215), .O(n9241[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_15 (.CI(n30367), .I0(n2942[13]), .I1(n2967[13]), 
            .CO(n30368));
    SB_CARRY state_23__I_0_add_2_9 (.CI(n30507), .I0(motor_state[7]), .I1(n1_adj_3898[7]), 
            .CO(n30508));
    SB_LUT4 add_628_14_lut (.I0(GND_net), .I1(n2942[12]), .I2(n2967[12]), 
            .I3(n30366), .O(duty_23__N_3478[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4587_14 (.CI(n31976), .I0(n8961[11]), .I1(GND_net), .CO(n31977));
    SB_LUT4 add_4587_13_lut (.I0(GND_net), .I1(n8961[10]), .I2(GND_net), 
            .I3(n31975), .O(n8944[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4587_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_8_lut (.I0(GND_net), .I1(motor_state[6]), 
            .I2(n1_adj_3898[6]), .I3(n30506), .O(\PID_CONTROLLER.err_23__N_3379 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_8 (.CI(n30506), .I0(motor_state[6]), .I1(n1_adj_3898[6]), 
            .CO(n30507));
    SB_LUT4 state_23__I_0_add_2_7_lut (.I0(GND_net), .I1(motor_state[5]), 
            .I2(n1_adj_3898[5]), .I3(n30505), .O(\PID_CONTROLLER.err_23__N_3379 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4587_13 (.CI(n31975), .I0(n8961[10]), .I1(GND_net), .CO(n31976));
    SB_CARRY add_4609_10 (.CI(n32215), .I0(n9258[7]), .I1(GND_net), .CO(n32216));
    SB_LUT4 add_4587_12_lut (.I0(GND_net), .I1(n8961[9]), .I2(GND_net), 
            .I3(n31974), .O(n8944[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4587_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_7 (.CI(n30505), .I0(motor_state[5]), .I1(n1_adj_3898[5]), 
            .CO(n30506));
    SB_LUT4 add_4609_9_lut (.I0(GND_net), .I1(n9258[6]), .I2(GND_net), 
            .I3(n32214), .O(n9241[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4587_12 (.CI(n31974), .I0(n8961[9]), .I1(GND_net), .CO(n31975));
    SB_LUT4 add_4587_11_lut (.I0(GND_net), .I1(n8961[8]), .I2(GND_net), 
            .I3(n31973), .O(n8944[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4587_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4587_11 (.CI(n31973), .I0(n8961[8]), .I1(GND_net), .CO(n31974));
    SB_LUT4 add_4587_10_lut (.I0(GND_net), .I1(n8961[7]), .I2(GND_net), 
            .I3(n31972), .O(n8944[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4587_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_9 (.CI(n32214), .I0(n9258[6]), .I1(GND_net), .CO(n32215));
    SB_LUT4 add_4609_8_lut (.I0(GND_net), .I1(n9258[5]), .I2(n536), .I3(n32213), 
            .O(n9241[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_8 (.CI(n32213), .I0(n9258[5]), .I1(n536), .CO(n32214));
    SB_LUT4 add_4609_7_lut (.I0(GND_net), .I1(n9258[4]), .I2(n463), .I3(n32212), 
            .O(n9241[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_7 (.CI(n32212), .I0(n9258[4]), .I1(n463), .CO(n32213));
    SB_LUT4 add_4609_6_lut (.I0(GND_net), .I1(n9258[3]), .I2(n390), .I3(n32211), 
            .O(n9241[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_6 (.CI(n32211), .I0(n9258[3]), .I1(n390), .CO(n32212));
    SB_CARRY add_4587_10 (.CI(n31972), .I0(n8961[7]), .I1(GND_net), .CO(n31973));
    SB_LUT4 add_4609_5_lut (.I0(GND_net), .I1(n9258[2]), .I2(n317), .I3(n32210), 
            .O(n9241[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_5 (.CI(n32210), .I0(n9258[2]), .I1(n317), .CO(n32211));
    SB_LUT4 add_4609_4_lut (.I0(GND_net), .I1(n9258[1]), .I2(n244), .I3(n32209), 
            .O(n9241[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_14 (.CI(n30366), .I0(n2942[12]), .I1(n2967[12]), 
            .CO(n30367));
    SB_LUT4 add_4587_9_lut (.I0(GND_net), .I1(n8961[6]), .I2(GND_net), 
            .I3(n31971), .O(n8944[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4587_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4609_4 (.CI(n32209), .I0(n9258[1]), .I1(n244), .CO(n32210));
    SB_CARRY add_4587_9 (.CI(n31971), .I0(n8961[6]), .I1(GND_net), .CO(n31972));
    SB_LUT4 add_4587_8_lut (.I0(GND_net), .I1(n8961[5]), .I2(n536_adj_3859), 
            .I3(n31970), .O(n8944[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4587_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_628_13_lut (.I0(GND_net), .I1(n2942[11]), .I2(n2967[11]), 
            .I3(n30365), .O(duty_23__N_3478[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4587_8 (.CI(n31970), .I0(n8961[5]), .I1(n536_adj_3859), 
            .CO(n31971));
    SB_LUT4 add_4609_3_lut (.I0(GND_net), .I1(n9258[0]), .I2(n171), .I3(n32208), 
            .O(n9241[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4587_7_lut (.I0(GND_net), .I1(n8961[4]), .I2(n463_adj_3860), 
            .I3(n31969), .O(n8944[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4587_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4587_7 (.CI(n31969), .I0(n8961[4]), .I1(n463_adj_3860), 
            .CO(n31970));
    SB_CARRY add_4609_3 (.CI(n32208), .I0(n9258[0]), .I1(n171), .CO(n32209));
    SB_LUT4 add_4609_2_lut (.I0(GND_net), .I1(n29_adj_3861), .I2(n98), 
            .I3(GND_net), .O(n9241[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4609_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_13 (.CI(n30365), .I0(n2942[11]), .I1(n2967[11]), 
            .CO(n30366));
    SB_CARRY add_4609_2 (.CI(GND_net), .I0(n29_adj_3861), .I1(n98), .CO(n32208));
    SB_LUT4 state_23__I_0_add_2_6_lut (.I0(GND_net), .I1(motor_state[4]), 
            .I2(n1_adj_3898[4]), .I3(n30504), .O(\PID_CONTROLLER.err_23__N_3379 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4587_6_lut (.I0(GND_net), .I1(n8961[3]), .I2(n390_adj_3863), 
            .I3(n31968), .O(n8944[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4587_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_628_12_lut (.I0(GND_net), .I1(n2942[10]), .I2(n2967[10]), 
            .I3(n30364), .O(duty_23__N_3478[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4608_17_lut (.I0(GND_net), .I1(n9241[14]), .I2(GND_net), 
            .I3(n32207), .O(n9223[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_12 (.CI(n30364), .I0(n2942[10]), .I1(n2967[10]), 
            .CO(n30365));
    SB_LUT4 add_628_11_lut (.I0(GND_net), .I1(n2942[9]), .I2(n2967[9]), 
            .I3(n30363), .O(duty_23__N_3478[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4608_16_lut (.I0(GND_net), .I1(n9241[13]), .I2(GND_net), 
            .I3(n32206), .O(n9223[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4608_16 (.CI(n32206), .I0(n9241[13]), .I1(GND_net), .CO(n32207));
    SB_CARRY add_4587_6 (.CI(n31968), .I0(n8961[3]), .I1(n390_adj_3863), 
            .CO(n31969));
    SB_LUT4 add_4608_15_lut (.I0(GND_net), .I1(n9241[12]), .I2(GND_net), 
            .I3(n32205), .O(n9223[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4608_15 (.CI(n32205), .I0(n9241[12]), .I1(GND_net), .CO(n32206));
    SB_LUT4 add_4587_5_lut (.I0(GND_net), .I1(n8961[2]), .I2(n317_adj_3864), 
            .I3(n31967), .O(n8944[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4587_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_11 (.CI(n30363), .I0(n2942[9]), .I1(n2967[9]), .CO(n30364));
    SB_LUT4 add_4608_14_lut (.I0(GND_net), .I1(n9241[11]), .I2(GND_net), 
            .I3(n32204), .O(n9223[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_628_10_lut (.I0(GND_net), .I1(n2942[8]), .I2(n2967[8]), 
            .I3(n30362), .O(duty_23__N_3478[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4608_14 (.CI(n32204), .I0(n9241[11]), .I1(GND_net), .CO(n32205));
    SB_CARRY add_4587_5 (.CI(n31967), .I0(n8961[2]), .I1(n317_adj_3864), 
            .CO(n31968));
    SB_LUT4 add_4608_13_lut (.I0(GND_net), .I1(n9241[10]), .I2(GND_net), 
            .I3(n32203), .O(n9223[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4608_13 (.CI(n32203), .I0(n9241[10]), .I1(GND_net), .CO(n32204));
    SB_LUT4 add_4608_12_lut (.I0(GND_net), .I1(n9241[9]), .I2(GND_net), 
            .I3(n32202), .O(n9223[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4608_12 (.CI(n32202), .I0(n9241[9]), .I1(GND_net), .CO(n32203));
    SB_LUT4 add_4587_4_lut (.I0(GND_net), .I1(n8961[1]), .I2(n244_adj_3865), 
            .I3(n31966), .O(n8944[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4587_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4587_4 (.CI(n31966), .I0(n8961[1]), .I1(n244_adj_3865), 
            .CO(n31967));
    SB_LUT4 add_4587_3_lut (.I0(GND_net), .I1(n8961[0]), .I2(n171_adj_3866), 
            .I3(n31965), .O(n8944[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4587_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4587_3 (.CI(n31965), .I0(n8961[0]), .I1(n171_adj_3866), 
            .CO(n31966));
    SB_LUT4 add_4587_2_lut (.I0(GND_net), .I1(n29_adj_3867), .I2(n98_adj_3868), 
            .I3(GND_net), .O(n8944[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4587_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_10 (.CI(n30362), .I0(n2942[8]), .I1(n2967[8]), .CO(n30363));
    SB_CARRY add_4587_2 (.CI(GND_net), .I0(n29_adj_3867), .I1(n98_adj_3868), 
            .CO(n31965));
    SB_CARRY state_23__I_0_add_2_6 (.CI(n30504), .I0(motor_state[4]), .I1(n1_adj_3898[4]), 
            .CO(n30505));
    SB_LUT4 add_4608_11_lut (.I0(GND_net), .I1(n9241[8]), .I2(GND_net), 
            .I3(n32201), .O(n9223[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4586_17_lut (.I0(GND_net), .I1(n8944[14]), .I2(GND_net), 
            .I3(n31964), .O(n8926[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4608_11 (.CI(n32201), .I0(n9241[8]), .I1(GND_net), .CO(n32202));
    SB_LUT4 add_4586_16_lut (.I0(GND_net), .I1(n8944[13]), .I2(GND_net), 
            .I3(n31963), .O(n8926[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_628_9_lut (.I0(GND_net), .I1(n2942[7]), .I2(n2967[7]), 
            .I3(n30361), .O(duty_23__N_3478[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_5_lut (.I0(GND_net), .I1(motor_state[3]), 
            .I2(n1_adj_3898[3]), .I3(n30503), .O(\PID_CONTROLLER.err_23__N_3379 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_9 (.CI(n30361), .I0(n2942[7]), .I1(n2967[7]), .CO(n30362));
    SB_LUT4 add_628_8_lut (.I0(GND_net), .I1(n2942[6]), .I2(n2967[6]), 
            .I3(n30360), .O(duty_23__N_3478[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_8 (.CI(n30360), .I0(n2942[6]), .I1(n2967[6]), .CO(n30361));
    SB_CARRY add_4586_16 (.CI(n31963), .I0(n8944[13]), .I1(GND_net), .CO(n31964));
    SB_LUT4 add_4608_10_lut (.I0(GND_net), .I1(n9241[7]), .I2(GND_net), 
            .I3(n32200), .O(n9223[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4586_15_lut (.I0(GND_net), .I1(n8944[12]), .I2(GND_net), 
            .I3(n31962), .O(n8926[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_5 (.CI(n30503), .I0(motor_state[3]), .I1(n1_adj_3898[3]), 
            .CO(n30504));
    SB_LUT4 add_628_7_lut (.I0(GND_net), .I1(n2942[5]), .I2(n2967[5]), 
            .I3(n30359), .O(duty_23__N_3478[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_7 (.CI(n30359), .I0(n2942[5]), .I1(n2967[5]), .CO(n30360));
    SB_LUT4 state_23__I_0_add_2_4_lut (.I0(GND_net), .I1(motor_state[2]), 
            .I2(n1_adj_3898[2]), .I3(n30502), .O(\PID_CONTROLLER.err_23__N_3379 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4608_10 (.CI(n32200), .I0(n9241[7]), .I1(GND_net), .CO(n32201));
    SB_CARRY add_4586_15 (.CI(n31962), .I0(n8944[12]), .I1(GND_net), .CO(n31963));
    SB_CARRY state_23__I_0_add_2_4 (.CI(n30502), .I0(motor_state[2]), .I1(n1_adj_3898[2]), 
            .CO(n30503));
    SB_LUT4 add_628_6_lut (.I0(GND_net), .I1(n2942[4]), .I2(n2967[4]), 
            .I3(n30358), .O(duty_23__N_3478[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4608_9_lut (.I0(GND_net), .I1(n9241[6]), .I2(GND_net), 
            .I3(n32199), .O(n9223[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4586_14_lut (.I0(GND_net), .I1(n8944[11]), .I2(GND_net), 
            .I3(n31961), .O(n8926[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_628_6 (.CI(n30358), .I0(n2942[4]), .I1(n2967[4]), .CO(n30359));
    SB_CARRY add_4586_14 (.CI(n31961), .I0(n8944[11]), .I1(GND_net), .CO(n31962));
    SB_CARRY add_4608_9 (.CI(n32199), .I0(n9241[6]), .I1(GND_net), .CO(n32200));
    SB_LUT4 add_4608_8_lut (.I0(GND_net), .I1(n9241[5]), .I2(n533_adj_3871), 
            .I3(n32198), .O(n9223[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4586_13_lut (.I0(GND_net), .I1(n8944[10]), .I2(GND_net), 
            .I3(n31960), .O(n8926[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4586_13 (.CI(n31960), .I0(n8944[10]), .I1(GND_net), .CO(n31961));
    SB_LUT4 state_23__I_0_add_2_3_lut (.I0(GND_net), .I1(motor_state[1]), 
            .I2(n1_adj_3898[1]), .I3(n30501), .O(\PID_CONTROLLER.err_23__N_3379 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_3 (.CI(n30501), .I0(motor_state[1]), .I1(n1_adj_3898[1]), 
            .CO(n30502));
    SB_LUT4 add_4586_12_lut (.I0(GND_net), .I1(n8944[9]), .I2(GND_net), 
            .I3(n31959), .O(n8926[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_2_lut (.I0(GND_net), .I1(motor_state[0]), 
            .I2(n1_adj_3898[0]), .I3(VCC_net), .O(\PID_CONTROLLER.err_23__N_3379 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_628_5_lut (.I0(GND_net), .I1(n2942[3]), .I2(n2967[3]), 
            .I3(n30357), .O(duty_23__N_3478[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_628_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_2 (.CI(VCC_net), .I0(motor_state[0]), .I1(n1_adj_3898[0]), 
            .CO(n30501));
    SB_CARRY add_4608_8 (.CI(n32198), .I0(n9241[5]), .I1(n533_adj_3871), 
            .CO(n32199));
    SB_CARRY add_4586_12 (.CI(n31959), .I0(n8944[9]), .I1(GND_net), .CO(n31960));
    SB_LUT4 add_4586_11_lut (.I0(GND_net), .I1(n8944[8]), .I2(GND_net), 
            .I3(n31958), .O(n8926[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4586_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4608_7_lut (.I0(GND_net), .I1(n9241[4]), .I2(n460), .I3(n32197), 
            .O(n9223[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4608_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_3736));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3735));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_3734));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_3733));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_3732));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_3731));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_3730));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_3729));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[2]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_3698));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3697));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_3696));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_3695));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_3694));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_3693));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_3691));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_3690));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_3689));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[3]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[4]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25086_2_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\Kp[1] ), .I3(\PID_CONTROLLER.err [19]), .O(n9076[0]));   // verilog/motorControl.v(42[17:23])
    defparam i25086_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3897[5]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17_adj_3874));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_3875));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_3876));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36251_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n43376));
    defparam i36251_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i36213_3_lut (.I0(n11_adj_3876), .I1(n9_adj_3875), .I2(n43376), 
            .I3(GND_net), .O(n43337));
    defparam i36213_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_346_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n46698));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_346_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i37256_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n46698), 
            .I2(IntegralLimit[7]), .I3(n43337), .O(n44381));
    defparam i37256_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i36790_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_3874), 
            .I2(IntegralLimit[9]), .I3(n44381), .O(n43915));
    defparam i36790_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_328_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n46680));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_328_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36704_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_3874), 
            .I2(IntegralLimit[9]), .I3(n9_adj_3875), .O(n43829));
    defparam i36704_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i36694_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n46680), 
            .I2(IntegralLimit[11]), .I3(n43829), .O(n43819));
    defparam i36694_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_321_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n46673));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_321_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36468_4_lut (.I0(n27_adj_3661), .I1(n15_adj_3679), .I2(n13_adj_3680), 
            .I3(n11_adj_3681), .O(n43593));
    defparam i36468_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i36493_4_lut (.I0(n21_adj_3676), .I1(n19_adj_3677), .I2(n17_adj_3678), 
            .I3(n9_adj_3683), .O(n43618));
    defparam i36493_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43_adj_3641), .I3(GND_net), 
            .O(n16_adj_3877));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i36422_2_lut (.I0(n43_adj_3641), .I1(n19_adj_3677), .I2(GND_net), 
            .I3(GND_net), .O(n43547));
    defparam i36422_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_3678), .I3(GND_net), 
            .O(n8_adj_3878));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_3877), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45_adj_3636), .I3(GND_net), 
            .O(n24_adj_3879));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i36531_2_lut (.I0(n7_adj_3687), .I1(n5_adj_3699), .I2(GND_net), 
            .I3(GND_net), .O(n43656));
    defparam i36531_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i37128_4_lut (.I0(n13_adj_3680), .I1(n11_adj_3681), .I2(n9_adj_3683), 
            .I3(n43656), .O(n44253));
    defparam i37128_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i37122_4_lut (.I0(n19_adj_3677), .I1(n17_adj_3678), .I2(n15_adj_3679), 
            .I3(n44253), .O(n44247));
    defparam i37122_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i37807_4_lut (.I0(n25_adj_3666), .I1(n23_adj_3671), .I2(n21_adj_3676), 
            .I3(n44247), .O(n44932));
    defparam i37807_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i37384_4_lut (.I0(n31_adj_3655), .I1(n29_adj_3659), .I2(n27_adj_3661), 
            .I3(n44932), .O(n44509));
    defparam i37384_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i37893_4_lut (.I0(n37_adj_3647), .I1(n35_adj_3650), .I2(n33_adj_3652), 
            .I3(n44509), .O(n45018));
    defparam i37893_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36794_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n46698), 
            .I2(IntegralLimit[7]), .I3(n11_adj_3876), .O(n43919));
    defparam i36794_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_315_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n46667));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_315_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i36620_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n46667), 
            .I2(IntegralLimit[14]), .I3(n43919), .O(n43745));
    defparam i36620_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_309_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n46661));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_309_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_3880));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36578_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n43703));
    defparam i36578_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_333_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n46685));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_333_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_3881));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_3880), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30_adj_3882));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i37452_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n46680), 
            .I2(IntegralLimit[11]), .I3(n43915), .O(n44577));
    defparam i37452_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i35962_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n46673), 
            .I2(IntegralLimit[13]), .I3(n44577), .O(n43086));
    defparam i35962_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_313_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n46665));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_313_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i37194_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n46665), 
            .I2(IntegralLimit[15]), .I3(n43086), .O(n44319));
    defparam i37194_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_339_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n46691));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_339_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i37653_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n46691), 
            .I2(IntegralLimit[17]), .I3(n44319), .O(n44778));
    defparam i37653_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_304_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n46656));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_304_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i37897_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n46656), 
            .I2(IntegralLimit[19]), .I3(n44778), .O(n45022));
    defparam i37897_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_301_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n46653));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_301_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_3883));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36535_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n43660));
    defparam i36535_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_3883), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_3884));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_3885));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i37595_3_lut (.I0(n6_adj_3885), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n44720));   // verilog/motorControl.v(39[10:34])
    defparam i37595_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i37596_3_lut (.I0(n44720), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n44721));   // verilog/motorControl.v(39[10:34])
    defparam i37596_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36541_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n46673), 
            .I2(IntegralLimit[21]), .I3(n43819), .O(n43666));
    defparam i36541_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i37482_4_lut (.I0(n24_adj_3884), .I1(n8_adj_3886), .I2(n46651), 
            .I3(n43660), .O(n44607));   // verilog/motorControl.v(39[10:34])
    defparam i37482_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i37479_3_lut (.I0(n44721), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n44604));   // verilog/motorControl.v(39[10:34])
    defparam i37479_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3454 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3_adj_3737), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_3887));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 i37587_3_lut (.I0(n4_adj_3887), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27_adj_3661), .I3(GND_net), .O(n44712));   // verilog/motorControl.v(39[38:63])
    defparam i37587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37588_3_lut (.I0(n44712), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29_adj_3659), .I3(GND_net), .O(n44713));   // verilog/motorControl.v(39[38:63])
    defparam i37588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33_adj_3652), .I3(GND_net), 
            .O(n12_adj_3888));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i36443_2_lut (.I0(n33_adj_3652), .I1(n15_adj_3679), .I2(GND_net), 
            .I3(GND_net), .O(n43568));
    defparam i36443_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_3680), .I3(GND_net), 
            .O(n10_adj_3889));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_3888), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35_adj_3650), .I3(GND_net), 
            .O(n30_adj_3890));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i36446_4_lut (.I0(n33_adj_3652), .I1(n31_adj_3655), .I2(n29_adj_3659), 
            .I3(n43593), .O(n43571));
    defparam i36446_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37823_4_lut (.I0(n30_adj_3890), .I1(n10_adj_3889), .I2(n35_adj_3650), 
            .I3(n43568), .O(n44948));   // verilog/motorControl.v(39[38:63])
    defparam i37823_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36753_3_lut (.I0(n44713), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31_adj_3655), .I3(GND_net), .O(n43878));   // verilog/motorControl.v(39[38:63])
    defparam i36753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37957_4_lut (.I0(n43878), .I1(n44948), .I2(n35_adj_3650), 
            .I3(n43571), .O(n45082));   // verilog/motorControl.v(39[38:63])
    defparam i37957_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i37958_3_lut (.I0(n45082), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37_adj_3647), .I3(GND_net), .O(n45083));   // verilog/motorControl.v(39[38:63])
    defparam i37958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37944_3_lut (.I0(n45083), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39_adj_3645), .I3(GND_net), .O(n45069));   // verilog/motorControl.v(39[38:63])
    defparam i37944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_3687), .I3(GND_net), 
            .O(n6_adj_3891));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i37589_3_lut (.I0(n6_adj_3891), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_3676), .I3(GND_net), .O(n44714));   // verilog/motorControl.v(39[38:63])
    defparam i37589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37590_3_lut (.I0(n44714), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_3671), .I3(GND_net), .O(n44715));   // verilog/motorControl.v(39[38:63])
    defparam i37590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36425_4_lut (.I0(n43_adj_3641), .I1(n25_adj_3666), .I2(n23_adj_3671), 
            .I3(n43618), .O(n43550));
    defparam i36425_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37484_4_lut (.I0(n24_adj_3879), .I1(n8_adj_3878), .I2(n45_adj_3636), 
            .I3(n43547), .O(n44609));   // verilog/motorControl.v(39[38:63])
    defparam i37484_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36751_3_lut (.I0(n44715), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_3666), .I3(GND_net), .O(n43876));   // verilog/motorControl.v(39[38:63])
    defparam i36751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36429_4_lut (.I0(n43_adj_3641), .I1(n41_adj_3643), .I2(n39_adj_3645), 
            .I3(n45018), .O(n43554));
    defparam i36429_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i37863_4_lut (.I0(n43876), .I1(n44609), .I2(n45_adj_3636), 
            .I3(n43550), .O(n44988));   // verilog/motorControl.v(39[38:63])
    defparam i37863_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36759_3_lut (.I0(n45069), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41_adj_3643), .I3(GND_net), .O(n43884));   // verilog/motorControl.v(39[38:63])
    defparam i36759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i37865_4_lut (.I0(n43884), .I1(n44988), .I2(n45_adj_3636), 
            .I3(n43554), .O(n44990));   // verilog/motorControl.v(39[38:63])
    defparam i37865_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_3892));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i37593_3_lut (.I0(n4_adj_3892), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n44718));   // verilog/motorControl.v(39[10:34])
    defparam i37593_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i37594_3_lut (.I0(n44718), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n44719));   // verilog/motorControl.v(39[10:34])
    defparam i37594_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36583_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n46661), 
            .I2(IntegralLimit[16]), .I3(n43745), .O(n43708));
    defparam i36583_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i37821_4_lut (.I0(n30_adj_3882), .I1(n10_adj_3881), .I2(n46685), 
            .I3(n43703), .O(n44946));   // verilog/motorControl.v(39[10:34])
    defparam i37821_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i37481_3_lut (.I0(n44719), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n28));   // verilog/motorControl.v(39[10:34])
    defparam i37481_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i37953_4_lut (.I0(n28), .I1(n44946), .I2(n46685), .I3(n43708), 
            .O(n45078));   // verilog/motorControl.v(39[10:34])
    defparam i37953_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i37954_3_lut (.I0(n45078), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n45079));   // verilog/motorControl.v(39[10:34])
    defparam i37954_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i37948_3_lut (.I0(n45079), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n45073));   // verilog/motorControl.v(39[10:34])
    defparam i37948_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36543_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n46653), 
            .I2(IntegralLimit[21]), .I3(n45022), .O(n43668));
    defparam i36543_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_299_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n46651));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_299_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i37859_4_lut (.I0(n44604), .I1(n44607), .I2(n46651), .I3(n43666), 
            .O(n44984));   // verilog/motorControl.v(39[10:34])
    defparam i37859_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36749_3_lut (.I0(n45073), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n43874));   // verilog/motorControl.v(39[10:34])
    defparam i36749_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i37866_3_lut (.I0(n44990), .I1(\PID_CONTROLLER.integral_23__N_3454 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3453 ));   // verilog/motorControl.v(39[38:63])
    defparam i37866_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i37861_4_lut (.I0(n43874), .I1(n44984), .I2(n46651), .I3(n43668), 
            .O(n44986));   // verilog/motorControl.v(39[10:34])
    defparam i37861_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_840_4_lut  (.I0(n44986), .I1(\PID_CONTROLLER.integral_23__N_3453 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3451 ));   // verilog/motorControl.v(39[10:63])
    defparam \PID_CONTROLLER.integral_23__I_840_4_lut .LUT_INIT = 16'h80c8;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty[4]), .I1(n257[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_3717));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty[5]), .I1(n257[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_3719));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty[6]), .I1(n257[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_3718));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_3627));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3626));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_3623));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_3621));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_3619));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i1_1_lut (.I0(setpoint[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[0]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i2_1_lut (.I0(setpoint[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[1]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_3871));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_3886));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_626_i5_3_lut (.I0(n155[4]), .I1(n1[4]), .I2(n256), .I3(GND_net), 
            .O(n2967[4]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 state_23__I_0_inv_0_i3_1_lut (.I0(setpoint[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[2]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_626_i6_3_lut (.I0(n155[5]), .I1(n1[5]), .I2(n256), .I3(GND_net), 
            .O(n2967[5]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_626_i7_3_lut (.I0(n155[6]), .I1(n1[6]), .I2(n256), .I3(GND_net), 
            .O(n2967[6]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 state_23__I_0_inv_0_i4_1_lut (.I0(setpoint[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[3]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_626_i8_3_lut (.I0(n155[7]), .I1(n1[7]), .I2(n256), .I3(GND_net), 
            .O(n2967[7]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_3868));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_3867));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_3866));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_3865));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_626_i9_3_lut (.I0(n155[8]), .I1(n1[8]), .I2(n256), .I3(GND_net), 
            .O(n2967[8]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317_adj_3864));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_626_i10_3_lut (.I0(n155[9]), .I1(n1[9]), .I2(n256), .I3(GND_net), 
            .O(n2967[9]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_626_i11_3_lut (.I0(n155[10]), .I1(n1[10]), .I2(n256), 
            .I3(GND_net), .O(n2967[10]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_3614));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_3863));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i5_1_lut (.I0(setpoint[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[4]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_3861));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_3860));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_626_i12_3_lut (.I0(n155[11]), .I1(n1[11]), .I2(n256), 
            .I3(GND_net), .O(n2967[11]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3612));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536_adj_3859));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i6_1_lut (.I0(setpoint[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[5]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i7_1_lut (.I0(setpoint[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[6]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_626_i13_3_lut (.I0(n155[12]), .I1(n1[12]), .I2(n256), 
            .I3(GND_net), .O(n2967[12]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i8_1_lut (.I0(setpoint[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[7]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_626_i14_3_lut (.I0(n155[13]), .I1(n1[13]), .I2(n256), 
            .I3(GND_net), .O(n2967[13]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_3610));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_3855));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_3854));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_3853));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i9_1_lut (.I0(setpoint[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[8]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_626_i15_3_lut (.I0(n155[14]), .I1(n1[14]), .I2(n256), 
            .I3(GND_net), .O(n2967[14]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_3851));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_626_i16_3_lut (.I0(n155[15]), .I1(n1[15]), .I2(n256), 
            .I3(GND_net), .O(n2967[15]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 state_23__I_0_inv_0_i10_1_lut (.I0(setpoint[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[9]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_3849));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_626_i17_3_lut (.I0(n155[16]), .I1(n1[16]), .I2(n256), 
            .I3(GND_net), .O(n2967[16]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i11_1_lut (.I0(setpoint[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[10]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_3847));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i12_1_lut (.I0(setpoint[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[11]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i13_1_lut (.I0(setpoint[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[12]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_3842));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_3839));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_626_i18_3_lut (.I0(n155[17]), .I1(n1[17]), .I2(n256), 
            .I3(GND_net), .O(n2967[17]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_3836));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3835));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177_adj_3834));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_3833));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_3832));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3831));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i14_1_lut (.I0(setpoint[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[13]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_3829));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_3828));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_3827));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542_adj_3826));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_626_i19_3_lut (.I0(n155[18]), .I1(n1[18]), .I2(n256), 
            .I3(GND_net), .O(n2967[18]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_626_i20_3_lut (.I0(n155[19]), .I1(n1[19]), .I2(n256), 
            .I3(GND_net), .O(n2967[19]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 state_23__I_0_inv_0_i15_1_lut (.I0(setpoint[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[14]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_626_i21_3_lut (.I0(n155[20]), .I1(n1[20]), .I2(n256), 
            .I3(GND_net), .O(n2967[20]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i16_1_lut (.I0(setpoint[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[15]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i17_1_lut (.I0(setpoint[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[16]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i18_1_lut (.I0(setpoint[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[17]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_626_i22_3_lut (.I0(n155[21]), .I1(n1[21]), .I2(n256), 
            .I3(GND_net), .O(n2967[21]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25208_2_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(\Ki[1] ), .I3(\PID_CONTROLLER.integral [19]), .O(n9373[0]));   // verilog/motorControl.v(42[26:37])
    defparam i25208_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i36261_3_lut_4_lut (.I0(duty[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty[2]), .O(n43386));   // verilog/motorControl.v(46[19:35])
    defparam i36261_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(GND_net), .O(n6_adj_3724));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_3821));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_3820));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_3819));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253_adj_3818));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_3817));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_626_i4_3_lut (.I0(n155[3]), .I1(PWMLimit[3]), .I2(n256), 
            .I3(GND_net), .O(n2967[3]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i4_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_3816));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_3815));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_3814));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_3813));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_626_i23_3_lut (.I0(n155[22]), .I1(n1[22]), .I2(n256), 
            .I3(GND_net), .O(n2967[22]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_626_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i19_1_lut (.I0(setpoint[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[18]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i20_1_lut (.I0(setpoint[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[19]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_3810));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3809));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_3808));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i21_1_lut (.I0(setpoint[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[20]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_3806));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_3805));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_3804));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_3803));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_3802));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3801));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_3800));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_3799));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_3798));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_3797));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_3796));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_3795));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_3794));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_3793));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_3792));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_3791));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_3790));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i22_1_lut (.I0(setpoint[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[21]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_3784));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_3783));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_3782));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i23_1_lut (.I0(setpoint[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[22]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_3780));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_3779));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_3778));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_3777));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_3776));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i24_1_lut (.I0(setpoint[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_3898[23]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_3774));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_3773));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_3772));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_3771));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_3770));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_3769));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_3768));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_3767));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_3766));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_3765));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_3762));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_3761));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_3760));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_626_i24_3_lut_3_lut (.I0(PWMLimit[23]), .I1(n256), .I2(n42910), 
            .I3(GND_net), .O(n2967[23]));   // verilog/motorControl.v(47[19:28])
    defparam mux_626_i24_3_lut_3_lut.LUT_INIT = 16'h7474;
    SB_LUT4 i36139_2_lut_4_lut (.I0(duty[21]), .I1(n257[21]), .I2(duty[9]), 
            .I3(n257[9]), .O(n43263));
    defparam i36139_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i36169_2_lut_4_lut (.I0(duty[16]), .I1(n257[16]), .I2(duty[7]), 
            .I3(n257[7]), .O(n43293));
    defparam i36169_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_3757));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_3756));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_3755));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_3754));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_3753));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_3752));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414_adj_3751));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_3750));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487_adj_3749));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560_adj_3748));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_3747));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_3746));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i24_3_lut (.I0(duty_23__N_3478[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[23]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i23_3_lut (.I0(duty_23__N_3478[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[22]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i22_3_lut (.I0(duty_23__N_3478[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[21]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i21_3_lut (.I0(duty_23__N_3478[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[20]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i20_3_lut (.I0(duty_23__N_3478[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[19]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i19_3_lut (.I0(duty_23__N_3478[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[18]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i18_3_lut (.I0(duty_23__N_3478[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[17]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i17_3_lut (.I0(duty_23__N_3478[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[16]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i16_3_lut (.I0(duty_23__N_3478[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[15]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i15_3_lut (.I0(duty_23__N_3478[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[14]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i14_3_lut (.I0(duty_23__N_3478[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[13]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i13_3_lut (.I0(duty_23__N_3478[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[12]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i12_3_lut (.I0(duty_23__N_3478[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[11]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i11_3_lut (.I0(duty_23__N_3478[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[10]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i10_3_lut (.I0(duty_23__N_3478[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[9]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i9_3_lut (.I0(duty_23__N_3478[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[8]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i8_3_lut (.I0(duty_23__N_3478[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[7]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i7_3_lut (.I0(duty_23__N_3478[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[6]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i6_3_lut (.I0(duty_23__N_3478[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[5]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i5_3_lut (.I0(duty_23__N_3478[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[4]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i4_3_lut (.I0(duty_23__N_3478[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[3]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i3_3_lut (.I0(duty_23__N_3478[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3502), .I3(GND_net), .O(duty_23__N_3355[2]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_3745));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_3744));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(PWMLimit[8]), 
            .I3(GND_net), .O(n8_adj_3628));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36263_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(PWMLimit[9]), 
            .I3(duty[9]), .O(n43388));
    defparam i36263_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(duty[9]), .I1(duty[21]), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n16_adj_3624));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(PWMLimit[6]), 
            .I3(GND_net), .O(n10_adj_3630));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i36291_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(PWMLimit[7]), 
            .I3(duty[7]), .O(n43416));
    defparam i36291_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(duty[7]), .I1(duty[16]), .I2(PWMLimit[16]), 
            .I3(GND_net), .O(n12_adj_3620));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344_adj_3743));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i38742_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n45865));   // verilog/motorControl.v(37[14] 56[8])
    defparam i38742_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i25068_3_lut_4_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n4_adj_3893), .I3(n9076[1]), .O(n6));   // verilog/motorControl.v(42[17:23])
    defparam i25068_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_855 (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n9076[1]), .I3(n4_adj_3893), .O(n9069[2]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_855.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_856 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n9076[0]), .I3(n29997), .O(n9069[1]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_856.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417_adj_3742));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_857 (.I0(n6), .I1(\Kp[4] ), .I2(n9076[2]), .I3(\PID_CONTROLLER.err [18]), 
            .O(n9069[3]));   // verilog/motorControl.v(42[17:23])
    defparam i2_4_lut_adj_857.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_3741));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_3740));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25060_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n29997), .I3(n9076[0]), .O(n4_adj_3893));   // verilog/motorControl.v(42[17:23])
    defparam i25060_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i138_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204_adj_3894));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25049_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n29997));   // verilog/motorControl.v(42[17:23])
    defparam i25049_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i25140_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n9087[0]));   // verilog/motorControl.v(42[17:23])
    defparam i25140_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i25047_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n9069[0]));   // verilog/motorControl.v(42[17:23])
    defparam i25047_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i25130_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n30074), .I3(n9087[0]), .O(n4_adj_3568));   // verilog/motorControl.v(42[17:23])
    defparam i25130_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_10_i89_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131_adj_3895));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i42_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62_adj_3896));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_858 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n9087[0]), .I3(n30074), .O(n9082[1]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_858.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_859 (.I0(n62_adj_3896), .I1(n131_adj_3895), 
            .I2(n9082[0]), .I3(n204_adj_3894), .O(n9076[1]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_859.LUT_INIT = 16'h8778;
    SB_LUT4 i25099_3_lut_4_lut (.I0(n62_adj_3896), .I1(n131_adj_3895), .I2(n204_adj_3894), 
            .I3(n9082[0]), .O(n4));   // verilog/motorControl.v(42[17:23])
    defparam i25099_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i25117_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n9082[0]));   // verilog/motorControl.v(42[17:23])
    defparam i25117_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i25119_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n30074));   // verilog/motorControl.v(42[17:23])
    defparam i25119_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i2_4_lut_adj_860 (.I0(n4), .I1(\Kp[3] ), .I2(n9082[1]), .I3(\PID_CONTROLLER.err [19]), 
            .O(n9076[2]));   // verilog/motorControl.v(42[17:23])
    defparam i2_4_lut_adj_860.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490_adj_3739));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_861 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(\PID_CONTROLLER.err [23]), 
            .I3(\PID_CONTROLLER.err [20]), .O(n12));   // verilog/motorControl.v(42[17:23])
    defparam i2_4_lut_adj_861.LUT_INIT = 16'h9c50;
    
endmodule
//
// Verilog Description of module \pwm(32000000,20000,32000000,23,1) 
//

module \pwm(32000000,20000,32000000,23,1)  (pwm_setpoint, GND_net, \half_duty_new[0] , 
            CLK_c, PIN_19_c_0, n19420, \half_duty[0][2] , n19421, 
            \half_duty[0][3] , n19422, \half_duty[0][4] , n19423, \half_duty[0][5] , 
            n19424, \half_duty[0][6] , n19425, \half_duty[0][7] , n19414, 
            \half_duty[0][1] , n1111, VCC_net, \half_duty_new[1] , \half_duty[0][0] , 
            \half_duty_new[2] , \half_duty_new[3] , \half_duty_new[4] , 
            \half_duty_new[5] , \half_duty_new[6] , \half_duty_new[7] , 
            n18810) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input [22:0]pwm_setpoint;
    input GND_net;
    output \half_duty_new[0] ;
    input CLK_c;
    output PIN_19_c_0;
    input n19420;
    output \half_duty[0][2] ;
    input n19421;
    output \half_duty[0][3] ;
    input n19422;
    output \half_duty[0][4] ;
    input n19423;
    output \half_duty[0][5] ;
    input n19424;
    output \half_duty[0][6] ;
    input n19425;
    output \half_duty[0][7] ;
    input n19414;
    output \half_duty[0][1] ;
    output n1111;
    input VCC_net;
    output \half_duty_new[1] ;
    output \half_duty[0][0] ;
    output \half_duty_new[2] ;
    output \half_duty_new[3] ;
    output \half_duty_new[4] ;
    output \half_duty_new[5] ;
    output \half_duty_new[6] ;
    output \half_duty_new[7] ;
    input n18810;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [22:0]n5875;
    
    wire n30577, n30578;
    wire [9:0]half_duty_new_9__N_664;
    
    wire pwm_out_0__N_582, n38158, n30576, n30575, n30574, n30573, 
        n30572, n30571;
    wire [10:0]n49;
    
    wire pause_counter_0__N_612;
    wire [10:0]\count[0] ;   // vhdl/pwm.vhd(51[11:16])
    
    wire pause_counter_0, n38146, n30300, pwm_out_0__N_586, n30299, 
        n10, n30298, n9, n30297, n8;
    wire [10:0]pwm_out_0__N_587;
    
    wire n30296, n4, n5, n3, n12, n1, n39870, n6, n2, n10_adj_3561, 
        n7, n9_adj_3562, n13, n12_adj_3563, n18, n3_adj_3564, n16, 
        n20, n30295, n30294, n30293, n30292, n30291, n30290, n31184, 
        n31183, n31182, n31181, n31180, n31179, n31178, n31177, 
        n31176, n31175, n30613, n30612, n30611, n30610, n30609, 
        n30608, n30607, n30606, n30605, n30604, n30603, n30602, 
        n30601, n30600, n30599, n30598, n30597, n30596, n30595, 
        n30594, n30593, n30592, n30591, n30590, n30589, n30588, 
        n30587, n30586, n30585, n30584, n30583, n30582, n30581, 
        n30580, n30579, n20_adj_3565, n19, n6_adj_3566;
    
    SB_LUT4 add_2004_9_lut (.I0(GND_net), .I1(pwm_setpoint[7]), .I2(pwm_setpoint[11]), 
            .I3(n30577), .O(n5875[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_9 (.CI(n30577), .I0(pwm_setpoint[7]), .I1(pwm_setpoint[11]), 
            .CO(n30578));
    SB_DFF half_duty_new_i1 (.Q(\half_duty_new[0] ), .C(CLK_c), .D(half_duty_new_9__N_664[0]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFFE pwm_out_0__39 (.Q(PIN_19_c_0), .C(CLK_c), .E(n38158), .D(pwm_out_0__N_582));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 add_2004_8_lut (.I0(GND_net), .I1(pwm_setpoint[6]), .I2(pwm_setpoint[10]), 
            .I3(n30576), .O(n5875[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_8 (.CI(n30576), .I0(pwm_setpoint[6]), .I1(pwm_setpoint[10]), 
            .CO(n30577));
    SB_LUT4 add_2004_7_lut (.I0(GND_net), .I1(pwm_setpoint[5]), .I2(pwm_setpoint[9]), 
            .I3(n30575), .O(n5875[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_7 (.CI(n30575), .I0(pwm_setpoint[5]), .I1(pwm_setpoint[9]), 
            .CO(n30576));
    SB_LUT4 add_2004_6_lut (.I0(GND_net), .I1(pwm_setpoint[4]), .I2(pwm_setpoint[8]), 
            .I3(n30574), .O(n5875[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_6 (.CI(n30574), .I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .CO(n30575));
    SB_LUT4 add_2004_5_lut (.I0(GND_net), .I1(pwm_setpoint[3]), .I2(pwm_setpoint[7]), 
            .I3(n30573), .O(n5875[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_5 (.CI(n30573), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[7]), 
            .CO(n30574));
    SB_DFF half_duty_0___i3 (.Q(\half_duty[0][2] ), .C(CLK_c), .D(n19420));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i4 (.Q(\half_duty[0][3] ), .C(CLK_c), .D(n19421));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i5 (.Q(\half_duty[0][4] ), .C(CLK_c), .D(n19422));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i6 (.Q(\half_duty[0][5] ), .C(CLK_c), .D(n19423));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i7 (.Q(\half_duty[0][6] ), .C(CLK_c), .D(n19424));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i8 (.Q(\half_duty[0][7] ), .C(CLK_c), .D(n19425));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 add_2004_4_lut (.I0(GND_net), .I1(pwm_setpoint[2]), .I2(pwm_setpoint[6]), 
            .I3(n30572), .O(n5875[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF half_duty_0___i2 (.Q(\half_duty[0][1] ), .C(CLK_c), .D(n19414));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_CARRY add_2004_4 (.CI(n30572), .I0(pwm_setpoint[2]), .I1(pwm_setpoint[6]), 
            .CO(n30573));
    SB_LUT4 add_2004_3_lut (.I0(GND_net), .I1(pwm_setpoint[1]), .I2(pwm_setpoint[5]), 
            .I3(n30571), .O(n5875[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_3 (.CI(n30571), .I0(pwm_setpoint[1]), .I1(pwm_setpoint[5]), 
            .CO(n30572));
    SB_LUT4 add_2004_2_lut (.I0(GND_net), .I1(pwm_setpoint[0]), .I2(pwm_setpoint[4]), 
            .I3(GND_net), .O(n5875[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_2 (.CI(GND_net), .I0(pwm_setpoint[0]), .I1(pwm_setpoint[4]), 
            .CO(n30571));
    SB_DFFESR count_0__1148__i10 (.Q(\count[0] [10]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[10]), .R(n1111));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1148__i9 (.Q(\count[0] [9]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[9]), .R(n1111));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1148__i8 (.Q(\count[0] [8]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[8]), .R(n1111));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1148__i7 (.Q(\count[0] [7]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[7]), .R(n1111));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1148__i6 (.Q(\count[0] [6]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[6]), .R(n1111));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1148__i5 (.Q(\count[0] [5]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[5]), .R(n1111));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1148__i4 (.Q(\count[0] [4]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[4]), .R(n1111));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1148__i3 (.Q(\count[0] [3]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[3]), .R(n1111));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1148__i2 (.Q(\count[0] [2]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[2]), .R(n1111));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1148__i1 (.Q(\count[0] [1]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[1]), .R(n1111));   // vhdl/pwm.vhd(77[18:26])
    SB_LUT4 i38727_2_lut (.I0(pause_counter_0), .I1(pwm_out_0__N_582), .I2(GND_net), 
            .I3(GND_net), .O(n38146));
    defparam i38727_2_lut.LUT_INIT = 16'h1111;
    SB_DFF pause_counter_0__38 (.Q(pause_counter_0), .C(CLK_c), .D(n38146));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFFESR count_0__1148__i0 (.Q(\count[0] [0]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[0]), .R(n1111));   // vhdl/pwm.vhd(77[18:26])
    SB_CARRY pwm_out_0__I_20_13 (.CI(n30300), .I0(GND_net), .I1(VCC_net), 
            .CO(pwm_out_0__N_586));
    SB_CARRY pwm_out_0__I_20_12 (.CI(n30299), .I0(VCC_net), .I1(VCC_net), 
            .CO(n30300));
    SB_LUT4 pwm_out_0__I_20_11_lut (.I0(\count[0] [9]), .I1(VCC_net), .I2(VCC_net), 
            .I3(n30298), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_11 (.CI(n30298), .I0(VCC_net), .I1(VCC_net), 
            .CO(n30299));
    SB_LUT4 pwm_out_0__I_20_10_lut (.I0(\count[0] [8]), .I1(GND_net), .I2(VCC_net), 
            .I3(n30297), .O(n9)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_10_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_10 (.CI(n30297), .I0(GND_net), .I1(VCC_net), 
            .CO(n30298));
    SB_LUT4 pause_counter_0__I_0_48_1_lut (.I0(pause_counter_0), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pause_counter_0__N_612));   // vhdl/pwm.vhd(72[7:27])
    defparam pause_counter_0__I_0_48_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 pwm_out_0__I_20_9_lut (.I0(\count[0] [7]), .I1(GND_net), .I2(pwm_out_0__N_587[7]), 
            .I3(n30296), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_9 (.CI(n30296), .I0(GND_net), .I1(pwm_out_0__N_587[7]), 
            .CO(n30297));
    SB_DFF half_duty_new_i2 (.Q(\half_duty_new[1] ), .C(CLK_c), .D(half_duty_new_9__N_664[1]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 i5_4_lut (.I0(n4), .I1(n5), .I2(n3), .I3(pwm_out_0__N_586), 
            .O(n12));   // vhdl/pwm.vhd(84[11:43])
    defparam i5_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i6_4_lut (.I0(n1), .I1(n12), .I2(n8), .I3(n9), .O(n39870));   // vhdl/pwm.vhd(84[11:43])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_4_lut (.I0(\count[0] [10]), .I1(n39870), .I2(n6), .I3(n2), 
            .O(n10_adj_3561));   // vhdl/pwm.vhd(84[11:43])
    defparam i4_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 i3_2_lut (.I0(n7), .I1(n10), .I2(GND_net), .I3(GND_net), 
            .O(n9_adj_3562));   // vhdl/pwm.vhd(84[11:43])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i38012_4_lut (.I0(n9_adj_3562), .I1(pause_counter_0), .I2(pwm_out_0__N_582), 
            .I3(n10_adj_3561), .O(n38158));
    defparam i38012_4_lut.LUT_INIT = 16'h0313;
    SB_LUT4 i2_4_lut (.I0(\half_duty[0][6] ), .I1(\half_duty[0][5] ), .I2(\count[0] [6]), 
            .I3(\count[0] [5]), .O(n13));   // vhdl/pwm.vhd(80[8:31])
    defparam i2_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_3_lut (.I0(\half_duty[0][3] ), .I1(\count[0] [10]), .I2(\count[0] [3]), 
            .I3(GND_net), .O(n12_adj_3563));   // vhdl/pwm.vhd(80[8:31])
    defparam i1_3_lut.LUT_INIT = 16'hdede;
    SB_LUT4 i7_4_lut (.I0(n13), .I1(\half_duty[0][7] ), .I2(\count[0] [9]), 
            .I3(\count[0] [7]), .O(n18));   // vhdl/pwm.vhd(80[8:31])
    defparam i7_4_lut.LUT_INIT = 16'hfbfe;
    SB_LUT4 half_duty_0__9__I_0_47_i3_2_lut (.I0(\half_duty[0][2] ), .I1(\count[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3564));   // vhdl/pwm.vhd(80[8:31])
    defparam half_duty_0__9__I_0_47_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_842 (.I0(\half_duty[0][1] ), .I1(\half_duty[0][0] ), 
            .I2(\count[0] [1]), .I3(\count[0] [0]), .O(n16));   // vhdl/pwm.vhd(80[8:31])
    defparam i5_4_lut_adj_842.LUT_INIT = 16'h7bde;
    SB_LUT4 i9_4_lut (.I0(\half_duty[0][4] ), .I1(n18), .I2(n12_adj_3563), 
            .I3(\count[0] [4]), .O(n20));   // vhdl/pwm.vhd(80[8:31])
    defparam i9_4_lut.LUT_INIT = 16'hfdfe;
    SB_LUT4 i10_4_lut (.I0(\count[0] [8]), .I1(n20), .I2(n16), .I3(n3_adj_3564), 
            .O(pwm_out_0__N_582));   // vhdl/pwm.vhd(80[8:31])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF half_duty_new_i3 (.Q(\half_duty_new[2] ), .C(CLK_c), .D(half_duty_new_9__N_664[2]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i4 (.Q(\half_duty_new[3] ), .C(CLK_c), .D(half_duty_new_9__N_664[3]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i5 (.Q(\half_duty_new[4] ), .C(CLK_c), .D(half_duty_new_9__N_664[4]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i6 (.Q(\half_duty_new[5] ), .C(CLK_c), .D(half_duty_new_9__N_664[5]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i7 (.Q(\half_duty_new[6] ), .C(CLK_c), .D(half_duty_new_9__N_664[6]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i8 (.Q(\half_duty_new[7] ), .C(CLK_c), .D(half_duty_new_9__N_664[7]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 pwm_out_0__I_20_8_lut (.I0(\count[0] [6]), .I1(VCC_net), .I2(pwm_out_0__N_587[6]), 
            .I3(n30295), .O(n7)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_8 (.CI(n30295), .I0(VCC_net), .I1(pwm_out_0__N_587[6]), 
            .CO(n30296));
    SB_LUT4 pwm_out_0__I_20_7_lut (.I0(\count[0] [5]), .I1(GND_net), .I2(pwm_out_0__N_587[5]), 
            .I3(n30294), .O(n6)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_7 (.CI(n30294), .I0(GND_net), .I1(pwm_out_0__N_587[5]), 
            .CO(n30295));
    SB_LUT4 pwm_out_0__I_20_6_lut (.I0(\count[0] [4]), .I1(GND_net), .I2(pwm_out_0__N_587[4]), 
            .I3(n30293), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_6 (.CI(n30293), .I0(GND_net), .I1(pwm_out_0__N_587[4]), 
            .CO(n30294));
    SB_LUT4 pwm_out_0__I_20_5_lut (.I0(\count[0] [3]), .I1(GND_net), .I2(pwm_out_0__N_587[3]), 
            .I3(n30292), .O(n4)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_5 (.CI(n30292), .I0(GND_net), .I1(pwm_out_0__N_587[3]), 
            .CO(n30293));
    SB_LUT4 pwm_out_0__I_20_4_lut (.I0(\count[0] [2]), .I1(GND_net), .I2(pwm_out_0__N_587[2]), 
            .I3(n30291), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_4 (.CI(n30291), .I0(GND_net), .I1(pwm_out_0__N_587[2]), 
            .CO(n30292));
    SB_LUT4 pwm_out_0__I_20_3_lut (.I0(\count[0] [1]), .I1(GND_net), .I2(pwm_out_0__N_587[1]), 
            .I3(n30290), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_3_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_3 (.CI(n30290), .I0(GND_net), .I1(pwm_out_0__N_587[1]), 
            .CO(n30291));
    SB_LUT4 pwm_out_0__I_20_2_lut (.I0(\count[0] [0]), .I1(GND_net), .I2(pwm_out_0__N_587[0]), 
            .I3(VCC_net), .O(n1)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_2_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_out_0__N_587[0]), 
            .CO(n30290));
    SB_DFF half_duty_0___i1 (.Q(\half_duty[0][0] ), .C(CLK_c), .D(n18810));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 count_0__1148_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [10]), 
            .I3(n31184), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1148_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 count_0__1148_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [9]), 
            .I3(n31183), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1148_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1148_add_4_11 (.CI(n31183), .I0(GND_net), .I1(\count[0] [9]), 
            .CO(n31184));
    SB_LUT4 count_0__1148_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [8]), 
            .I3(n31182), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1148_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1148_add_4_10 (.CI(n31182), .I0(GND_net), .I1(\count[0] [8]), 
            .CO(n31183));
    SB_LUT4 count_0__1148_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [7]), 
            .I3(n31181), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1148_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1148_add_4_9 (.CI(n31181), .I0(GND_net), .I1(\count[0] [7]), 
            .CO(n31182));
    SB_LUT4 count_0__1148_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [6]), 
            .I3(n31180), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1148_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1148_add_4_8 (.CI(n31180), .I0(GND_net), .I1(\count[0] [6]), 
            .CO(n31181));
    SB_LUT4 count_0__1148_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [5]), 
            .I3(n31179), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1148_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1148_add_4_7 (.CI(n31179), .I0(GND_net), .I1(\count[0] [5]), 
            .CO(n31180));
    SB_LUT4 count_0__1148_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [4]), 
            .I3(n31178), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1148_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1148_add_4_6 (.CI(n31178), .I0(GND_net), .I1(\count[0] [4]), 
            .CO(n31179));
    SB_LUT4 count_0__1148_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [3]), 
            .I3(n31177), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1148_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1148_add_4_5 (.CI(n31177), .I0(GND_net), .I1(\count[0] [3]), 
            .CO(n31178));
    SB_LUT4 count_0__1148_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [2]), 
            .I3(n31176), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1148_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1148_add_4_4 (.CI(n31176), .I0(GND_net), .I1(\count[0] [2]), 
            .CO(n31177));
    SB_LUT4 count_0__1148_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [1]), 
            .I3(n31175), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1148_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1148_add_4_3 (.CI(n31175), .I0(GND_net), .I1(\count[0] [1]), 
            .CO(n31176));
    SB_LUT4 count_0__1148_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1148_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1148_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\count[0] [0]), 
            .CO(n31175));
    SB_LUT4 add_1996_24_lut (.I0(GND_net), .I1(n5875[22]), .I2(pwm_setpoint[22]), 
            .I3(n30613), .O(half_duty_new_9__N_664[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1996_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1996_23_lut (.I0(GND_net), .I1(n5875[21]), .I2(pwm_setpoint[21]), 
            .I3(n30612), .O(half_duty_new_9__N_664[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1996_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1996_23 (.CI(n30612), .I0(n5875[21]), .I1(pwm_setpoint[21]), 
            .CO(n30613));
    SB_LUT4 add_1996_22_lut (.I0(GND_net), .I1(n5875[20]), .I2(pwm_setpoint[20]), 
            .I3(n30611), .O(half_duty_new_9__N_664[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1996_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1996_22 (.CI(n30611), .I0(n5875[20]), .I1(pwm_setpoint[20]), 
            .CO(n30612));
    SB_LUT4 add_1996_21_lut (.I0(GND_net), .I1(n5875[19]), .I2(pwm_setpoint[19]), 
            .I3(n30610), .O(half_duty_new_9__N_664[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1996_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1996_21 (.CI(n30610), .I0(n5875[19]), .I1(pwm_setpoint[19]), 
            .CO(n30611));
    SB_LUT4 add_1996_20_lut (.I0(GND_net), .I1(n5875[18]), .I2(pwm_setpoint[18]), 
            .I3(n30609), .O(half_duty_new_9__N_664[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1996_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1996_20 (.CI(n30609), .I0(n5875[18]), .I1(pwm_setpoint[18]), 
            .CO(n30610));
    SB_LUT4 add_1996_19_lut (.I0(GND_net), .I1(n5875[17]), .I2(pwm_setpoint[17]), 
            .I3(n30608), .O(half_duty_new_9__N_664[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1996_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1996_19 (.CI(n30608), .I0(n5875[17]), .I1(pwm_setpoint[17]), 
            .CO(n30609));
    SB_LUT4 add_1996_18_lut (.I0(GND_net), .I1(n5875[16]), .I2(pwm_setpoint[16]), 
            .I3(n30607), .O(half_duty_new_9__N_664[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1996_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1996_18 (.CI(n30607), .I0(n5875[16]), .I1(pwm_setpoint[16]), 
            .CO(n30608));
    SB_LUT4 add_1996_17_lut (.I0(GND_net), .I1(n5875[15]), .I2(pwm_setpoint[15]), 
            .I3(n30606), .O(half_duty_new_9__N_664[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1996_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1996_17 (.CI(n30606), .I0(n5875[15]), .I1(pwm_setpoint[15]), 
            .CO(n30607));
    SB_CARRY add_1996_16 (.CI(n30605), .I0(n5875[14]), .I1(pwm_setpoint[14]), 
            .CO(n30606));
    SB_CARRY add_1996_15 (.CI(n30604), .I0(n5875[13]), .I1(pwm_setpoint[13]), 
            .CO(n30605));
    SB_CARRY add_1996_14 (.CI(n30603), .I0(n5875[12]), .I1(pwm_setpoint[12]), 
            .CO(n30604));
    SB_CARRY add_1996_13 (.CI(n30602), .I0(n5875[11]), .I1(pwm_setpoint[11]), 
            .CO(n30603));
    SB_CARRY add_1996_12 (.CI(n30601), .I0(n5875[10]), .I1(pwm_setpoint[10]), 
            .CO(n30602));
    SB_CARRY add_1996_11 (.CI(n30600), .I0(n5875[9]), .I1(pwm_setpoint[9]), 
            .CO(n30601));
    SB_CARRY add_1996_10 (.CI(n30599), .I0(n5875[8]), .I1(pwm_setpoint[8]), 
            .CO(n30600));
    SB_CARRY add_1996_9 (.CI(n30598), .I0(n5875[7]), .I1(pwm_setpoint[7]), 
            .CO(n30599));
    SB_CARRY add_1996_8 (.CI(n30597), .I0(n5875[6]), .I1(pwm_setpoint[6]), 
            .CO(n30598));
    SB_CARRY add_1996_7 (.CI(n30596), .I0(n5875[5]), .I1(pwm_setpoint[5]), 
            .CO(n30597));
    SB_CARRY add_1996_6 (.CI(n30595), .I0(n5875[4]), .I1(pwm_setpoint[4]), 
            .CO(n30596));
    SB_CARRY add_1996_5 (.CI(n30594), .I0(n5875[3]), .I1(pwm_setpoint[3]), 
            .CO(n30595));
    SB_CARRY add_1996_4 (.CI(n30593), .I0(n5875[2]), .I1(pwm_setpoint[2]), 
            .CO(n30594));
    SB_CARRY add_1996_3 (.CI(n30592), .I0(n5875[1]), .I1(pwm_setpoint[1]), 
            .CO(n30593));
    SB_CARRY add_1996_2 (.CI(GND_net), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[0]), 
            .CO(n30592));
    SB_LUT4 add_2004_23_lut (.I0(GND_net), .I1(pwm_setpoint[21]), .I2(GND_net), 
            .I3(n30591), .O(n5875[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2004_22_lut (.I0(GND_net), .I1(pwm_setpoint[20]), .I2(GND_net), 
            .I3(n30590), .O(n5875[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_22 (.CI(n30590), .I0(pwm_setpoint[20]), .I1(GND_net), 
            .CO(n30591));
    SB_LUT4 add_2004_21_lut (.I0(GND_net), .I1(pwm_setpoint[19]), .I2(GND_net), 
            .I3(n30589), .O(n5875[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_21 (.CI(n30589), .I0(pwm_setpoint[19]), .I1(GND_net), 
            .CO(n30590));
    SB_LUT4 add_2004_20_lut (.I0(GND_net), .I1(pwm_setpoint[18]), .I2(pwm_setpoint[22]), 
            .I3(n30588), .O(n5875[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_20 (.CI(n30588), .I0(pwm_setpoint[18]), .I1(pwm_setpoint[22]), 
            .CO(n30589));
    SB_LUT4 add_2004_19_lut (.I0(GND_net), .I1(pwm_setpoint[17]), .I2(pwm_setpoint[21]), 
            .I3(n30587), .O(n5875[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_19 (.CI(n30587), .I0(pwm_setpoint[17]), .I1(pwm_setpoint[21]), 
            .CO(n30588));
    SB_LUT4 add_2004_18_lut (.I0(GND_net), .I1(pwm_setpoint[16]), .I2(pwm_setpoint[20]), 
            .I3(n30586), .O(n5875[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_18 (.CI(n30586), .I0(pwm_setpoint[16]), .I1(pwm_setpoint[20]), 
            .CO(n30587));
    SB_LUT4 add_2004_17_lut (.I0(GND_net), .I1(pwm_setpoint[15]), .I2(pwm_setpoint[19]), 
            .I3(n30585), .O(n5875[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_17 (.CI(n30585), .I0(pwm_setpoint[15]), .I1(pwm_setpoint[19]), 
            .CO(n30586));
    SB_LUT4 add_2004_16_lut (.I0(GND_net), .I1(pwm_setpoint[14]), .I2(pwm_setpoint[18]), 
            .I3(n30584), .O(n5875[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_16 (.CI(n30584), .I0(pwm_setpoint[14]), .I1(pwm_setpoint[18]), 
            .CO(n30585));
    SB_LUT4 add_2004_15_lut (.I0(GND_net), .I1(pwm_setpoint[13]), .I2(pwm_setpoint[17]), 
            .I3(n30583), .O(n5875[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_15 (.CI(n30583), .I0(pwm_setpoint[13]), .I1(pwm_setpoint[17]), 
            .CO(n30584));
    SB_LUT4 add_2004_14_lut (.I0(GND_net), .I1(pwm_setpoint[12]), .I2(pwm_setpoint[16]), 
            .I3(n30582), .O(n5875[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_14 (.CI(n30582), .I0(pwm_setpoint[12]), .I1(pwm_setpoint[16]), 
            .CO(n30583));
    SB_LUT4 add_2004_13_lut (.I0(GND_net), .I1(pwm_setpoint[11]), .I2(pwm_setpoint[15]), 
            .I3(n30581), .O(n5875[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_13 (.CI(n30581), .I0(pwm_setpoint[11]), .I1(pwm_setpoint[15]), 
            .CO(n30582));
    SB_LUT4 add_2004_12_lut (.I0(GND_net), .I1(pwm_setpoint[10]), .I2(pwm_setpoint[14]), 
            .I3(n30580), .O(n5875[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_12 (.CI(n30580), .I0(pwm_setpoint[10]), .I1(pwm_setpoint[14]), 
            .CO(n30581));
    SB_LUT4 add_2004_11_lut (.I0(GND_net), .I1(pwm_setpoint[9]), .I2(pwm_setpoint[13]), 
            .I3(n30579), .O(n5875[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_11 (.CI(n30579), .I0(pwm_setpoint[9]), .I1(pwm_setpoint[13]), 
            .CO(n30580));
    SB_LUT4 add_2004_10_lut (.I0(GND_net), .I1(pwm_setpoint[8]), .I2(pwm_setpoint[12]), 
            .I3(n30578), .O(n5875[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2004_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2004_10 (.CI(n30578), .I0(pwm_setpoint[8]), .I1(pwm_setpoint[12]), 
            .CO(n30579));
    SB_LUT4 half_duty_0__9__I_0_i7_1_lut (.I0(\half_duty[0][6] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[6]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i8_1_lut (.I0(\half_duty[0][7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[7]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_4_lut (.I0(\count[0] [6]), .I1(\count[0] [0]), .I2(\count[0] [10]), 
            .I3(\count[0] [1]), .O(n20_adj_3565));
    defparam i8_4_lut.LUT_INIT = 16'hbfff;
    SB_LUT4 i7_4_lut_adj_843 (.I0(pause_counter_0), .I1(\count[0] [9]), 
            .I2(\count[0] [8]), .I3(\count[0] [7]), .O(n19));
    defparam i7_4_lut_adj_843.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_3_lut_adj_844 (.I0(\count[0] [4]), .I1(n19), .I2(n20_adj_3565), 
            .I3(GND_net), .O(n6_adj_3566));
    defparam i1_3_lut_adj_844.LUT_INIT = 16'h0202;
    SB_LUT4 i4_4_lut_adj_845 (.I0(\count[0] [5]), .I1(\count[0] [2]), .I2(\count[0] [3]), 
            .I3(n6_adj_3566), .O(n1111));
    defparam i4_4_lut_adj_845.LUT_INIT = 16'h8000;
    SB_LUT4 half_duty_0__9__I_0_i1_1_lut (.I0(\half_duty[0][0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[0]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i2_1_lut (.I0(\half_duty[0][1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[1]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i3_1_lut (.I0(\half_duty[0][2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[2]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i4_1_lut (.I0(\half_duty[0][3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[3]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i5_1_lut (.I0(\half_duty[0][4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[4]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i6_1_lut (.I0(\half_duty[0][5] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[5]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i6_1_lut.LUT_INIT = 16'h5555;
    
endmodule
