// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Thu Dec  5 20:29:53 2019
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, PIN_1, PIN_2, PIN_3, PIN_4, 
            PIN_5, PIN_6, PIN_7, PIN_8, PIN_9, PIN_10, PIN_11, 
            PIN_12, PIN_13, PIN_14, PIN_15, PIN_16, PIN_17, PIN_18, 
            PIN_19, PIN_20, PIN_21, PIN_22, PIN_23, PIN_24) /* synthesis syn_preserve=0, syn_noprune=0, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input PIN_1 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(6[9:14])
    input PIN_2 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(7[9:14])
    inout PIN_3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(8[9:14])
    inout PIN_4 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(9[9:14])
    inout PIN_5 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input PIN_6 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input PIN_7 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    output PIN_8 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(13[9:14])
    input PIN_9 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(14[9:14])
    input PIN_10 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(15[9:15])
    output PIN_11 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(16[9:15])
    inout PIN_12 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(17[9:15])
    input PIN_13 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(18[9:15])
    input PIN_14 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(19[9:15])
    input PIN_15 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(20[9:15])
    input PIN_16 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(21[9:15])
    input PIN_17 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(22[9:15])
    input PIN_18 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(23[9:15])
    output PIN_19 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(24[9:15])
    output PIN_20 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(25[9:15])
    output PIN_21 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(26[9:15])
    output PIN_22 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(27[9:15])
    output PIN_23 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(28[9:15])
    output PIN_24 /* synthesis .original_dir=IN_OUT */ ;   // verilog/TinyFPGA_B.v(29[9:15])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire LED_c /* synthesis SET_AS_NETWORK=LED_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(4[10:13])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire GND_net, VCC_net, PIN_1_c_1, PIN_2_c_0, PIN_6_c_1, PIN_7_c_0, 
        PIN_8_c, PIN_11_c, PIN_13_c, PIN_19_c_0, PIN_20_c, PIN_21_c, 
        PIN_22_c, PIN_23_c;
    wire [31:0]communication_counter;   // verilog/TinyFPGA_B.v(45[9:30])
    wire [23:0]color;   // verilog/TinyFPGA_B.v(46[12:17])
    
    wire blink, hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(129[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(130[21:25])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position;   // verilog/TinyFPGA_B.v(167[22:39])
    wire [23:0]encoder1_position;   // verilog/TinyFPGA_B.v(168[22:39])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(169[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(170[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(171[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(172[22:24])
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(174[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(175[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(176[22:35])
    
    wire n4483;
    wire [23:0]gearBoxRatio;   // verilog/TinyFPGA_B.v(178[22:34])
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(207[22:33])
    
    wire n24190, n6050, n6049, n6048, n6047, n6046, n6045, n6044, 
        n6043, n6042, n6003;
    wire [7:0]color_23__N_164;
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    
    wire n1170, n29889, n1164, n15864, n29888, n4, n28322, n29887, 
        n1481, n29886, n28321, n10, n29885, blink_N_255, n20, 
        n18, n16;
    wire [22:0]pwm_setpoint_22__N_57;
    
    wire PIN_13_N_105, n29884, n41122, n41078, n28137, n28320;
    wire [31:0]motor_state_23__N_106;
    wire [24:0]displacement_23__N_229;
    wire [23:0]displacement_23__N_80;
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire start, \neo_pixel_transmitter.done ;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n28319, n29883, n29882, n29881, n28318, n29880, n28317, 
        n28136;
    wire [3:0]state_3__N_362;
    
    wire n36071, n29879, n28135, n28316;
    wire [31:0]one_wire_N_513;
    
    wire n29878, n28134, n28315, n28314, n28313, n29877, n28312, 
        n29876, n29875, n28133, n28311, n28310, n29874, n6005, 
        n28309, n29873, n29872, n29871, n28308, n75, n28307, n29870, 
        n28306, n28305, n29869, n63, n3006, n28304, n3005, n3004, 
        n29868, n29867, n29866, n29865, n15983, n6070, n6103, 
        n6102, n6099, n6098, n6097, n28303, n1258, n2945_adj_4654, 
        n2947_adj_4655, n2943_adj_4656, n2941, n2939, n2937, n2935, 
        n3133, n3003, n3002, n58, n6096, n70, n6095, n17458, 
        n56, n55, n64, n3001, n1184, n3000, n1318, n1319, n1320, 
        n248, n249, n29864, n2999, n2998, n2997, n65, n2996, 
        n2995, n2994, n2993, n2966, n62, n29863, n4593, n6094, 
        n6091, n6090, n6088, n6119, n6118, n6117, n6116, n6115, 
        n6110, n6109, n6108, n6107, n63_adj_4657, n29862, n60, 
        n28302, n2965, n2964, n2963, n2962, n2961, n2960, n2959, 
        n2958, n2957, n2956, n2955, n2954, n2953, n2952, n2951, 
        n2950, n2949, n2948, n2947, n2946, n2945, n2944, n2943, 
        n28301, n28300, n28299, n939, n938, n919, n918, n917, 
        n916, n915, n914, n1158, n1157, n1156, n1155, n1154, 
        n1153, n1152, n1151, n1553, n1552, n1551, n1550, n41772, 
        n33631;
    wire [9:0]half_duty_new;   // vhdl/pwm.vhd(53[12:25])
    wire [9:0]\half_duty[0] ;   // vhdl/pwm.vhd(55[11:20])
    
    wire n28122, n15980, n28298, n61, n15, n59, n1549, n1548, 
        n1547, n3, n4_adj_4658, n5, n6, n7, n8, n9, n10_adj_4659, 
        n11, n12, n13, n14, n15_adj_4660, n16_adj_4661, n17, n18_adj_4662, 
        n19, n20_adj_4663, n21, n22, n23, n24, n25, n11_adj_4664, 
        rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(90[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(94[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(94[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(94[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(94[12:19])
    
    wire n42067, n28297;
    wire [7:0]\data_in_frame[24] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[22] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(95[12:25])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(96[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(96[12:26])
    
    wire n28121, n15977, n41076;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(101[12:33])
    
    wire tx_active;
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(111[11:16])
    
    wire n28120, n1125, n1124, n1123, n6012, n1122, n1121, n122, 
        n1120;
    wire [31:0]\FRAME_MATCHER.state_31__N_2661 ;
    
    wire n28119, n28118, n28117, n28296, n28116, n28115, n28295, 
        n41766, n28294, n28293, n28292, n41764, n28114, n28113, 
        n28112, n28291, n28111, n28290, n28289, n28288, n28287, 
        n53, n54, n369, n15_adj_4665, n28286, n6004, n28110, n28109, 
        n28285, n28284, n28108, n28107, n28106, n28105, n28104, 
        n28103, n28102, n788, n42075, n28283, n28282, n28281, 
        n28280, n28279, n28278, n35996, n28277, n28101, n28276, 
        n28275, n28274, n28273, n28272, n41752, n28271, n21_adj_4666, 
        n72, n28270, n41750, n41748, n28269, n15974, n28268, n15971, 
        n15966, n15996, n28, n41883, n27, n26, n34343, n25_adj_4667, 
        n32167, n2, n15942, n6_adj_4668, n15910, n27919, n15904, 
        n27918, n27917, n27916, n8_adj_4669, n15901, n27915, n41740, 
        n37483, n35983, n15897, n15893, n16086, n6_adj_4670, n41738, 
        n19670, n29, n41734, n2957_adj_4671, n41732, n3894, n15883, 
        n41722, n41718, n15880, n42338, n15877, n42317, n41709, 
        n15851, n42342, n24984, n4_adj_4672, n2774, n6001, n4698, 
        n15_adj_4673, n4720, n29063, n29062, n29061, n29060, n29059, 
        n29058, n29057, n29056, n29055, n29054, n29053, n29052, 
        n29051, n17934, n17933, n17932, n17931, n17930, n17929, 
        n17928, n17927, n17926, n17925, n17924, n17923, n17922, 
        n17921, n17920, n17919, n17918, n17917, n17916, n17915, 
        n17914, n17913, n17912, n17911, n17910, n17909, n17908, 
        n17907, n17906, n17905, n17904, n17903, n17902, n17901, 
        n17900, n17899, n17898, n17897, n17896, n17895, n17894, 
        n17893, n17892, n17891, n17890, n17889, n17888, n17887, 
        n17886, n17885, n17884, n17883, n17882, n17881, n17880, 
        n17879, n17878, n17877, n17876, n17875, n17874, n17873, 
        n17872, n17871, n17870, n17869, n17868, n17867, n17866, 
        n17865, n17864, n17863, n17862, n17861, n17860, n17859, 
        n17858, n17857, n17856, n17855, n17854, n17853, n17852, 
        n17851, n17850, n17849, n17848, n17847, n17846, n17845, 
        n17844, n17843, n17842, n17841, n17840, n17839, n17838, 
        n17837, n17836, n17835, n17834, n17833, n17832, n17831, 
        n17830, n17829, n17828, n17827, n17826, n17825, n17824, 
        n17823, n17822, n17821, n17820, n17819, n17818, n17817, 
        n17816, n17815, n17814, n17813, n17812, n17811, n17810, 
        n17809, n17808, n17807, n17806, n17805, n17804, n17803, 
        n17802, n17801, n17800, n17799, n17798, n17797, n17796, 
        n17795, n17794, n17793, n17792, n17791, n17790, n17789, 
        n17788, n17787, n17786, n17785, n17784, n17783, n17782, 
        n17781, n17780, n17779, n17778, n17777, n17776, n17775, 
        n17774, n17773, n17772, n17771, n17770, n17769, n17768, 
        n17767, n17766, n17765, n17764, n17763, n17762, n17761, 
        n17760, n17759, n17758, n17757, n17756, n17755, n17754, 
        n17753, n17752, n17751, n17750, n17749, n17748, n17747, 
        n17746, n17745, n17744, n17743, n17742, n17741, n17740, 
        n17739, n17738, n17737, n17736, n17735, n17734, n17733, 
        n17732, n17731, n17730, n17729, n17728, n17727, n17726, 
        n17725, n17724, n17723, n17722, n17721, n17720, n17719, 
        n17718, n6011, n6010, n6009, n42336, n807, n806, n1418, 
        n1419, n786, n785, n784, n783, n1525, n1524, n1523, 
        n1522, n1521, n1520, n1519, n1518, n1517, n1516, n1085, 
        n29050, n6029, n6028, n6027, n6026, n6025, n6024, n6023, 
        n6022, n672, n671, n5945, n5947, n5948, n5950, n29049, 
        n17717, n650, n649, n648, n1058, n1057, n1056, n1055, 
        n1054, n1053, n1052, n17716, n17714, n17713, n17712, n17711, 
        n17710, n17709, n17708, n17707, n17706, n17705, n17704, 
        n17703, n17702, n17701, n17700, n17699, n17698, n17697, 
        n17696, n17695, n17694, n17693, n17692, n33619, n29048, 
        n17687, n17686, n17685, n78, n29047, n17684, n41053, n6039, 
        n6038, n6037, n6055, n6000, n66, n29046, n6054, n558, 
        n29045, n29044, n29043, n25734, n25736, n29042, n28227, 
        n28226, n28225, n28224, n28223, n28222, n29041, n29040, 
        n34409, n29_adj_4674, n29039, n29038, n29037, n35975, n35, 
        n29036, n35966, n42101, n29035, n29034, n77, n29033, n29032, 
        n29031, n29030, n29029, n29028, n29027, n29026, n29025, 
        n29024, n17683, n29023, n29022, n29021, n29020, n29019, 
        n29018, n29017, n15957, n29016, n29015, n29014, n29013, 
        n29012, n29011, n17682, n29010, n42325, n29009, n29008, 
        n74, n29007, n29006, n1283, n29005, n29004, n17681, n29003, 
        n29002, n29001, n29000, n28999, n28998, n28997, n28996, 
        n28995, n28994, n28993, n28992, n28991, n28990, n28989, 
        n28988, n6217, n5_adj_4675, n4451, n28987, n28986, n28985, 
        n28984, n28983, n28982, n4409, n28981, n28980, n28979, 
        n28978, n28977, n4408, n4407, n4406, n4405, n4404, n4403, 
        n4402, n4401, n4400, n4399, n4398, n4397, n4396, n4395, 
        n28976, n28975, n28974, n28973, n28972, n28971, n28970, 
        n28969, n28968, n28967, n28966, n28965, n28964, n28963, 
        n28962, n28961, n28960, n28959, n42335, n17680, n17679, 
        n17678, n17677, n17676, n17675, n17674, n17673, n17672, 
        n17671, n17670, n17669, n17668, n17667, n1025, quadA_debounced, 
        quadB_debounced, count_enable, n1024, n17666, n1257, n1450, 
        n1448, n1449, n10_adj_4676, n25779, n28958, n4394, n4393, 
        n4392, n4391, n4390, n4389, n4388, n4387, n4386, n1256, 
        n9_adj_4677, n1023, n534, n533, n1382, n1022, n1021, quadA_debounced_adj_4678, 
        quadB_debounced_adj_4679, count_enable_adj_4680, n28957, n28956, 
        n17665, n17664, n28955, n17663, n28954, n28953, n28952, 
        n8_adj_4681, n57, n7_adj_4682, n3016, n3015, n3014, n3013, 
        n3012, n3011, n3010, n3009, n3008, n3007, n511, n510, 
        n28951, n6_adj_4683, n17376, n1453, n1454, n1451, n1452, 
        n1456, n17662, n1457, n1455, n28950, n1458, n28949, r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n28948, n17661, n17660, n17659, n17658, n17657, n17656, 
        n33621, n28947, n33623, n28946, n28945, n5999, n5998, 
        n5997, n5996, n5995, n6015, n6014, n28944, n28943, n17637, 
        n28942, n28941, n28940, n41018, n28939, n28938;
    wire [2:0]r_SM_Main_adj_5400;   // verilog/uart_tx.v(31[16:25])
    wire [8:0]r_Clock_Count_adj_5401;   // verilog/uart_tx.v(32[16:29])
    wire [2:0]r_Bit_Index_adj_5402;   // verilog/uart_tx.v(33[16:27])
    
    wire n313, n314, n315, n3_adj_4689, n17625, n17623, n17622, 
        n17621, n17620, n17619, n17618, n17617, n28937, n17616, 
        n33633, n28936, n28935, n28934, n28933, n28932, n28931, 
        n28930, n33635, n17608, n17607, n17606, n316, n317, n318, 
        n319, n320, n28929, n28928, n28927, n28926, n28925, n28924;
    wire [1:0]reg_B;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n17605, n33641, n28923, n28922, n28921;
    wire [1:0]reg_B_adj_5411;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[19:24])
    
    wire n17598, n17597, n17596, n17594, n28920, n28919, n28918, 
        n28917, n28916, n28915, n28914, n28913, n17593, n17591, 
        n17590, n28912, n15960, n28911, n28910, n28909, n17589, 
        n28908, n28907, n28906, n17588, n17587, n33647, n28905, 
        n5_adj_4692, n28904, n28903, n4_adj_4693, n3_adj_4694, n28902, 
        n28901, n28900, n28899, n28898, n28897, n28896, n33649, 
        n28895, n9_adj_4695, n28894, n28893, n8_adj_4696, n28892, 
        n28891, n28890, n28889, n33651, n33653, n13_adj_4697, n28888, 
        n28887, n12_adj_4698, n28886, n28885, n28884, n28883, n28882, 
        n28881, n33655, n20_adj_4699, n19_adj_4700, n18_adj_4701, 
        n28880, n28879, n17_adj_4702, n16_adj_4703, n1255, n15994, 
        n28878, n35676, n33657, n68, n28877, n28876, n28875, n28874, 
        n28873, n16000, n28872, n28871, n28870, n33659, n28869, 
        n28868, n28867, n33661, n28866, n1321, n28865, n28864, 
        n4_adj_4704, n33663, n71, n28863, n28862, n97, n28861, 
        n28860, n28859, n28858, n28857, n1325, n28856, n1324, 
        n13302, n28855, n28854, n1323, n28853, n28852, n33665, 
        n33667, n1354, n1353, n1352, n28851, n1351, n1350, n15874, 
        n28850, n28849, n82, n42878, n28848, n28847, n28846, n81, 
        n80, n79, n28845, n1358, n1357, n1356, n1355, n28844, 
        n28843, n28842, n33669, n33671, n96, n95, n94, n93, 
        n92, n91, n90, n89, n88, n87, n86, n85, n84, n1322, 
        n986, n28841, n28840, n28839, n28838, n28837, n28836, 
        n28835, n28834, n393, n28833, n99, n28832, n28831, n6219, 
        n6218, n28830, n1417, n33673, n28829, n392, n1254, n28828, 
        n28827, n33675, n67, n1349, n6127, n28826, n6112, n28825, 
        n28824, n28823, n28822, n1554, n958, n957, n956, n955, 
        n954, n6101, n6100, n6093, n6092, n6089, n6120, n6114, 
        n953, n28821, n28820, n17541, n73, n17540, n28819, n28818, 
        n7_adj_4705, n6_adj_4706, n28817, n28816, n69, n1253, n1252, 
        n1251, n83, n11_adj_4707, n10_adj_4708, n28815, n28814, 
        n6111, n17537, n1250, n15_adj_4709, n14_adj_4710, n42, n41, 
        n40, n8950, n39, n98, n25_adj_4711, n24_adj_4712, n23_adj_4713, 
        n22_adj_4714, n28813, n28812, n34421, n224, n6113, n28811, 
        n28810, n28809, n28808, n28807, n37, n42333, n28806, n28805, 
        n36, n28804, n1425, n28803, n28802, n1424, n1423, n4_adj_4715, 
        n28801, n28800, n28799, n28798, n28797, n28796, n28795, 
        n28794, n28793, n12_adj_4716, n13_adj_4717, n14_adj_4718, 
        n15_adj_4719, n16_adj_4720, n17_adj_4721, n18_adj_4722, n19_adj_4723, 
        n20_adj_4724, n21_adj_4725, n22_adj_4726, n23_adj_4727, n24_adj_4728, 
        n25_adj_4729, n28792, n28791, n29_adj_4730, n884, n42561, 
        n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
        n1051, n1052_adj_4731, n1053_adj_4732, n1054_adj_4733, n1055_adj_4734, 
        n1056_adj_4735, n1057_adj_4736, n1058_adj_4737, n1059, n1060, 
        n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, 
        n5964, n5965, n5966, n5967, n5968, n5969, n855, n852, 
        n1169, n1170_adj_4738, n1171, n1172, n1173, n1174, n1175, 
        n44342, n1193, n1194, n36026, n34978, n1292, n1293, n1294, 
        n1295, n1296, n1297, n1298, n1299, n1316, n1317, n5983, 
        n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, 
        n28790, n1412, n1413, n1414, n1415, n1416, n1417_adj_4739, 
        n1418_adj_4740, n1419_adj_4741, n1420, n18307, n41613, n28789, 
        n28788, n1436, n1437, n28787, n28786, n28785, n28784, 
        n28783, n28782, n28781, n28780, n36012, n28779, n28778, 
        n35969, n28777, n28776, n28775, n749, n748, n746, n1529, 
        n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, 
        n1538, n1553_adj_4742, n1554_adj_4743, n28774, n36058, n28773, 
        n28772, n28771, n28770, n42328, n6016, n6017, n6018, n6019, 
        n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, 
        n1651, n1652, n1653, n1667, n1668, n28769, n35948, n28768, 
        n28767, n28766, n28765, n28764, n28763, n6030, n6031, 
        n6032, n6033, n6034, n28762, n28761, n18259, n18258, n1754, 
        n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, 
        n1763, n1764, n1765, n18256, n18255, n18254, n18253, n18252, 
        n18251, n1778, n1779, n18250, n18249, n18248, n18247, 
        n18246, n18245, n18244, n18243, n18242, n18241, n18240, 
        n18239, n1862, n1863, n1864, n1865, n1866, n1867, n1868, 
        n1869, n1870, n1871, n1872, n1873, n1874, n1886, n1887, 
        n18238, n18237, n18236, n18235, n18234, n18233, n18232, 
        n18231, n18230, n18229, n6056, n6057, n6058, n6059, n6060, 
        n6061, n6062, n6063, n6064, n6065, n6066, n6067, n35936, 
        n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, 
        n1975, n1976, n1977, n1978, n1979, n1980, n18223, n41571, 
        n18222, n1991, n1992, n28760, n18215, n6071, n6072, n6073, 
        n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, 
        n6082, n6083, n6084, n6085, n18213, n18212, n2069, n2070, 
        n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, 
        n2079, n2080, n2081, n2082, n2083, n2093, n2094, n28759, 
        n28758, n43572, n43575, n43578, n43581, n18203, n6104, 
        n3452, n3453, n3454, n3455, n3456, n3458, n18202, n18201, 
        n18200, n18199, n2168, n2169, n2170, n2171, n2172, n2173, 
        n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, 
        n2182, n2183, n18198, n18197, n18196, n18195, n2192, n2193, 
        n18194, n18193, n18192, n18191, n18190, n18189, n18188, 
        n18187, n18186, n18185, n6121, n6122, n6123, n6124, n6167, 
        n6190, n16003, n6214, n18184, n18183, n18182, n2264, n2265, 
        n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, 
        n2274, n2275, n2276, n2277, n2278, n2279, n2280, n18181, 
        n18179, n18178, n2288, n2289, n18177, n18176, n18175, 
        n40975, n18174, n18173, n40971, n6128, n6129, n6130, n6131, 
        n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, 
        n6140, n6141, n6142, n6143, n6144, n6145, n18172, n18171, 
        n18170, n2357, n2358, n2359, n2360, n2361, n2362, n2363, 
        n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, 
        n2372, n2373, n2374, n18169, n18168, n18167, n2381, n2382, 
        n18166, n18165, n18164, n18163, n18162, n6148, n6149, 
        n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, 
        n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, 
        n6166, n18161, n2447, n2448, n2449, n2450, n2451, n2452, 
        n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, 
        n2461, n2462, n2463, n2464, n2465, n18160, n18159, n2471, 
        n2472, n18158, n18157, n28757, n12_adj_4744, n6170, n6171, 
        n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, 
        n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, 
        n6188, n6189, n18156, n18155, n18154, n2534, n2535, n2536, 
        n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, 
        n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, 
        n2553, n42341, n2558, n2559, n18153, n18152, n28756, n28755, 
        n28754, n28753, n28752, n28751, n28750, n18151, n6193, 
        n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, 
        n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, 
        n6210, n6211, n6212, n6213, n2618, n2619, n2620, n2621, 
        n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, 
        n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, 
        n2638, n2642, n2643, n18150, n6220, n6221, n6222, n6223, 
        n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, 
        n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, 
        n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, 
        n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, 
        n2715, n2716, n2717, n2718, n2719, n2720, n3362, n2723, 
        n2724, n17011, n28749, n3360, n2777, n2798, n2799, n28213, 
        n2801, n2802, n41555, n42099, n28212, n18149, n18148, 
        n18147, n18146, n18145, n18144, n18143, n18142, n18141, 
        n18140, n18139, n18138, n18137, n42326, n3357, n3356, 
        n3355, n3354, n3353, n3351, n3346, n3344, n3343, n3340, 
        n3337, n18136, n18135, n18134, n28748, n28747, n28746, 
        n3330, n28745, n28744, n18133, n28743, n18132, n18131, 
        n3325, n3324, n28742, n28741, n3323, n3322, n28740, n3321, 
        n3320, n3319, n18130, n18129, n18128, n18127, n18126, 
        n3318, n3317, n3316, n3315, n3314, n3313, n3312, n3311, 
        n28739, n3310, n3309, n3308, n3307, n3306, n28738, n3305, 
        n42725, n3304, n3303, n3302, n3301, n3300, n28737, n3299, 
        n28736, n3298, n28735, n28734, n28733, n28732, n28731, 
        n28730, n28729, n17513, n17256, n17250, n18021, n18020, 
        n17510, n63_adj_4745, n1422, n41561, n3263, n28728, n17203, 
        n3258, n3257, n3256, n3255, n3254, n3253, n3252, n3251, 
        n3250, n3249, n3248, n3247, n3246, n17506, n3245, n17385, 
        n3244, n3243, n3242, n3241, n3240, n3239, n3238, n3237, 
        n3236, n3235, n3234, n3233, n3232, n3231, n17505, n3230, 
        n18019, n3225, n3224, n1421, n3223, n18018, n3222, n3221, 
        n3220, n3219, n3218, n3217, n3216, n3215, n3214, n3213, 
        n3212, n17503, n3211, n3210, n3209, n3208, n3207, n3206, 
        n3205, n3204, n3203, n3202, n3201, n3200, n3199, n28727, 
        n28726, n6002, n3164, n28725, n3158, n3157, n3156, n3155, 
        n3154, n3153, n3152, n3151, n3150, n3149, n3148, n3147, 
        n3146, n3145, n3144, n3143, n3142, n3141, n3140, n3139, 
        n3138, n3137, n3136, n3135, n41551, n28724, n28723, n28722, 
        n42434, n28721, n40963, n42603, n28720, n40957, n42851, 
        n28719, n3134, n6_adj_4746, n42115, n28718, n42147, n3132, 
        n3131, n3125, n3124, n42876, n3123, n3122, n3121, n42872, 
        n3120, n3119, n3118, n3117, n3116, n3115, n3114, n3113, 
        n3112, n3111, n3110, n3109, n3108, n3107, n3106, n3105, 
        n3104, n3103, n3102, n3101, n3100, n3065, n28717, n3058, 
        n3057, n3056, n3055, n3054, n28716, n3053, n3052, n28715, 
        n28714, n3051, n28713, n28712, n3050, n3049, n3048, n28711, 
        n3047, n3046, n28710, n28709, n3045, n28708, n3044, n3043, 
        n3042, n3041, n3040, n3039, n3038, n3037, n3036, n3035, 
        n3034, n3033, n3032, n42868, n3025, n3024, n3023, n3022, 
        n3021, n3020, n3019, n3018, n3017, n3016_adj_4747, n3015_adj_4748, 
        n3014_adj_4749, n3013_adj_4750, n3012_adj_4751, n3011_adj_4752, 
        n3010_adj_4753, n3009_adj_4754, n3008_adj_4755, n3007_adj_4756, 
        n3006_adj_4757, n3005_adj_4758, n3004_adj_4759, n3003_adj_4760, 
        n3002_adj_4761, n3001_adj_4762, n2966_adj_4763, n28707, n2958_adj_4764, 
        n2957_adj_4765, n5_adj_4766, n2956_adj_4767, n2955_adj_4768, 
        n2954_adj_4769, n2953_adj_4770, n2952_adj_4771, n2951_adj_4772, 
        n2950_adj_4773, n2949_adj_4774, n28706, n2948_adj_4775, n28705, 
        n2946_adj_4776, n28704, n2944_adj_4777, n28703, n2942, n28702, 
        n2940, n28701, n2938, n28700, n2936, n6013, n2934, n2933, 
        n42867, n2925, n2924, n2923, n2922, n2921, n2920, n2919, 
        n2918, n2917, n2916, n2915, n2914, n2913, n2912, n2911, 
        n2910, n2909, n2908, n2907, n2906, n2905, n2904, n2903, 
        n2902, n28699, n40949, n42_adj_4778, n42117, n33, n32, 
        n31, n30, n35991, n36038, n1912, n1913, n1914, n1915, 
        n1916, n1917, n1918, n1919, n1920, n1921, n1953, n1922, 
        n1954, n1923, n1955, n1924, n1956, n1925, n1957, n1958, 
        n1943, n28698, n1944, n1976_adj_4779, n1945, n1946, n1947, 
        n1948, n33629, n1949, n1950, n1951, n1952, n3358, n134, 
        n135, n136, n137, n138, n139, n140, n141, n142, n143, 
        n144, n145, n146, n147, n148, n149, n150, n151, n152, 
        n153, n154, n155, n156, n157, n158, n159, n160, n161, 
        n162, n163, n164, n165, n28697, n1877, n36089, n1844, 
        n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, 
        n1853, n1854, n1855, n1856, n1857, n1858, n29_adj_4780, 
        n28_adj_4781, n27_adj_4782, n26_adj_4783, n25_adj_4784, n24_adj_4785, 
        n23_adj_4786, n22_adj_4787, n21_adj_4788, n20_adj_4789, n19_adj_4790, 
        n18_adj_4791, n17_adj_4792, n16_adj_4793, n15_adj_4794, n14_adj_4795, 
        n13_adj_4796, n12_adj_4797, n11_adj_4798, n10_adj_4799, n9_adj_4800, 
        n8_adj_4801, n7_adj_4802, n6_adj_4803, n5_adj_4804, n4_adj_4805, 
        n3_adj_4806, n28696, n2858, n2857, n2856, n2855, n2854, 
        n2853, n2852, n2851, n2850, n2849, n2848, n2847, n2846, 
        n42854, n2845, n2844, n2843, n2842, n2841, n2840, n2839, 
        n2838, n2837, n2836, n1745, n1746, n1747, n1748, n1749, 
        n1750, n1751, n1752, n1753, n1754_adj_4807, n1755_adj_4808, 
        n1756_adj_4809, n1757_adj_4810, n1758_adj_4811, n42141, n42852, 
        n28695, n1778_adj_4812, n33617, n1813, n1814, n1815, n1816, 
        n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, 
        n1825, n2867, n2834, n2835, n1714, n1715, n1716, n1717, 
        n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, 
        n28694, n1679, n1646_adj_4813, n1647_adj_4814, n1648_adj_4815, 
        n1649_adj_4816, n1650_adj_4817, n1651_adj_4818, n1652_adj_4819, 
        n1653_adj_4820, n1654, n1655, n1656, n1657, n1658, n33643, 
        n33645, n17445, n17444, n17500, n17497, n17494, n17491, 
        n5946, n42846, n1615, n1616, n1617, n2824, n1618, n1619, 
        n1620, n1621, n1622, n1623, n1225, n1624, n1224, n1625, 
        n1223, n1222, n1221, n1220, n1219, n2825, n28693, n1580, 
        n2823, n17488, n17485, n2819, n2822, n2820, n2821, n2818, 
        n1557, n1558, n2814, n28211, n2817, n2815, n2816, n1555, 
        n1556, n2813, n2812, n2811, n2810, n2809, n2808, n2807, 
        n2806, n2805, n2804, n2803, n28692, n40_adj_4821, n42_adj_4822, 
        n44, n45, n42135, n2768, n28691, n42840, n28690, n2758, 
        n2757, n2756, n2755, n2754, n2753, n2752, n2751, n2750, 
        n2749, n2748, n2747, n2746, n2745, n2744, n2743, n2742, 
        n2741, n2740, n2739, n2738, n2737, n2736, n2735, n42875, 
        n2725, n2724_adj_4823, n2723_adj_4824, n2722, n2721, n2720_adj_4825, 
        n2719_adj_4826, n2718_adj_4827, n2717_adj_4828, n2716_adj_4829, 
        n2715_adj_4830, n2714_adj_4831, n28689, n2713_adj_4832, n2712_adj_4833, 
        n2711_adj_4834, n2710_adj_4835, n2709_adj_4836, n2708_adj_4837, 
        n2707_adj_4838, n2706_adj_4839, n2705_adj_4840, n2704_adj_4841, 
        n6041, n2669, n28688, n2658, n2657, n2656, n2655, n2654, 
        n2653, n2652, n2651, n28687, n44_adj_4842, n2650, n2649, 
        n2648, n2647, n2646, n2645, n2644, n2643_adj_4843, n2642_adj_4844, 
        n2641, n2640, n2639, n2638_adj_4845, n2637_adj_4846, n2636_adj_4847, 
        n6040, n2625_adj_4848, n2624_adj_4849, n2623_adj_4850, n2622_adj_4851, 
        n2621_adj_4852, n2620_adj_4853, n2619_adj_4854, n2618_adj_4855, 
        n2617, n2616, n2615, n2614, n2613, n2612, n2611, n2610, 
        n2609, n2608, n2607, n2606, n2605, n28686, n46, n42871, 
        n2570, n28685, n28684, n28683, n2558_adj_4856, n2557, n2556, 
        n2555, n2554, n2553_adj_4857, n2552_adj_4858, n2551_adj_4859, 
        n2550_adj_4860, n2549_adj_4861, n2548_adj_4862, n2547_adj_4863, 
        n2546_adj_4864, n2545_adj_4865, n2544_adj_4866, n2543_adj_4867, 
        n2542_adj_4868, n2541_adj_4869, n2540_adj_4870, n2539_adj_4871, 
        n2538_adj_4872, n2537_adj_4873, n2525, n28682, n40928, n2524, 
        n2523, n2522, n2521, n2520, n2519, n2518, n2517, n2516, 
        n2515, n2514, n2513, n28681, n2512, n28680, n2511, n28679, 
        n2510, n2509, n2508, n2507, n2506, n2471_adj_4874, n28678, 
        n2458_adj_4875, n2457_adj_4876, n2456_adj_4877, n2455_adj_4878, 
        n2454_adj_4879, n1420_adj_4880, n2453_adj_4881, n2452_adj_4882, 
        n2451_adj_4883, n2450_adj_4884, n2449_adj_4885, n2448_adj_4886, 
        n2447_adj_4887, n2446, n2445, n2444, n2443, n2442, n2441, 
        n2440, n2439, n2438, n41601, n2_adj_4888, n3_adj_4889, n4_adj_4890, 
        n5_adj_4891, n6_adj_4892, n7_adj_4893, n8_adj_4894, n9_adj_4895, 
        n10_adj_4896, n11_adj_4897, n12_adj_4898, n13_adj_4899, n14_adj_4900, 
        n15_adj_4901, n16_adj_4902, n17_adj_4903, n18_adj_4904, n19_adj_4905, 
        n20_adj_4906, n21_adj_4907, n22_adj_4908, n23_adj_4909, n24_adj_4910, 
        n25_adj_4911, n2_adj_4912, n3_adj_4913, n4_adj_4914, n5_adj_4915, 
        n6_adj_4916, n7_adj_4917, n8_adj_4918, n9_adj_4919, n10_adj_4920, 
        n11_adj_4921, n12_adj_4922, n13_adj_4923, n14_adj_4924, n15_adj_4925, 
        n16_adj_4926, n17_adj_4927, n18_adj_4928, n19_adj_4929, n20_adj_4930, 
        n21_adj_4931, n22_adj_4932, n23_adj_4933, n24_adj_4934, n25_adj_4935, 
        n2425, n2424, n2423, n2422, n2421, n2420, n2419, n2418, 
        n2417, n2416, n2415, n2414, n2413, n2412, n2411, n2410, 
        n2409, n2408, n2407, n28677, n38, n40_adj_4936, n42_adj_4937, 
        n43, n13_adj_4938, n2372_adj_4939, n28676, n2358_adj_4940, 
        n2357_adj_4941, n2356, n2355, n2354, n2353, n2352, n2351, 
        n2350, n2349, n28675, n36_adj_4942, n38_adj_4943, n40_adj_4944, 
        n41_adj_4945, n42623, n2348, n2347, n2346, n2345, n2344, 
        n2343, n2342, n2341, n2340, n2339, n2325, n2324, n2323, 
        n2322, n2321, n2320, n2319, n2318, n2317, n2316, n2315, 
        n2314, n2313, n2312, n2311, n2310, n2309, n2308, n28674, 
        n34, n36_adj_4946, n38_adj_4947, n39_adj_4948, n41_adj_4949, 
        n43_adj_4950, n44_adj_4951, n45_adj_4952, n42155, n42849, 
        n42807, n41507, n2273_adj_4953, n28673, n28672, n32_adj_4954, 
        n34_adj_4955, n37_adj_4956, n39_adj_4957, n41_adj_4958, n42605, 
        n43_adj_4959, n42157, n2258, n2257, n2256, n2255, n2254, 
        n2253, n2252, n2251, n2250, n2249, n2248, n2247, n2246, 
        n2245, n2244, n2243, n2242, n2241, n2240, n2225, n2224, 
        n2223, n2222, n28671, n30_adj_4960, n31_adj_4961, n32_adj_4962, 
        n33_adj_4963, n34_adj_4964, n35_adj_4965, n37_adj_4966, n39_adj_4967, 
        n41_adj_4968, n42_adj_4969, n43_adj_4970, n45_adj_4971, n42788, 
        n2221, n2220, n2219, n2218, n2217, n2216, n28670, n2215, 
        n2214, n2213, n2212, n2211, n2210, n2209, n41839, n40905, 
        n36533, n28669, n40901, n28_adj_4972, n29_adj_4973, n30_adj_4974, 
        n31_adj_4975, n32_adj_4976, n33_adj_4977, n35_adj_4978, n37_adj_4979, 
        n42597, n39_adj_4980, n40_adj_4981, n41_adj_4982, n43_adj_4983, 
        n42595, n42753, n40899, n2174_adj_4984, n28668, n2158, n2157, 
        n2156, n2155, n2154, n2153, n2152, n28667, n26_adj_4985, 
        n27_adj_4986, n28_adj_4987, n29_adj_4988, n30_adj_4989, n31_adj_4990, 
        n33_adj_4991, n35_adj_4992, n42593, n37_adj_4993, n38_adj_4994, 
        n39_adj_4995, n41_adj_4996, n42415, n42869, n2151, n2150, 
        n2149, n2148, n2147, n2146, n2145, n2144, n2143, n2142, 
        n2141, n28210, n28666, n28665, n2125, n2124, n2123, n2122, 
        n28664, n40891, n24_adj_4997, n25_adj_4998, n26_adj_4999, 
        n27_adj_5000, n28_adj_5001, n29_adj_5002, n30_adj_5003, n31_adj_5004, 
        n32_adj_5005, n33_adj_5006, n35_adj_5007, n36_adj_5008, n37_adj_5009, 
        n39_adj_5010, n42417, n2121, n2120, n2119, n2118, n2117, 
        n2116, n2115, n2114, n2113, n2112, n2111, n2110, n40889, 
        n40887, n28663, n22_adj_5011, n23_adj_5012, n24_adj_5013, 
        n25_adj_5014, n26_adj_5015, n27_adj_5016, n28_adj_5017, n29_adj_5018, 
        n30_adj_5019, n31_adj_5020, n33_adj_5021, n34_adj_5022, n35_adj_5023, 
        n37_adj_5024, n39_adj_5025, n42570, n41_adj_5026, n43_adj_5027, 
        n42425, n42711, n15963, n41835, n33639, n2075_adj_5028, 
        n28662, n28661, n20_adj_5029, n21_adj_5030, n22_adj_5031, 
        n23_adj_5032, n24_adj_5033, n25_adj_5034, n26_adj_5035, n27_adj_5036, 
        n28_adj_5037, n29_adj_5038, n31_adj_5039, n32_adj_5040, n33_adj_5041, 
        n35_adj_5042, n37_adj_5043, n42558, n39_adj_5044, n41_adj_5045, 
        n42731, n28209, n43569, n28208, n2058, n2057, n2056, n2055, 
        n2054, n2053, n2052, n2051, n2050, n2049, n28660, n18_adj_5046, 
        n19_adj_5047, n20_adj_5048, n21_adj_5049, n22_adj_5050, n23_adj_5051, 
        n24_adj_5052, n25_adj_5053, n26_adj_5054, n27_adj_5055, n29_adj_5056, 
        n30_adj_5057, n31_adj_5058, n33_adj_5059, n35_adj_5060, n42783, 
        n37_adj_5061, n39_adj_5062, n41_adj_5063, n43_adj_5064, n45_adj_5065, 
        n42427, n2048, n2047, n2046, n2045, n2044, n2043, n2042, 
        n28659, n16_adj_5066, n17_adj_5067, n18_adj_5068, n19_adj_5069, 
        n20_adj_5070, n21_adj_5071, n22_adj_5072, n23_adj_5073, n25_adj_5074, 
        n27_adj_5075, n28_adj_5076, n29_adj_5077, n31_adj_5078, n33_adj_5079, 
        n35_adj_5080, n37_adj_5081, n39_adj_5082, n41_adj_5083, n43_adj_5084, 
        n42806, n2025, n2024, n2023, n2022, n2021, n2020, n2019, 
        n2018, n2017, n2016, n28658, n14_adj_5085, n16_adj_5086, 
        n17_adj_5087, n18_adj_5088, n19_adj_5089, n20_adj_5090, n21_adj_5091, 
        n22_adj_5092, n23_adj_5093, n25_adj_5094, n26_adj_5095, n27_adj_5096, 
        n29_adj_5097, n31_adj_5098, n33_adj_5099, n35_adj_5100, n37_adj_5101, 
        n42337, n39_adj_5102, n40_adj_5103, n41_adj_5104, n43_adj_5105, 
        n45_adj_5106, n42755, n2015, n2014, n2013, n2012, n2011, 
        n28657, n12_adj_5107, n14_adj_5108, n15_adj_5109, n16_adj_5110, 
        n17_adj_5111, n18_adj_5112, n19_adj_5113, n20_adj_5114, n21_adj_5115, 
        n23_adj_5116, n24_adj_5117, n25_adj_5118, n27_adj_5119, n29_adj_5120, 
        n31_adj_5121, n42792, n33_adj_5122, n35_adj_5123, n42572, 
        n37_adj_5124, n38_adj_5125, n39_adj_5126, n41_adj_5127, n43_adj_5128, 
        n42726, n40867, n28656, n10_adj_5129, n12_adj_5130, n13_adj_5131, 
        n14_adj_5132, n15_adj_5133, n16_adj_5134, n17_adj_5135, n18_adj_5136, 
        n19_adj_5137, n21_adj_5138, n22_adj_5139, n23_adj_5140, n25_adj_5141, 
        n27_adj_5142, n29_adj_5143, n42794, n31_adj_5144, n33_adj_5145, 
        n42564, n35_adj_5146, n36_adj_5147, n37_adj_5148, n39_adj_5149, 
        n41_adj_5150, n42796, n42881, n28655, n28654, n8_adj_5151, 
        n10_adj_5152, n11_adj_5153, n12_adj_5154, n13_adj_5155, n14_adj_5156, 
        n15_adj_5157, n16_adj_5158, n17_adj_5159, n19_adj_5160, n20_adj_5161, 
        n21_adj_5162, n23_adj_5163, n25_adj_5164, n42560, n27_adj_5165, 
        n29_adj_5166, n31_adj_5167, n42727, n33_adj_5168, n34_adj_5169, 
        n35_adj_5170, n37_adj_5171, n39_adj_5172, n42456, n41_adj_5173, 
        n42777, n43_adj_5174, n44_adj_5175, n45_adj_5176, n42458, 
        n42803, n28653, n6_adj_5177, n8_adj_5178, n9_adj_5179, n10_adj_5180, 
        n11_adj_5181, n12_adj_5182, n13_adj_5183, n14_adj_5184, n15_adj_5185, 
        n17_adj_5186, n19_adj_5187, n21_adj_5188, n23_adj_5189, n24_adj_5190, 
        n25_adj_5191, n27_adj_5192, n29_adj_5193, n31_adj_5194, n32_adj_5195, 
        n33_adj_5196, n35_adj_5197, n37_adj_5198, n42723, n28652, 
        n40856, n4_adj_5199, n6_adj_5200, n7_adj_5201, n8_adj_5202, 
        n9_adj_5203, n10_adj_5204, n11_adj_5205, n12_adj_5206, n13_adj_5207, 
        n15_adj_5208, n16_adj_5209, n17_adj_5210, n19_adj_5211, n21_adj_5212, 
        n42327, n23_adj_5213, n24_adj_5214, n25_adj_5215, n27_adj_5216, 
        n29_adj_5217, n30_adj_5218, n31_adj_5219, n33_adj_5220, n35_adj_5221, 
        n37_adj_5222, n39_adj_5223, n41_adj_5224, n43_adj_5225, n45_adj_5226, 
        n42761, n18017, n28207, n28651, n5973, n5974, n5975, n5976, 
        n5977, n5978, n5979, n5980, n5992, n5962, n5963, n18016, 
        n18015, n28206, n28205, n16_adj_5227, n36097, n5954, n5955, 
        n5956, n5957, n5958, n5959, n11_adj_5228, n10_adj_5229, 
        n28650, n10_adj_5230, n42853, n42799, n42797, n28649, n28648, 
        n28647, n28646, n28645, n28644, n42759, n42369, n24_adj_5231, 
        n36043, n22_adj_5232, n20_adj_5233, n12_adj_5234, n28643, 
        n28642, n28641, n28640, n28639, n28638, n28637, n28636, 
        n28635, n16_adj_5235, n28195, n33589, n33601, n33595, n42781, 
        n41479, n41471, n37_adj_5236, n35_adj_5237, n34_adj_5238, 
        n32_adj_5239, n31_adj_5240, n25_adj_5241, n5_adj_5242, n42883, 
        n41452, n41446, n41440, n8_adj_5243, n43830, n42730, n42724, 
        n28_adj_5244, n41436, n42133, n41430, n42722, n42721, n26_adj_5245, 
        n24_adj_5246, n41426, n19_adj_5247, n16_adj_5248, n42716, 
        n36006, n43694, n3209_adj_5249, n28194, n28193, n18014, 
        n13_adj_5250, n11_adj_5251, n40846, n42790, n42708, n42706, 
        n28192, n40842, n28191, n36105, n42679, n28190, n28189, 
        n42662, n42661, n15987, n36053, n36008, n28188, n36556, 
        n42153, n28187, n43565, n36110, n42652, n41390, n4_adj_5252, 
        n41385, n42651, n42559, n42793, n42644, n42643, n10249, 
        n10248, n10247, n10246, n10245, n42636, n10244, n41375, 
        n6_adj_5253, n42634, n40836, n41368, n42618, n42617, n42472, 
        n41363, n11_adj_5254, n42610, n42609, n42606, n42604, n42602, 
        n42601, n42598, n42594, n42557, n38_adj_5255, n37_adj_5256, 
        n42590, n36_adj_5257, n42589, n42791, n41329, n35_adj_5258, 
        n15740, n41326, n41324, n33_adj_5259, n42189, n41321, n42573, 
        n26_adj_5260, n42569, n41314, n42565, n22_adj_5261, n42464, 
        n34_adj_5262, n33_adj_5263, n34989, n32_adj_5264, n42462, 
        n31_adj_5265, n30_adj_5266, n42453, n42451, n42191, n42447, 
        n42553, n41296, n42441, n42430, n36526, n42412, n15889, 
        n42408, n42404, n40828, n42398, n42552, n28570, n28569, 
        n28568, n28567, n28566, n28565, n3_adj_5267, n28564, n28563, 
        n28562, n42484, n28561, n28560, n28559, n28558, n28557, 
        n28556, n41276, n28555, n28554, n28553, n28186, n28185, 
        n41274, n28552, n28551, n28550, n40824, n42884, n28549, 
        n28548, n41272, n42549, n28547, n28546, n28545, n42787, 
        n41270, n41268, n28544, n28543, n28542, n41258, n28541, 
        n28540, n41244, n41242, n28539, n28538, n28184, n28537, 
        n2_adj_5268, n28536, n4_adj_5269, n28535, n28534, n28533, 
        n28532, n41819, n42544, n36076, n28531, n28530, n41238, 
        n28529, n28528, n28527, n24824, n28526, n5949, n41226, 
        n5953, n42541, n41877, n5972, n41222, n6008, n28525, n28524, 
        n6053, n42665, n40820, n42767, n41216, n40818, n40815, 
        n40805, n42882, n41212, n40798, n40794, n40780, n8_adj_5270, 
        n7_adj_5271, n28523, n38429, n4_adj_5272, n38425, n42547, 
        n28522, n28521, n28520, n42786, n28519, n28518, n2_adj_5273, 
        n28517, n28516, n35946, n40747, n40746, n40745, n40744, 
        n40743, n40742, n40740, n28183, n38401, n42536, n28515, 
        n18_adj_5274, n40730, n40728, n42490, n40726, n40725, n40724, 
        n2_adj_5275, n3_adj_5276, n4_adj_5277, n5_adj_5278, n6_adj_5279, 
        n7_adj_5280, n8_adj_5281, n9_adj_5282, n10_adj_5283, n11_adj_5284, 
        n12_adj_5285, n13_adj_5286, n14_adj_5287, n15_adj_5288, n16_adj_5289, 
        n17_adj_5290, n18_adj_5291, n19_adj_5292, n20_adj_5293, n21_adj_5294, 
        n22_adj_5295, n23_adj_5296, n24_adj_5297, n25_adj_5298, n26_adj_5299, 
        n27_adj_5300, n28_adj_5301, n29_adj_5302, n30_adj_5303, n31_adj_5304, 
        n32_adj_5305, n33_adj_5306, n28514, n28513, n28512, n28511, 
        n28510, n40723, n28509, n28508, n28507, n28506, n28505, 
        n28504, n28503, n28502, n28501, n28500, n28499, n28498, 
        n28497, n35940, n28496, n28495, n28494, n28493, n28492, 
        n28182, n47, n40722, n46_adj_5307, n40721, n43_adj_5308, 
        n42_adj_5309, n40_adj_5310, n28491, n28490, n28489, n28488, 
        n39_adj_5311, n28487, n28486, n28181, n38_adj_5312, n28485, 
        n40720, n28484, n28483, n32_adj_5313, n28482, n28481, n28480, 
        n28479, n28478, n28477, n40719, n28476, n40718, n40717, 
        n28475, n28474, n28473, n28472, n40716, n28471, n28470, 
        n40715, n40714, n28469, n28468, n28467, n28180, n28466, 
        n28465, n28464, n28463, n28462, n28461, n28460, n28459, 
        n40713, n22_adj_5314, n40712, n40711, n19_adj_5315, n40710, 
        n18_adj_5316, n28458, n28457, n28456, n28455, n28454, n28453, 
        n15_adj_5317, n40709, n28452, n28451, n28450, n28179, n28449, 
        n28448, n28447, n28446, n28445, n42880, n28444, n40708, 
        n40707, n28443, n28442, n28441, n28440, n28439, n28438, 
        n28437, n35942, n28436, n28435, n28434, n40706, n28433, 
        n28432, n28431, n40772, n24794, n28430, n24918, n32_adj_5318, 
        n40705, n31_adj_5319, n28178, n30_adj_5320, n29_adj_5321, 
        n28_adj_5322, n40704, n42500, n42782, n28429, n28428, n28427, 
        n28426, n40703, n28425, n40702, n40701, n40700, n28424, 
        n40699, n28423, n28422, n28421, n42249, n28420, n28419, 
        n40770, n28418, n28417, n28416, n28415, n28414, n28413, 
        n28412, n28411, n28410, n28177, n28409, n28408, n40698, 
        n28407, n28406, n28405, n28404, n24782, n28403, n28402, 
        n28401, n28400, n28399, n28176, n42681, n28398, n28397, 
        n28396, n42780, n40690, n40689, n28395, n28394, n28393, 
        n28392, n28175, n28391, n28390, n28389, n28388, n28387, 
        n38277, n28386, n28385, n28174, n28384, n28383, n28382, 
        n28381, n23989, n28380, n28379, n28378, n28377, n28376, 
        n28375, n28374, n28373, n28372, n28371, n28370, n28369, 
        n28368, n28367, n28366, n28365, n28364, n28363, n28362, 
        n28361, n28360, n28173, n28172, n28359, n28171, n28170, 
        n28358, n28357, n28356, n28355, n28354, n28169, n2_adj_5323, 
        n28353, n28352, n28351, n28168, n28167, n28166, n28350, 
        n28349, n28348, n28347, n28346, n28345, n28344, n38596, 
        n28343, n28342, n28341, n40674, n41969, n28340, n28339, 
        n28338, n28337, n28336, n41979, n28335, n28334, n28333, 
        n28332, n28331, n28330, n28142, n28329, n28328, n28141, 
        n28140, n28139, n28327, n35873, n28326, n28325, n28324, 
        n35865, n28323, n42779, n28138, n29892, n29891, n29890, 
        n38205, n38575, n35825, n36342, n38562, n42348, n38171, 
        n34167, n40768, n42506, n38513, n38143, n38137, n38133, 
        n35833, n40651, n34225, n38109, n38107, n38105, n38103, 
        n30_adj_5324, n29_adj_5325, n28_adj_5326, n27_adj_5327, n38101, 
        n38099, n18_adj_5328, n34267, n34315, n3_adj_5329, n38059, 
        n38057, n35644, n38051, n38049, n38047, n37132, n35463, 
        n17_adj_5330, n38031, n38027, n47_adj_5331, n16_adj_5332, 
        n36518, n38464, n35626, n35562, n26_adj_5333, n24_adj_5334, 
        n22_adj_5335, n18_adj_5336, n46_adj_5337, n5_adj_5338, n37622, 
        n38584, n34419, n28_adj_5339, n43653, n5_adj_5340, n42347, 
        n13_adj_5341, n40756, n40_adj_5342, n39_adj_5343, n38_adj_5344, 
        n44_adj_5345, n43_adj_5346, n37_adj_5347, n42_adj_5348, n41_adj_5349, 
        n40_adj_5350, n38_adj_5351, n30_adj_5352, n26_adj_5353, n35_adj_5354, 
        n34_adj_5355, n28_adj_5356, n43635, n40620, n40619, n40616, 
        n42775, n41061, n37785, n6_adj_5357, n37783, n16_adj_5358, 
        n42307, n16_adj_5359, n37725;
    
    VCC i2 (.Y(VCC_net));
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[0]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_LUT4 i18_4_lut (.I0(n3247), .I1(n3253), .I2(n3245), .I3(n3244), 
            .O(n43_adj_5308));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF h2_56 (.Q(PIN_21_c), .C(clk32MHz), .D(hall2));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(clk32MHz), .D(displacement_23__N_80[0]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_IO hall2_input (.PACKAGE_PIN(PIN_4), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(PIN_5), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(PIN_12), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), 
          .D_OUT_1(GND_net), .D_OUT_0(tx_o)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i13008_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n36556), 
            .I3(GND_net), .O(n17747));   // verilog/coms.v(127[12] 295[6])
    defparam i13008_3_lut.LUT_INIT = 16'hacac;
    SB_DFF h3_57 (.Q(PIN_22_c), .C(clk32MHz), .D(hall3));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF dir_61 (.Q(PIN_23_c), .C(clk32MHz), .D(duty[23]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_LUT4 div_46_unary_minus_2_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4918), .I3(n28816), .O(n8_adj_4696)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15_4_lut (.I0(n3234), .I1(n3237), .I2(n3238), .I3(n3239), 
            .O(n40_adj_5310));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_IO PIN_2_pad (.PACKAGE_PIN(PIN_2), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_2_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_2_pad.PIN_TYPE = 6'b000001;
    defparam PIN_2_pad.PULLUP = 1'b0;
    defparam PIN_2_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_2_pad.IO_STANDARD = "SB_LVCMOS";
    neopixel nx (.\neo_pixel_transmitter.done (\neo_pixel_transmitter.done ), 
            .clk32MHz(clk32MHz), .\state_3__N_362[1] (state_3__N_362[1]), 
            .\state[1] (state[1]), .n40674(n40674), .GND_net(GND_net), 
            .bit_ctr({bit_ctr}), .VCC_net(VCC_net), .n33653(n33653), .n33655(n33655), 
            .n33657(n33657), .n33659(n33659), .n33661(n33661), .n33663(n33663), 
            .n33665(n33665), .n33635(n33635), .n33639(n33639), .n33641(n33641), 
            .n33643(n33643), .n33645(n33645), .n33647(n33647), .n18307(n18307), 
            .n33589(n33589), .n33673(n33673), .n33623(n33623), .n33667(n33667), 
            .n33669(n33669), .n33671(n33671), .n33649(n33649), .n33651(n33651), 
            .n33631(n33631), .n33633(n33633), .n33595(n33595), .n18212(n18212), 
            .n33601(n33601), .n33621(n33621), .timer({timer}), .n40726(n40726), 
            .n25779(n25779), .n40725(n40725), .n40724(n40724), .n40723(n40723), 
            .n40722(n40722), .n40721(n40721), .n40720(n40720), .n40719(n40719), 
            .n3209(n3209_adj_5249), .n40718(n40718), .n40717(n40717), 
            .n40716(n40716), .n40715(n40715), .n40714(n40714), .n40713(n40713), 
            .n33619(n33619), .n33617(n33617), .n33629(n33629), .n17687(n17687), 
            .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), .n17686(n17686), 
            .n17685(n17685), .n17684(n17684), .n17683(n17683), .n17682(n17682), 
            .n17681(n17681), .n17680(n17680), .n17679(n17679), .n17678(n17678), 
            .n17677(n17677), .n17676(n17676), .n17675(n17675), .n17674(n17674), 
            .n17673(n17673), .n17672(n17672), .n17671(n17671), .n17670(n17670), 
            .n17669(n17669), .n17668(n17668), .n17667(n17667), .n17666(n17666), 
            .n17665(n17665), .n17664(n17664), .n17663(n17663), .n17662(n17662), 
            .n17661(n17661), .n17660(n17660), .n17659(n17659), .n17658(n17658), 
            .n17657(n17657), .start(start), .\one_wire_N_513[9] (one_wire_N_513[9]), 
            .\one_wire_N_513[10] (one_wire_N_513[10]), .\one_wire_N_513[6] (one_wire_N_513[6]), 
            .\one_wire_N_513[8] (one_wire_N_513[8]), .n11(n11_adj_5254), 
            .\one_wire_N_513[11] (one_wire_N_513[11]), .n4451(n4451), .n1164(n1164), 
            .\state[0] (state[0]), .n4483(n4483), .n40712(n40712), .n35873(n35873), 
            .n40709(n40709), .n40708(n40708), .n17625(n17625), .\state_3__N_362[0] (state_3__N_362[0]), 
            .n17203(n17203), .n35833(n35833), .n40704(n40704), .n40703(n40703), 
            .n17458(n17458), .PIN_8_c(PIN_8_c), .n37483(n37483), .n40702(n40702), 
            .n40700(n40700), .n33675(n33675), .n17444(n17444), .n40699(n40699), 
            .n40698(n40698), .n40707(n40707), .n40706(n40706), .n40701(n40701), 
            .n40711(n40711), .n40710(n40710), .n40705(n40705), .n40619(n40619), 
            .n40620(n40620), .n40616(n40616), .n24984(n24984), .n24782(n24782), 
            .n24824(n24824), .n36533(n36533)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(76[10] 82[2])
    SB_IO hall1_input (.PACKAGE_PIN(PIN_3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis lattice_noprune=1, syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY rem_4_add_849_3 (.CI(n29032), .I0(n1257), .I1(VCC_net), .CO(n29033));
    SB_LUT4 i21_4_lut (.I0(n3240), .I1(n42_adj_5309), .I2(n32_adj_5313), 
            .I3(n3241), .O(n46_adj_5307));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_add_849_2_lut (.I0(GND_net), .I1(n1258), .I2(GND_net), 
            .I3(VCC_net), .O(n1325)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_2 (.CI(VCC_net), .I0(n1258), .I1(GND_net), 
            .CO(n29032));
    SB_LUT4 div_46_unary_minus_4_inv_0_i3_1_lut (.I0(gearBoxRatio[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4909));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY div_46_unary_minus_2_add_3_19 (.CI(n28816), .I0(GND_net), .I1(n8_adj_4918), 
            .CO(n28817));
    SB_LUT4 i13009_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n36556), 
            .I3(GND_net), .O(n17748));   // verilog/coms.v(127[12] 295[6])
    defparam i13009_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_2_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4919), .I3(n28815), .O(n9_adj_4695)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_18 (.CI(n28815), .I0(GND_net), .I1(n9_adj_4919), 
            .CO(n28816));
    SB_LUT4 i13010_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n36556), 
            .I3(GND_net), .O(n17749));   // verilog/coms.v(127[12] 295[6])
    defparam i13010_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut (.I0(n1164), .I1(n40674), .I2(state[0]), .I3(n4451), 
            .O(n25779));   // verilog/neopixel.v(35[12] 117[6])
    defparam i1_4_lut.LUT_INIT = 16'h0535;
    SB_LUT4 div_46_unary_minus_2_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4920), .I3(n28814), .O(n10_adj_4708)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_17 (.CI(n28814), .I0(GND_net), .I1(n10_adj_4920), 
            .CO(n28815));
    SB_LUT4 i13011_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n36556), 
            .I3(GND_net), .O(n17750));   // verilog/coms.v(127[12] 295[6])
    defparam i13011_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i14_4_lut (.I0(n3232), .I1(n3235), .I2(n3233), .I3(n3236), 
            .O(n39_adj_5311));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n43_adj_5308), .I1(n3246), .I2(n38_adj_5312), 
            .I3(n3249), .O(n47));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_unary_minus_4_inv_0_i4_1_lut (.I0(gearBoxRatio[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n22_adj_4908));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i5_1_lut (.I0(gearBoxRatio[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4907));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i6_1_lut (.I0(gearBoxRatio[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4906));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i24_4_lut (.I0(n47), .I1(n39_adj_5311), .I2(n46_adj_5307), 
            .I3(n40_adj_5310), .O(n3263));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13012_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n36556), 
            .I3(GND_net), .O(n17751));   // verilog/coms.v(127[12] 295[6])
    defparam i13012_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_add_1184_16_lut (.I0(n1778_adj_4812), .I1(n1745), .I2(VCC_net), 
            .I3(n29031), .O(n1844)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_46_unary_minus_2_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4921), .I3(n28813), .O(n11_adj_4707)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_15_lut (.I0(GND_net), .I1(n1746), .I2(VCC_net), 
            .I3(n29030), .O(n1813)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_15 (.CI(n29030), .I0(n1746), .I1(VCC_net), 
            .CO(n29031));
    SB_LUT4 rem_4_add_1184_14_lut (.I0(GND_net), .I1(n1747), .I2(VCC_net), 
            .I3(n29029), .O(n1814)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_16 (.CI(n28813), .I0(GND_net), .I1(n11_adj_4921), 
            .CO(n28814));
    SB_LUT4 div_46_unary_minus_2_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4922), .I3(n28812), .O(n12_adj_4698)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_14 (.CI(n29029), .I0(n1747), .I1(VCC_net), 
            .CO(n29030));
    SB_CARRY div_46_unary_minus_2_add_3_15 (.CI(n28812), .I0(GND_net), .I1(n12_adj_4922), 
            .CO(n28813));
    SB_LUT4 div_46_unary_minus_2_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4923), .I3(n28811), .O(n13_adj_4697)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_13_lut (.I0(GND_net), .I1(n1748), .I2(VCC_net), 
            .I3(n29028), .O(n1815)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_13 (.CI(n29028), .I0(n1748), .I1(VCC_net), 
            .CO(n29029));
    SB_CARRY div_46_unary_minus_2_add_3_14 (.CI(n28811), .I0(GND_net), .I1(n13_adj_4923), 
            .CO(n28812));
    SB_LUT4 div_46_unary_minus_2_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4924), .I3(n28810), .O(n14_adj_4710)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_12_lut (.I0(GND_net), .I1(n1749), .I2(VCC_net), 
            .I3(n29027), .O(n1816)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_13 (.CI(n28810), .I0(GND_net), .I1(n14_adj_4924), 
            .CO(n28811));
    SB_CARRY rem_4_add_1184_12 (.CI(n29027), .I0(n1749), .I1(VCC_net), 
            .CO(n29028));
    SB_LUT4 div_46_unary_minus_2_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4925), .I3(n28809), .O(n15_adj_4709)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_11_lut (.I0(GND_net), .I1(n1750), .I2(VCC_net), 
            .I3(n29026), .O(n1817)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_12 (.CI(n28809), .I0(GND_net), .I1(n15_adj_4925), 
            .CO(n28810));
    SB_CARRY rem_4_add_1184_11 (.CI(n29026), .I0(n1750), .I1(VCC_net), 
            .CO(n29027));
    SB_LUT4 div_46_unary_minus_2_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4926), .I3(n28808), .O(n16_adj_4703)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_11 (.CI(n28808), .I0(GND_net), .I1(n16_adj_4926), 
            .CO(n28809));
    SB_LUT4 rem_4_add_1184_10_lut (.I0(GND_net), .I1(n1751), .I2(VCC_net), 
            .I3(n29025), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4927), .I3(n28807), .O(n17_adj_4702)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_10 (.CI(n29025), .I0(n1751), .I1(VCC_net), 
            .CO(n29026));
    SB_CARRY div_46_unary_minus_2_add_3_10 (.CI(n28807), .I0(GND_net), .I1(n17_adj_4927), 
            .CO(n28808));
    SB_LUT4 rem_4_add_1184_9_lut (.I0(GND_net), .I1(n1752), .I2(VCC_net), 
            .I3(n29024), .O(n1819)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4928), .I3(n28806), .O(n18_adj_4701)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_9 (.CI(n29024), .I0(n1752), .I1(VCC_net), 
            .CO(n29025));
    SB_CARRY div_46_unary_minus_2_add_3_9 (.CI(n28806), .I0(GND_net), .I1(n18_adj_4928), 
            .CO(n28807));
    SB_LUT4 div_46_unary_minus_2_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4929), .I3(n28805), .O(n19_adj_4700)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_8_lut (.I0(GND_net), .I1(n1753), .I2(VCC_net), 
            .I3(n29023), .O(n1820)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_8 (.CI(n29023), .I0(n1753), .I1(VCC_net), 
            .CO(n29024));
    SB_CARRY div_46_unary_minus_2_add_3_8 (.CI(n28805), .I0(GND_net), .I1(n19_adj_4929), 
            .CO(n28806));
    SB_LUT4 rem_4_add_1184_7_lut (.I0(GND_net), .I1(n1754_adj_4807), .I2(GND_net), 
            .I3(n29022), .O(n1821)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4930), .I3(n28804), .O(n20_adj_4699)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_7 (.CI(n28804), .I0(GND_net), .I1(n20_adj_4930), 
            .CO(n28805));
    SB_CARRY rem_4_add_1184_7 (.CI(n29022), .I0(n1754_adj_4807), .I1(GND_net), 
            .CO(n29023));
    SB_LUT4 div_46_unary_minus_2_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4931), .I3(n28803), .O(n21_adj_4666)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_6_lut (.I0(GND_net), .I1(n1755_adj_4808), .I2(GND_net), 
            .I3(n29021), .O(n1822)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_6 (.CI(n28803), .I0(GND_net), .I1(n21_adj_4931), 
            .CO(n28804));
    SB_CARRY rem_4_add_1184_6 (.CI(n29021), .I0(n1755_adj_4808), .I1(GND_net), 
            .CO(n29022));
    SB_LUT4 div_46_unary_minus_2_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4932), .I3(n28802), .O(n22_adj_4714)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1184_5_lut (.I0(GND_net), .I1(n1756_adj_4809), .I2(VCC_net), 
            .I3(n29020), .O(n1823)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_5 (.CI(n28802), .I0(GND_net), .I1(n22_adj_4932), 
            .CO(n28803));
    SB_LUT4 i13013_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n36556), 
            .I3(GND_net), .O(n17752));   // verilog/coms.v(127[12] 295[6])
    defparam i13013_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13014_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n36556), 
            .I3(GND_net), .O(n17753));   // verilog/coms.v(127[12] 295[6])
    defparam i13014_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i2148_3_lut (.I0(n3155), .I1(n3222), .I2(n3164), .I3(GND_net), 
            .O(n3254));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13015_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n36556), 
            .I3(GND_net), .O(n17754));   // verilog/coms.v(127[12] 295[6])
    defparam i13015_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13016_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n36556), 
            .I3(GND_net), .O(n17755));   // verilog/coms.v(127[12] 295[6])
    defparam i13016_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_4_inv_0_i7_1_lut (.I0(gearBoxRatio[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4905));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2215_3_lut (.I0(n3254), .I1(n3321), .I2(n3263), .I3(GND_net), 
            .O(n3353));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2215_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13017_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n36556), 
            .I3(GND_net), .O(n17756));   // verilog/coms.v(127[12] 295[6])
    defparam i13017_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13018_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n36556), 
            .I3(GND_net), .O(n17757));   // verilog/coms.v(127[12] 295[6])
    defparam i13018_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_4_inv_0_i8_1_lut (.I0(gearBoxRatio[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4904));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13019_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n36556), 
            .I3(GND_net), .O(n17758));   // verilog/coms.v(127[12] 295[6])
    defparam i13019_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13020_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n36556), 
            .I3(GND_net), .O(n17759));   // verilog/coms.v(127[12] 295[6])
    defparam i13020_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13021_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n36556), 
            .I3(GND_net), .O(n17760));   // verilog/coms.v(127[12] 295[6])
    defparam i13021_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13022_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n36556), 
            .I3(GND_net), .O(n17761));   // verilog/coms.v(127[12] 295[6])
    defparam i13022_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_4_inv_0_i9_1_lut (.I0(gearBoxRatio[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4903));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13023_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n36556), 
            .I3(GND_net), .O(n17762));   // verilog/coms.v(127[12] 295[6])
    defparam i13023_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_4_inv_0_i10_1_lut (.I0(gearBoxRatio[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4902));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13024_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n36556), 
            .I3(GND_net), .O(n17763));   // verilog/coms.v(127[12] 295[6])
    defparam i13024_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_4_inv_0_i11_1_lut (.I0(gearBoxRatio[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4901));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13025_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n36556), 
            .I3(GND_net), .O(n17764));   // verilog/coms.v(127[12] 295[6])
    defparam i13025_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1262_3_lut (.I0(n1853), .I1(n1920), .I2(n1877), .I3(GND_net), 
            .O(n1952));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1262_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13026_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n36556), 
            .I3(GND_net), .O(n17765));   // verilog/coms.v(127[12] 295[6])
    defparam i13026_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1259_3_lut (.I0(n1850), .I1(n1917), .I2(n1877), .I3(GND_net), 
            .O(n1949));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1259_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13027_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n36556), 
            .I3(GND_net), .O(n17766));   // verilog/coms.v(127[12] 295[6])
    defparam i13027_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1260_3_lut (.I0(n1851), .I1(n1918), .I2(n1877), .I3(GND_net), 
            .O(n1950));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1260_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13028_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n36556), 
            .I3(GND_net), .O(n17767));   // verilog/coms.v(127[12] 295[6])
    defparam i13028_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1258_3_lut (.I0(n1849), .I1(n1916), .I2(n1877), .I3(GND_net), 
            .O(n1948));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1258_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1263_3_lut (.I0(n1854), .I1(n1921), .I2(n1877), .I3(GND_net), 
            .O(n1953));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1263_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1261_3_lut (.I0(n1852), .I1(n1919), .I2(n1877), .I3(GND_net), 
            .O(n1951));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1261_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1256_3_lut (.I0(n1847), .I1(n1914), .I2(n1877), .I3(GND_net), 
            .O(n1946));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1256_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13029_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n36556), 
            .I3(GND_net), .O(n17768));   // verilog/coms.v(127[12] 295[6])
    defparam i13029_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1255_3_lut (.I0(n1846), .I1(n1913), .I2(n1877), .I3(GND_net), 
            .O(n1945));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1255_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1254_3_lut (.I0(n1845), .I1(n1912), .I2(n1877), .I3(GND_net), 
            .O(n1944));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1254_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF color__i11 (.Q(color[11]), .C(LED_c), .D(n18223));   // verilog/TinyFPGA_B.v(51[8] 74[4])
    SB_DFF color__i12 (.Q(color[12]), .C(LED_c), .D(n32167));   // verilog/TinyFPGA_B.v(51[8] 74[4])
    SB_LUT4 i13030_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17769));   // verilog/coms.v(127[12] 295[6])
    defparam i13030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13031_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17770));   // verilog/coms.v(127[12] 295[6])
    defparam i13031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1265_3_lut (.I0(n1856), .I1(n1923), .I2(n1877), .I3(GND_net), 
            .O(n1955));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1265_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF color__i10 (.Q(color[10]), .C(LED_c), .D(n18222));   // verilog/TinyFPGA_B.v(51[8] 74[4])
    SB_DFF color__i9 (.Q(color[9]), .C(LED_c), .D(n18215));   // verilog/TinyFPGA_B.v(51[8] 74[4])
    SB_LUT4 rem_4_i1264_3_lut (.I0(n1855), .I1(n1922), .I2(n1877), .I3(GND_net), 
            .O(n1954));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1264_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1257_3_lut (.I0(n1848), .I1(n1915), .I2(n1877), .I3(GND_net), 
            .O(n1947));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1257_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1267_3_lut (.I0(n1858), .I1(n1925), .I2(n1877), .I3(GND_net), 
            .O(n1957));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1267_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1266_3_lut (.I0(n1857), .I1(n1924), .I2(n1877), .I3(GND_net), 
            .O(n1956));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1266_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(n1956), .I1(n1957), .I2(n1958), .I3(GND_net), 
            .O(n35991));
    defparam i1_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut (.I0(n1947), .I1(n1954), .I2(n35991), .I3(n1955), 
            .O(n15_adj_5317));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i3_4_lut.LUT_INIT = 16'heaaa;
    SB_LUT4 i13032_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17771));   // verilog/coms.v(127[12] 295[6])
    defparam i13032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut (.I0(n1944), .I1(n1945), .I2(n1943), .I3(n1946), 
            .O(n19_adj_5315));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(n1951), .I1(n1953), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_5316));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut (.I0(n19_adj_5315), .I1(n15_adj_5317), .I2(n1948), 
            .I3(n1950), .O(n22_adj_5314));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n1949), .I1(n22_adj_5314), .I2(n18_adj_5316), 
            .I3(n1952), .O(n1976_adj_4779));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 unary_minus_28_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_mux_3_i17_3_lut (.I0(communication_counter[16]), .I1(n17_adj_4792), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1958));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1768_3_lut_3_lut (.I0(n2642), .I1(n6207), .I2(n2632), 
            .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1768_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13169_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n13302), .I3(GND_net), .O(n17908));   // verilog/coms.v(127[12] 295[6])
    defparam i13169_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1184_5 (.CI(n29020), .I0(n1756_adj_4809), .I1(VCC_net), 
            .CO(n29021));
    SB_LUT4 div_46_unary_minus_4_inv_0_i12_1_lut (.I0(gearBoxRatio[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4900));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13033_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17772));   // verilog/coms.v(127[12] 295[6])
    defparam i13033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i13_1_lut (.I0(gearBoxRatio[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4899));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13034_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17773));   // verilog/coms.v(127[12] 295[6])
    defparam i13034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1755_3_lut_3_lut (.I0(n2642), .I1(n6194), .I2(n2619), 
            .I3(GND_net), .O(n2700));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1755_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13035_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17774));   // verilog/coms.v(127[12] 295[6])
    defparam i13035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i14_1_lut (.I0(gearBoxRatio[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_4898));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i15_1_lut (.I0(gearBoxRatio[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4897));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13036_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17775));   // verilog/coms.v(127[12] 295[6])
    defparam i13036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13037_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17776));   // verilog/coms.v(127[12] 295[6])
    defparam i13037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13038_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17777));   // verilog/coms.v(127[12] 295[6])
    defparam i13038_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13039_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17778));   // verilog/coms.v(127[12] 295[6])
    defparam i13039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1754_3_lut_3_lut (.I0(n2642), .I1(n6193), .I2(n2618), 
            .I3(GND_net), .O(n2699));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1754_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1757_3_lut_3_lut (.I0(n2642), .I1(n6196), .I2(n2621), 
            .I3(GND_net), .O(n2702));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1757_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13040_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17779));   // verilog/coms.v(127[12] 295[6])
    defparam i13040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13041_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17780));   // verilog/coms.v(127[12] 295[6])
    defparam i13041_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1758_3_lut_3_lut (.I0(n2642), .I1(n6197), .I2(n2622), 
            .I3(GND_net), .O(n2703));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1758_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1756_3_lut_3_lut (.I0(n2642), .I1(n6195), .I2(n2620), 
            .I3(GND_net), .O(n2701));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1756_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_4_inv_0_i16_1_lut (.I0(gearBoxRatio[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4896));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13042_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17781));   // verilog/coms.v(127[12] 295[6])
    defparam i13042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13043_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17782));   // verilog/coms.v(127[12] 295[6])
    defparam i13043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13044_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17783));   // verilog/coms.v(127[12] 295[6])
    defparam i13044_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13045_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17784));   // verilog/coms.v(127[12] 295[6])
    defparam i13045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13170_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n13302), .I3(GND_net), .O(n17909));   // verilog/coms.v(127[12] 295[6])
    defparam i13170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4933), .I3(n28801), .O(n23_adj_4713)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13046_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17785));   // verilog/coms.v(127[12] 295[6])
    defparam i13046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13047_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17786));   // verilog/coms.v(127[12] 295[6])
    defparam i13047_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i17_1_lut (.I0(gearBoxRatio[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4895));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13048_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17787));   // verilog/coms.v(127[12] 295[6])
    defparam i13048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13049_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17788));   // verilog/coms.v(127[12] 295[6])
    defparam i13049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1761_3_lut_3_lut (.I0(n2642), .I1(n6200), .I2(n2625), 
            .I3(GND_net), .O(n2706));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1761_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13050_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17789));   // verilog/coms.v(127[12] 295[6])
    defparam i13050_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13051_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17790));   // verilog/coms.v(127[12] 295[6])
    defparam i13051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13052_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17791));   // verilog/coms.v(127[12] 295[6])
    defparam i13052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13053_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17792));   // verilog/coms.v(127[12] 295[6])
    defparam i13053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1184_4_lut (.I0(GND_net), .I1(n1757_adj_4810), .I2(VCC_net), 
            .I3(n29019), .O(n1824)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1184_4 (.CI(n29019), .I0(n1757_adj_4810), .I1(VCC_net), 
            .CO(n29020));
    SB_LUT4 div_46_unary_minus_4_inv_0_i18_1_lut (.I0(gearBoxRatio[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4894));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13171_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n13302), .I3(GND_net), .O(n17910));   // verilog/coms.v(127[12] 295[6])
    defparam i13171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13172_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n13302), .I3(GND_net), .O(n17911));   // verilog/coms.v(127[12] 295[6])
    defparam i13172_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13054_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17793));   // verilog/coms.v(127[12] 295[6])
    defparam i13054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13055_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17794));   // verilog/coms.v(127[12] 295[6])
    defparam i13055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13173_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n13302), .I3(GND_net), .O(n17912));   // verilog/coms.v(127[12] 295[6])
    defparam i13173_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1184_3_lut (.I0(GND_net), .I1(n1758_adj_4811), .I2(GND_net), 
            .I3(n29018), .O(n1825)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1184_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13056_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17795));   // verilog/coms.v(127[12] 295[6])
    defparam i13056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13057_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17796));   // verilog/coms.v(127[12] 295[6])
    defparam i13057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13058_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17797));   // verilog/coms.v(127[12] 295[6])
    defparam i13058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13059_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17798));   // verilog/coms.v(127[12] 295[6])
    defparam i13059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13174_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n13302), .I3(GND_net), .O(n17913));   // verilog/coms.v(127[12] 295[6])
    defparam i13174_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_46_unary_minus_2_add_3_4 (.CI(n28801), .I0(GND_net), .I1(n23_adj_4933), 
            .CO(n28802));
    SB_LUT4 i13060_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17799));   // verilog/coms.v(127[12] 295[6])
    defparam i13060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13061_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n13302), .I3(GND_net), .O(n17800));   // verilog/coms.v(127[12] 295[6])
    defparam i13061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13175_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n13302), .I3(GND_net), .O(n17914));   // verilog/coms.v(127[12] 295[6])
    defparam i13175_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13062_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n13302), .I3(GND_net), .O(n17801));   // verilog/coms.v(127[12] 295[6])
    defparam i13062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13176_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n13302), .I3(GND_net), .O(n17915));   // verilog/coms.v(127[12] 295[6])
    defparam i13176_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13063_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n13302), .I3(GND_net), .O(n17802));   // verilog/coms.v(127[12] 295[6])
    defparam i13063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i19_1_lut (.I0(gearBoxRatio[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4893));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13064_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n13302), .I3(GND_net), .O(n17803));   // verilog/coms.v(127[12] 295[6])
    defparam i13064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13177_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n13302), .I3(GND_net), .O(n17916));   // verilog/coms.v(127[12] 295[6])
    defparam i13177_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13065_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n13302), .I3(GND_net), .O(n17804));   // verilog/coms.v(127[12] 295[6])
    defparam i13065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13066_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n13302), .I3(GND_net), .O(n17805));   // verilog/coms.v(127[12] 295[6])
    defparam i13066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13178_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n13302), .I3(GND_net), .O(n17917));   // verilog/coms.v(127[12] 295[6])
    defparam i13178_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13167_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n13302), .I3(GND_net), .O(n17906));   // verilog/coms.v(127[12] 295[6])
    defparam i13167_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13179_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n13302), .I3(GND_net), .O(n17918));   // verilog/coms.v(127[12] 295[6])
    defparam i13179_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1184_3 (.CI(n29018), .I0(n1758_adj_4811), .I1(GND_net), 
            .CO(n29019));
    SB_LUT4 div_46_unary_minus_2_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4934), .I3(n28800), .O(n24_adj_4712)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13180_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n13302), .I3(GND_net), .O(n17919));   // verilog/coms.v(127[12] 295[6])
    defparam i13180_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13181_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n13302), .I3(GND_net), .O(n17920));   // verilog/coms.v(127[12] 295[6])
    defparam i13181_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13182_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n13302), .I3(GND_net), .O(n17921));   // verilog/coms.v(127[12] 295[6])
    defparam i13182_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1762_3_lut_3_lut (.I0(n2642), .I1(n6201), .I2(n2626), 
            .I3(GND_net), .O(n2707));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1762_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13183_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n13302), .I3(GND_net), .O(n17922));   // verilog/coms.v(127[12] 295[6])
    defparam i13183_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1759_3_lut_3_lut (.I0(n2642), .I1(n6198), .I2(n2623), 
            .I3(GND_net), .O(n2704));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1759_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13168_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n13302), .I3(GND_net), .O(n17907));   // verilog/coms.v(127[12] 295[6])
    defparam i13168_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13184_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n13302), .I3(GND_net), .O(n17923));   // verilog/coms.v(127[12] 295[6])
    defparam i13184_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13067_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n13302), .I3(GND_net), .O(n17806));   // verilog/coms.v(127[12] 295[6])
    defparam i13067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13185_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n13302), .I3(GND_net), .O(n17924));   // verilog/coms.v(127[12] 295[6])
    defparam i13185_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13186_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n13302), .I3(GND_net), .O(n17925));   // verilog/coms.v(127[12] 295[6])
    defparam i13186_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13187_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n13302), .I3(GND_net), .O(n17926));   // verilog/coms.v(127[12] 295[6])
    defparam i13187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1766_3_lut_3_lut (.I0(n2642), .I1(n6205), .I2(n2630), 
            .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1766_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13068_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n13302), .I3(GND_net), .O(n17807));   // verilog/coms.v(127[12] 295[6])
    defparam i13068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1767_3_lut_3_lut (.I0(n2642), .I1(n6206), .I2(n2631), 
            .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1767_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13188_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n13302), .I3(GND_net), .O(n17927));   // verilog/coms.v(127[12] 295[6])
    defparam i13188_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13189_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n4593), .I3(GND_net), .O(n17928));   // verilog/coms.v(127[12] 295[6])
    defparam i13189_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_46_unary_minus_2_add_3_3 (.CI(n28800), .I0(GND_net), .I1(n24_adj_4934), 
            .CO(n28801));
    SB_LUT4 i13190_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n4593), .I3(GND_net), .O(n17929));   // verilog/coms.v(127[12] 295[6])
    defparam i13190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13191_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n4593), .I3(GND_net), .O(n17930));   // verilog/coms.v(127[12] 295[6])
    defparam i13191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i20_1_lut (.I0(gearBoxRatio[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4892));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 PIN_13_I_0_1_lut (.I0(PIN_13_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(PIN_13_N_105));   // verilog/TinyFPGA_B.v(189[10:15])
    defparam PIN_13_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1760_3_lut_3_lut (.I0(n2642), .I1(n6199), .I2(n2624), 
            .I3(GND_net), .O(n2705));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1760_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_4_inv_0_i21_1_lut (.I0(gearBoxRatio[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4891));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13192_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n4593), .I3(GND_net), .O(n17931));   // verilog/coms.v(127[12] 295[6])
    defparam i13192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13193_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n4593), .I3(GND_net), .O(n17932));   // verilog/coms.v(127[12] 295[6])
    defparam i13193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13194_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n4593), .I3(GND_net), .O(n17933));   // verilog/coms.v(127[12] 295[6])
    defparam i13194_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1184_2 (.CI(VCC_net), .I0(n1858), .I1(VCC_net), 
            .CO(n29018));
    SB_LUT4 rem_4_add_1251_17_lut (.I0(n1877), .I1(n1844), .I2(VCC_net), 
            .I3(n29017), .O(n1943)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_46_unary_minus_2_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4935), .I3(VCC_net), .O(n25_adj_4711)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_16_lut (.I0(GND_net), .I1(n1845), .I2(VCC_net), 
            .I3(n29016), .O(n1912)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4935), 
            .CO(n28800));
    SB_CARRY rem_4_add_1251_16 (.CI(n29016), .I0(n1845), .I1(VCC_net), 
            .CO(n29017));
    SB_LUT4 rem_4_add_1251_15_lut (.I0(GND_net), .I1(n1846), .I2(VCC_net), 
            .I3(n29015), .O(n1913)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_25_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(n2_adj_4888), .I3(n28799), .O(n77)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_46_unary_minus_4_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4889), .I3(n28798), .O(n53)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_15 (.CI(n29015), .I0(n1846), .I1(VCC_net), 
            .CO(n29016));
    SB_LUT4 rem_4_add_1251_14_lut (.I0(GND_net), .I1(n1847), .I2(VCC_net), 
            .I3(n29014), .O(n1914)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_24 (.CI(n28798), .I0(GND_net), .I1(n3_adj_4889), 
            .CO(n28799));
    SB_LUT4 rem_4_i1870_3_lut (.I0(n2749), .I1(n2816), .I2(n2768), .I3(GND_net), 
            .O(n2848));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1870_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1775_3_lut_3_lut (.I0(n2642), .I1(n6214), .I2(n1064), 
            .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1775_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1251_14 (.CI(n29014), .I0(n1847), .I1(VCC_net), 
            .CO(n29015));
    SB_LUT4 div_46_unary_minus_4_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4890), .I3(n28797), .O(n54)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_13_lut (.I0(GND_net), .I1(n1848), .I2(VCC_net), 
            .I3(n29013), .O(n1915)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1765_3_lut_3_lut (.I0(n2642), .I1(n6204), .I2(n2629), 
            .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1765_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1874_rep_29_3_lut (.I0(n2753), .I1(n2820), .I2(n2768), 
            .I3(GND_net), .O(n2852));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1874_rep_29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1866_3_lut (.I0(n2745), .I1(n2812), .I2(n2768), .I3(GND_net), 
            .O(n2844));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1866_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1251_13 (.CI(n29013), .I0(n1848), .I1(VCC_net), 
            .CO(n29014));
    SB_CARRY div_46_unary_minus_4_add_3_23 (.CI(n28797), .I0(GND_net), .I1(n4_adj_4890), 
            .CO(n28798));
    SB_LUT4 rem_4_add_1251_12_lut (.I0(GND_net), .I1(n1849), .I2(VCC_net), 
            .I3(n29012), .O(n1916)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4891), .I3(n28796), .O(n55)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1764_3_lut_3_lut (.I0(n2642), .I1(n6203), .I2(n2628), 
            .I3(GND_net), .O(n2709));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1764_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY div_46_unary_minus_4_add_3_22 (.CI(n28796), .I0(GND_net), .I1(n5_adj_4891), 
            .CO(n28797));
    SB_CARRY rem_4_add_1251_12 (.CI(n29012), .I0(n1849), .I1(VCC_net), 
            .CO(n29013));
    SB_LUT4 rem_4_add_1251_11_lut (.I0(GND_net), .I1(n1850), .I2(VCC_net), 
            .I3(n29011), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4892), .I3(n28795), .O(n56)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1865_3_lut (.I0(n2744), .I1(n2811), .I2(n2768), .I3(GND_net), 
            .O(n2843));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1865_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1251_11 (.CI(n29011), .I0(n1850), .I1(VCC_net), 
            .CO(n29012));
    SB_CARRY div_46_unary_minus_4_add_3_21 (.CI(n28795), .I0(GND_net), .I1(n6_adj_4892), 
            .CO(n28796));
    SB_LUT4 rem_4_i1871_3_lut (.I0(n2750), .I1(n2817), .I2(n2768), .I3(GND_net), 
            .O(n2849));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1871_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1773_3_lut_3_lut (.I0(n2642), .I1(n6212), .I2(n2637), 
            .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1773_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1875_3_lut (.I0(n2754), .I1(n2821), .I2(n2768), .I3(GND_net), 
            .O(n2853));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1875_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1774_3_lut_3_lut (.I0(n2642), .I1(n6213), .I2(n2638), 
            .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1774_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1251_10_lut (.I0(GND_net), .I1(n1851), .I2(VCC_net), 
            .I3(n29010), .O(n1918)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1872_3_lut (.I0(n2751), .I1(n2818), .I2(n2768), .I3(GND_net), 
            .O(n2850));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1872_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1251_10 (.CI(n29010), .I0(n1851), .I1(VCC_net), 
            .CO(n29011));
    SB_LUT4 div_46_unary_minus_4_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4893), .I3(n28794), .O(n57)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1772_3_lut_3_lut (.I0(n2642), .I1(n6211), .I2(n2636), 
            .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1772_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1863_3_lut (.I0(n2742), .I1(n2809), .I2(n2768), .I3(GND_net), 
            .O(n2841));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1863_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1862_3_lut (.I0(n2741), .I1(n2808), .I2(n2768), .I3(GND_net), 
            .O(n2840));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1862_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1867_3_lut (.I0(n2746), .I1(n2813), .I2(n2768), .I3(GND_net), 
            .O(n2845));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1867_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1869_rep_35_3_lut (.I0(n2748), .I1(n2815), .I2(n2768), 
            .I3(GND_net), .O(n2847));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1869_rep_35_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1770_3_lut_3_lut (.I0(n2642), .I1(n6209), .I2(n2634), 
            .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1770_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i34861_3_lut (.I0(n2747), .I1(n2814), .I2(n2768), .I3(GND_net), 
            .O(n2846));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i34861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34858_3_lut (.I0(n2653), .I1(n2720_adj_4825), .I2(n2669), 
            .I3(GND_net), .O(n2752));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i34858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34859_3_lut (.I0(n2752), .I1(n2819), .I2(n2768), .I3(GND_net), 
            .O(n2851));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i34859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1857_3_lut (.I0(n2736), .I1(n2803), .I2(n2768), .I3(GND_net), 
            .O(n2835));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1251_9_lut (.I0(GND_net), .I1(n1852), .I2(VCC_net), 
            .I3(n29009), .O(n1919)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_9 (.CI(n29009), .I0(n1852), .I1(VCC_net), 
            .CO(n29010));
    SB_CARRY div_46_unary_minus_4_add_3_20 (.CI(n28794), .I0(GND_net), .I1(n7_adj_4893), 
            .CO(n28795));
    SB_LUT4 div_46_i1769_3_lut_3_lut (.I0(n2642), .I1(n6208), .I2(n2633), 
            .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1769_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1861_3_lut (.I0(n2740), .I1(n2807), .I2(n2768), .I3(GND_net), 
            .O(n2839));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1861_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1251_8_lut (.I0(GND_net), .I1(n1853), .I2(VCC_net), 
            .I3(n29008), .O(n1920)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_4894), .I3(n28793), .O(n58)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_8 (.CI(n29008), .I0(n1853), .I1(VCC_net), 
            .CO(n29009));
    SB_CARRY div_46_unary_minus_4_add_3_19 (.CI(n28793), .I0(GND_net), .I1(n8_adj_4894), 
            .CO(n28794));
    SB_LUT4 rem_4_i1859_3_lut (.I0(n2738), .I1(n2805), .I2(n2768), .I3(GND_net), 
            .O(n2837));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1860_3_lut (.I0(n2739), .I1(n2806), .I2(n2768), .I3(GND_net), 
            .O(n2838));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1860_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1858_3_lut (.I0(n2737), .I1(n2804), .I2(n2768), .I3(GND_net), 
            .O(n2836));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_4895), .I3(n28792), .O(n59)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_7_lut (.I0(GND_net), .I1(n1854), .I2(GND_net), 
            .I3(n29007), .O(n1921)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_18 (.CI(n28792), .I0(GND_net), .I1(n9_adj_4895), 
            .CO(n28793));
    SB_LUT4 div_46_unary_minus_4_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_4896), .I3(n28791), .O(n60)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1877_3_lut (.I0(n2756), .I1(n2823), .I2(n2768), .I3(GND_net), 
            .O(n2855));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1877_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1876_3_lut (.I0(n2755), .I1(n2822), .I2(n2768), .I3(GND_net), 
            .O(n2854));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1876_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1864_3_lut (.I0(n2743), .I1(n2810), .I2(n2768), .I3(GND_net), 
            .O(n2842));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1864_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1798_3_lut (.I0(n2645), .I1(n2712_adj_4833), .I2(n2669), 
            .I3(GND_net), .O(n2744));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1798_3_lut.LUT_INIT = 16'hcaca;
    SB_IO PIN_1_pad (.PACKAGE_PIN(PIN_1), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_1_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_1_pad.PIN_TYPE = 6'b000001;
    defparam PIN_1_pad.PULLUP = 1'b0;
    defparam PIN_1_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_1_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 rem_4_i1803_3_lut (.I0(n2650), .I1(n2717_adj_4828), .I2(n2669), 
            .I3(GND_net), .O(n2749));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1804_3_lut (.I0(n2651), .I1(n2718_adj_4827), .I2(n2669), 
            .I3(GND_net), .O(n2750));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1802_3_lut (.I0(n2649), .I1(n2716_adj_4829), .I2(n2669), 
            .I3(GND_net), .O(n2748));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1802_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1805_3_lut (.I0(n2652), .I1(n2719_adj_4826), .I2(n2669), 
            .I3(GND_net), .O(n2751));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1805_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1792_3_lut (.I0(n2639), .I1(n2706_adj_4839), .I2(n2669), 
            .I3(GND_net), .O(n2738));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1792_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1791_3_lut (.I0(n2638_adj_4845), .I1(n2705_adj_4840), 
            .I2(n2669), .I3(GND_net), .O(n2737));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1790_3_lut (.I0(n2637_adj_4846), .I1(n2704_adj_4841), 
            .I2(n2669), .I3(GND_net), .O(n2736));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1796_3_lut (.I0(n2643_adj_4843), .I1(n2710_adj_4835), 
            .I2(n2669), .I3(GND_net), .O(n2742));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1796_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1794_3_lut (.I0(n2641), .I1(n2708_adj_4837), .I2(n2669), 
            .I3(GND_net), .O(n2740));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1794_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1795_3_lut (.I0(n2642_adj_4844), .I1(n2709_adj_4836), 
            .I2(n2669), .I3(GND_net), .O(n2741));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1795_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1793_3_lut (.I0(n2640), .I1(n2707_adj_4838), .I2(n2669), 
            .I3(GND_net), .O(n2739));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1793_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1763_3_lut_3_lut (.I0(n2642), .I1(n6202), .I2(n2627), 
            .I3(GND_net), .O(n2708));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1763_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1809_3_lut (.I0(n2656), .I1(n2723_adj_4824), .I2(n2669), 
            .I3(GND_net), .O(n2755));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1808_3_lut (.I0(n2655), .I1(n2722), .I2(n2669), .I3(GND_net), 
            .O(n2754));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1808_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_46_unary_minus_4_add_3_17 (.CI(n28791), .I0(GND_net), .I1(n10_adj_4896), 
            .CO(n28792));
    SB_LUT4 div_46_i1771_3_lut_3_lut (.I0(n2642), .I1(n6210), .I2(n2635), 
            .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1771_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1251_7 (.CI(n29007), .I0(n1854), .I1(GND_net), 
            .CO(n29008));
    SB_LUT4 rem_4_add_1251_6_lut (.I0(GND_net), .I1(n1855), .I2(GND_net), 
            .I3(n29006), .O(n1922)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_4897), .I3(n28790), .O(n61)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_16 (.CI(n28790), .I0(GND_net), .I1(n11_adj_4897), 
            .CO(n28791));
    SB_LUT4 div_46_unary_minus_4_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_4898), .I3(n28789), .O(n62)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_6 (.CI(n29006), .I0(n1855), .I1(GND_net), 
            .CO(n29007));
    SB_LUT4 rem_4_add_1251_5_lut (.I0(GND_net), .I1(n1856), .I2(VCC_net), 
            .I3(n29005), .O(n1923)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_5 (.CI(n29005), .I0(n1856), .I1(VCC_net), 
            .CO(n29006));
    SB_CARRY div_46_unary_minus_4_add_3_15 (.CI(n28789), .I0(GND_net), .I1(n12_adj_4898), 
            .CO(n28790));
    SB_LUT4 div_46_unary_minus_4_inv_0_i22_1_lut (.I0(gearBoxRatio[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4890));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_24_pad (.PACKAGE_PIN(PIN_24), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_24_pad.PIN_TYPE = 6'b011001;
    defparam PIN_24_pad.PULLUP = 1'b0;
    defparam PIN_24_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_24_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_23_pad (.PACKAGE_PIN(PIN_23), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_23_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_23_pad.PIN_TYPE = 6'b011001;
    defparam PIN_23_pad.PULLUP = 1'b0;
    defparam PIN_23_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_23_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_22_pad (.PACKAGE_PIN(PIN_22), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_22_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_22_pad.PIN_TYPE = 6'b011001;
    defparam PIN_22_pad.PULLUP = 1'b0;
    defparam PIN_22_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_22_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_6_pad (.PACKAGE_PIN(PIN_6), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_6_c_1)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_6_pad.PIN_TYPE = 6'b000001;
    defparam PIN_6_pad.PULLUP = 1'b0;
    defparam PIN_6_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_6_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 rem_4_i1797_3_lut (.I0(n2644), .I1(n2711_adj_4834), .I2(n2669), 
            .I3(GND_net), .O(n2743));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1797_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1251_4_lut (.I0(GND_net), .I1(n1857), .I2(VCC_net), 
            .I3(n29004), .O(n1924)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_4899), .I3(n28788), .O(n63)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_14 (.CI(n28788), .I0(GND_net), .I1(n13_adj_4899), 
            .CO(n28789));
    SB_CARRY rem_4_add_1251_4 (.CI(n29004), .I0(n1857), .I1(VCC_net), 
            .CO(n29005));
    SB_LUT4 div_46_unary_minus_4_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_4900), .I3(n28787), .O(n64)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1251_3_lut (.I0(GND_net), .I1(n1858), .I2(GND_net), 
            .I3(n29003), .O(n1925)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1251_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1251_3 (.CI(n29003), .I0(n1858), .I1(GND_net), 
            .CO(n29004));
    SB_CARRY div_46_unary_minus_4_add_3_13 (.CI(n28787), .I0(GND_net), .I1(n14_adj_4900), 
            .CO(n28788));
    SB_LUT4 rem_4_i1801_3_lut (.I0(n2648), .I1(n2715_adj_4830), .I2(n2669), 
            .I3(GND_net), .O(n2747));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1807_3_lut (.I0(n2654), .I1(n2721), .I2(n2669), .I3(GND_net), 
            .O(n2753));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1799_3_lut (.I0(n2646), .I1(n2713_adj_4832), .I2(n2669), 
            .I3(GND_net), .O(n2745));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1799_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1251_2 (.CI(VCC_net), .I0(n1958), .I1(VCC_net), 
            .CO(n29003));
    SB_LUT4 rem_4_add_1318_18_lut (.I0(n1976_adj_4779), .I1(n1943), .I2(VCC_net), 
            .I3(n29002), .O(n2042)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_46_unary_minus_4_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_4901), .I3(n28786), .O(n65)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1800_3_lut (.I0(n2647), .I1(n2714_adj_4831), .I2(n2669), 
            .I3(GND_net), .O(n2746));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1800_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_46_unary_minus_4_add_3_12 (.CI(n28786), .I0(GND_net), .I1(n15_adj_4901), 
            .CO(n28787));
    SB_LUT4 div_46_unary_minus_4_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_4902), .I3(n28785), .O(n66)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1318_17_lut (.I0(GND_net), .I1(n1944), .I2(VCC_net), 
            .I3(n29001), .O(n2011)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1730_3_lut (.I0(n2545_adj_4865), .I1(n2612), .I2(n2570), 
            .I3(GND_net), .O(n2644));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1730_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_46_unary_minus_4_add_3_11 (.CI(n28785), .I0(GND_net), .I1(n16_adj_4902), 
            .CO(n28786));
    SB_LUT4 div_46_unary_minus_4_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_4903), .I3(n28784), .O(n67)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1222_add_4_33_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[31]), .I3(n28570), .O(n134)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_17 (.CI(n29001), .I0(n1944), .I1(VCC_net), 
            .CO(n29002));
    SB_CARRY div_46_unary_minus_4_add_3_10 (.CI(n28784), .I0(GND_net), .I1(n17_adj_4903), 
            .CO(n28785));
    SB_LUT4 communication_counter_1222_add_4_32_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[30]), .I3(n28569), .O(n135)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1729_3_lut (.I0(n2544_adj_4866), .I1(n2611), .I2(n2570), 
            .I3(GND_net), .O(n2643_adj_4843));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1729_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1222_add_4_32 (.CI(n28569), .I0(GND_net), 
            .I1(communication_counter[30]), .CO(n28570));
    SB_LUT4 communication_counter_1222_add_4_31_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[29]), .I3(n28568), .O(n136)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1222_add_4_31 (.CI(n28568), .I0(GND_net), 
            .I1(communication_counter[29]), .CO(n28569));
    SB_LUT4 communication_counter_1222_add_4_30_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[28]), .I3(n28567), .O(n137)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13195_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n4593), .I3(GND_net), .O(n17934));   // verilog/coms.v(127[12] 295[6])
    defparam i13195_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1222_add_4_30 (.CI(n28567), .I0(GND_net), 
            .I1(communication_counter[28]), .CO(n28568));
    SB_LUT4 communication_counter_1222_add_4_29_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[27]), .I3(n28566), .O(n138)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1222_add_4_29 (.CI(n28566), .I0(GND_net), 
            .I1(communication_counter[27]), .CO(n28567));
    SB_LUT4 rem_4_i1728_3_lut (.I0(n2543_adj_4867), .I1(n2610), .I2(n2570), 
            .I3(GND_net), .O(n2642_adj_4844));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1728_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13069_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position[16]), 
            .I2(n13302), .I3(GND_net), .O(n17808));   // verilog/coms.v(127[12] 295[6])
    defparam i13069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13070_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position[17]), 
            .I2(n13302), .I3(GND_net), .O(n17809));   // verilog/coms.v(127[12] 295[6])
    defparam i13070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1735_3_lut (.I0(n2550_adj_4860), .I1(n2617), .I2(n2570), 
            .I3(GND_net), .O(n2649));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1735_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13071_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position[18]), 
            .I2(n13302), .I3(GND_net), .O(n17810));   // verilog/coms.v(127[12] 295[6])
    defparam i13071_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13072_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position[19]), 
            .I2(n13302), .I3(GND_net), .O(n17811));   // verilog/coms.v(127[12] 295[6])
    defparam i13072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i23_1_lut (.I0(gearBoxRatio[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4889));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_4904), .I3(n28783), .O(n68)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1732_3_lut (.I0(n2547_adj_4863), .I1(n2614), .I2(n2570), 
            .I3(GND_net), .O(n2646));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_inv_0_i24_1_lut (.I0(gearBoxRatio[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n2_adj_4888));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 communication_counter_1222_add_4_28_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[26]), .I3(n28565), .O(n139)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1222_add_4_28 (.CI(n28565), .I0(GND_net), 
            .I1(communication_counter[26]), .CO(n28566));
    SB_LUT4 communication_counter_1222_add_4_27_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[25]), .I3(n28564), .O(n140)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_9 (.CI(n28783), .I0(GND_net), .I1(n18_adj_4904), 
            .CO(n28784));
    SB_CARRY communication_counter_1222_add_4_27 (.CI(n28564), .I0(GND_net), 
            .I1(communication_counter[25]), .CO(n28565));
    SB_LUT4 communication_counter_1222_add_4_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[24]), .I3(n28563), .O(n141)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13073_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position[20]), 
            .I2(n13302), .I3(GND_net), .O(n17812));   // verilog/coms.v(127[12] 295[6])
    defparam i13073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13074_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position[21]), 
            .I2(n13302), .I3(GND_net), .O(n17813));   // verilog/coms.v(127[12] 295[6])
    defparam i13074_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1222_add_4_26 (.CI(n28563), .I0(GND_net), 
            .I1(communication_counter[24]), .CO(n28564));
    SB_LUT4 div_46_unary_minus_4_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_4905), .I3(n28782), .O(n69)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_8 (.CI(n28782), .I0(GND_net), .I1(n19_adj_4905), 
            .CO(n28783));
    SB_LUT4 communication_counter_1222_add_4_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[23]), .I3(n28562), .O(n142)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1318_16_lut (.I0(GND_net), .I1(n1945), .I2(VCC_net), 
            .I3(n29000), .O(n2012)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1222_add_4_25 (.CI(n28562), .I0(GND_net), 
            .I1(communication_counter[23]), .CO(n28563));
    SB_LUT4 div_46_unary_minus_4_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_4906), .I3(n28781), .O(n70)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_16 (.CI(n29000), .I0(n1945), .I1(VCC_net), 
            .CO(n29001));
    SB_LUT4 i13075_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position[22]), 
            .I2(n13302), .I3(GND_net), .O(n17814));   // verilog/coms.v(127[12] 295[6])
    defparam i13075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13076_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position[23]), 
            .I2(n13302), .I3(GND_net), .O(n17815));   // verilog/coms.v(127[12] 295[6])
    defparam i13076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4935));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_1318_15_lut (.I0(GND_net), .I1(n1946), .I2(VCC_net), 
            .I3(n28999), .O(n2013)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_15 (.CI(n28999), .I0(n1946), .I1(VCC_net), 
            .CO(n29000));
    SB_LUT4 communication_counter_1222_add_4_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[22]), .I3(n28561), .O(n143)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13077_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position[8]), 
            .I2(n13302), .I3(GND_net), .O(n17816));   // verilog/coms.v(127[12] 295[6])
    defparam i13077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1318_14_lut (.I0(GND_net), .I1(n1947), .I2(VCC_net), 
            .I3(n28998), .O(n2014)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_7 (.CI(n28781), .I0(GND_net), .I1(n20_adj_4906), 
            .CO(n28782));
    SB_CARRY rem_4_add_1318_14 (.CI(n28998), .I0(n1947), .I1(VCC_net), 
            .CO(n28999));
    SB_LUT4 rem_4_add_1318_13_lut (.I0(GND_net), .I1(n1948), .I2(VCC_net), 
            .I3(n28997), .O(n2015)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_4_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_4907), .I3(n28780), .O(n71)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_6 (.CI(n28780), .I0(GND_net), .I1(n21_adj_4907), 
            .CO(n28781));
    SB_LUT4 div_46_unary_minus_4_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_4908), .I3(n28779), .O(n72)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1222_add_4_24 (.CI(n28561), .I0(GND_net), 
            .I1(communication_counter[22]), .CO(n28562));
    SB_LUT4 communication_counter_1222_add_4_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[21]), .I3(n28560), .O(n144)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13078_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position[9]), 
            .I2(n13302), .I3(GND_net), .O(n17817));   // verilog/coms.v(127[12] 295[6])
    defparam i13078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1192_3_lut (.I0(n1751), .I1(n1818), .I2(n1778_adj_4812), 
            .I3(GND_net), .O(n1850));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1192_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1222_add_4_23 (.CI(n28560), .I0(GND_net), 
            .I1(communication_counter[21]), .CO(n28561));
    SB_LUT4 rem_4_i653_3_lut (.I0(n956), .I1(n1023), .I2(n986), .I3(GND_net), 
            .O(n1055));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13079_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position[10]), 
            .I2(n13302), .I3(GND_net), .O(n17818));   // verilog/coms.v(127[12] 295[6])
    defparam i13079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1222_add_4_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[20]), .I3(n28559), .O(n145)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13080_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position[11]), 
            .I2(n13302), .I3(GND_net), .O(n17819));   // verilog/coms.v(127[12] 295[6])
    defparam i13080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1191_3_lut (.I0(n1750), .I1(n1817), .I2(n1778_adj_4812), 
            .I3(GND_net), .O(n1849));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1191_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1187_3_lut (.I0(n1746), .I1(n1813), .I2(n1778_adj_4812), 
            .I3(GND_net), .O(n1845));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1187_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13081_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position[12]), 
            .I2(n13302), .I3(GND_net), .O(n17820));   // verilog/coms.v(127[12] 295[6])
    defparam i13081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1737_3_lut (.I0(n2552_adj_4858), .I1(n2619_adj_4854), 
            .I2(n2570), .I3(GND_net), .O(n2651));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1737_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1731_3_lut (.I0(n2546_adj_4864), .I1(n2613), .I2(n2570), 
            .I3(GND_net), .O(n2645));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1731_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13082_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position[13]), 
            .I2(n13302), .I3(GND_net), .O(n17821));   // verilog/coms.v(127[12] 295[6])
    defparam i13082_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1318_13 (.CI(n28997), .I0(n1948), .I1(VCC_net), 
            .CO(n28998));
    SB_LUT4 rem_4_add_1318_12_lut (.I0(GND_net), .I1(n1949), .I2(VCC_net), 
            .I3(n28996), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13083_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position[14]), 
            .I2(n13302), .I3(GND_net), .O(n17822));   // verilog/coms.v(127[12] 295[6])
    defparam i13083_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_46_unary_minus_4_add_3_5 (.CI(n28779), .I0(GND_net), .I1(n22_adj_4908), 
            .CO(n28780));
    SB_CARRY communication_counter_1222_add_4_22 (.CI(n28559), .I0(GND_net), 
            .I1(communication_counter[20]), .CO(n28560));
    SB_LUT4 communication_counter_1222_add_4_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[19]), .I3(n28558), .O(n146)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1222_add_4_21 (.CI(n28558), .I0(GND_net), 
            .I1(communication_counter[19]), .CO(n28559));
    SB_LUT4 i13084_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position[15]), 
            .I2(n13302), .I3(GND_net), .O(n17823));   // verilog/coms.v(127[12] 295[6])
    defparam i13084_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1193_3_lut (.I0(n1752), .I1(n1819), .I2(n1778_adj_4812), 
            .I3(GND_net), .O(n1851));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1193_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1318_12 (.CI(n28996), .I0(n1949), .I1(VCC_net), 
            .CO(n28997));
    SB_LUT4 rem_4_i1190_3_lut (.I0(n1749), .I1(n1816), .I2(n1778_adj_4812), 
            .I3(GND_net), .O(n1848));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1190_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_4909), .I3(n28778), .O(n73)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13085_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position[0]), 
            .I2(n13302), .I3(GND_net), .O(n17824));   // verilog/coms.v(127[12] 295[6])
    defparam i13085_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1318_11_lut (.I0(GND_net), .I1(n1950), .I2(VCC_net), 
            .I3(n28995), .O(n2017)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_11 (.CI(n28995), .I0(n1950), .I1(VCC_net), 
            .CO(n28996));
    SB_LUT4 rem_4_i1733_3_lut (.I0(n2548_adj_4862), .I1(n2615), .I2(n2570), 
            .I3(GND_net), .O(n2647));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1733_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1318_10_lut (.I0(GND_net), .I1(n1951), .I2(VCC_net), 
            .I3(n28994), .O(n2018)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_4_add_3_4 (.CI(n28778), .I0(GND_net), .I1(n23_adj_4909), 
            .CO(n28779));
    SB_LUT4 i13086_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position[1]), 
            .I2(n13302), .I3(GND_net), .O(n17825));   // verilog/coms.v(127[12] 295[6])
    defparam i13086_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_4910), .I3(n28777), .O(n74)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1189_3_lut (.I0(n1748), .I1(n1815), .I2(n1778_adj_4812), 
            .I3(GND_net), .O(n1847));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1188_3_lut (.I0(n1747), .I1(n1814), .I2(n1778_adj_4812), 
            .I3(GND_net), .O(n1846));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1188_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1318_10 (.CI(n28994), .I0(n1951), .I1(VCC_net), 
            .CO(n28995));
    SB_CARRY div_46_unary_minus_4_add_3_3 (.CI(n28777), .I0(GND_net), .I1(n24_adj_4910), 
            .CO(n28778));
    SB_LUT4 rem_4_i1734_rep_42_3_lut (.I0(n2549_adj_4861), .I1(n2616), .I2(n2570), 
            .I3(GND_net), .O(n2648));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1734_rep_42_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13087_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position[2]), 
            .I2(n13302), .I3(GND_net), .O(n17826));   // verilog/coms.v(127[12] 295[6])
    defparam i13087_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1194_3_lut (.I0(n1753), .I1(n1820), .I2(n1778_adj_4812), 
            .I3(GND_net), .O(n1852));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1738_3_lut (.I0(n2553_adj_4857), .I1(n2620_adj_4853), 
            .I2(n2570), .I3(GND_net), .O(n2652));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1738_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_4_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_4911), .I3(VCC_net), .O(n75)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_4_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1318_9_lut (.I0(GND_net), .I1(n1952), .I2(VCC_net), 
            .I3(n28993), .O(n2019)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13088_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position[3]), 
            .I2(n13302), .I3(GND_net), .O(n17827));   // verilog/coms.v(127[12] 295[6])
    defparam i13088_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1318_9 (.CI(n28993), .I0(n1952), .I1(VCC_net), 
            .CO(n28994));
    SB_LUT4 i13089_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position[4]), 
            .I2(n13302), .I3(GND_net), .O(n17828));   // verilog/coms.v(127[12] 295[6])
    defparam i13089_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY div_46_unary_minus_4_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n25_adj_4911), 
            .CO(n28777));
    SB_LUT4 rem_4_i1195_3_lut (.I0(n1754_adj_4807), .I1(n1821), .I2(n1778_adj_4812), 
            .I3(GND_net), .O(n1853));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1199_3_lut (.I0(n1758_adj_4811), .I1(n1825), .I2(n1778_adj_4812), 
            .I3(GND_net), .O(n1857));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13090_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position[5]), 
            .I2(n13302), .I3(GND_net), .O(n17829));   // verilog/coms.v(127[12] 295[6])
    defparam i13090_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13091_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position[6]), 
            .I2(n13302), .I3(GND_net), .O(n17830));   // verilog/coms.v(127[12] 295[6])
    defparam i13091_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13092_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position[7]), 
            .I2(n13302), .I3(GND_net), .O(n17831));   // verilog/coms.v(127[12] 295[6])
    defparam i13092_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13093_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position[16]), 
            .I2(n13302), .I3(GND_net), .O(n17832));   // verilog/coms.v(127[12] 295[6])
    defparam i13093_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1921_27_lut (.I0(n2867), .I1(n2834), .I2(VCC_net), 
            .I3(n28776), .O(n2933)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_i1197_3_lut (.I0(n1756_adj_4809), .I1(n1823), .I2(n1778_adj_4812), 
            .I3(GND_net), .O(n1855));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1196_3_lut (.I0(n1755_adj_4808), .I1(n1822), .I2(n1778_adj_4812), 
            .I3(GND_net), .O(n1854));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1198_3_lut (.I0(n1757_adj_4810), .I1(n1824), .I2(n1778_adj_4812), 
            .I3(GND_net), .O(n1856));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1318_8_lut (.I0(GND_net), .I1(n1953), .I2(VCC_net), 
            .I3(n28992), .O(n2020)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13094_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position[17]), 
            .I2(n13302), .I3(GND_net), .O(n17833));   // verilog/coms.v(127[12] 295[6])
    defparam i13094_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(n1856), .I1(n1858), .I2(GND_net), .I3(GND_net), 
            .O(n38277));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 rem_4_add_1921_26_lut (.I0(GND_net), .I1(n2835), .I2(VCC_net), 
            .I3(n28775), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1725 (.I0(n1854), .I1(n38277), .I2(n1855), .I3(n1857), 
            .O(n36006));
    defparam i1_4_lut_adj_1725.LUT_INIT = 16'ha080;
    SB_CARRY rem_4_add_1921_26 (.CI(n28775), .I0(n2835), .I1(VCC_net), 
            .CO(n28776));
    SB_LUT4 rem_4_i652_3_lut (.I0(n955), .I1(n1022), .I2(n986), .I3(GND_net), 
            .O(n1054));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i652_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1318_8 (.CI(n28992), .I0(n1953), .I1(VCC_net), 
            .CO(n28993));
    SB_LUT4 rem_4_add_1318_7_lut (.I0(GND_net), .I1(n1954), .I2(GND_net), 
            .I3(n28991), .O(n2021)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_25_lut (.I0(GND_net), .I1(n2836), .I2(VCC_net), 
            .I3(n28774), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_25 (.CI(n28774), .I0(n2836), .I1(VCC_net), 
            .CO(n28775));
    SB_CARRY rem_4_add_1318_7 (.CI(n28991), .I0(n1954), .I1(GND_net), 
            .CO(n28992));
    SB_LUT4 i13095_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position[18]), 
            .I2(n13302), .I3(GND_net), .O(n17834));   // verilog/coms.v(127[12] 295[6])
    defparam i13095_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1222_add_4_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[18]), .I3(n28557), .O(n147)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1222_add_4_20 (.CI(n28557), .I0(GND_net), 
            .I1(communication_counter[18]), .CO(n28558));
    SB_LUT4 rem_4_add_1921_24_lut (.I0(GND_net), .I1(n2837), .I2(VCC_net), 
            .I3(n28773), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1318_6_lut (.I0(GND_net), .I1(n1955), .I2(GND_net), 
            .I3(n28990), .O(n2022)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_24 (.CI(n28773), .I0(n2837), .I1(VCC_net), 
            .CO(n28774));
    SB_LUT4 rem_4_add_1921_23_lut (.I0(GND_net), .I1(n2838), .I2(VCC_net), 
            .I3(n28772), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_6 (.CI(n28990), .I0(n1955), .I1(GND_net), 
            .CO(n28991));
    SB_LUT4 i13096_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position[19]), 
            .I2(n13302), .I3(GND_net), .O(n17835));   // verilog/coms.v(127[12] 295[6])
    defparam i13096_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13097_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position[20]), 
            .I2(n13302), .I3(GND_net), .O(n17836));   // verilog/coms.v(127[12] 295[6])
    defparam i13097_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i26_3_lut (.I0(communication_counter[25]), .I1(n8_adj_4801), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1058));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1736_3_lut (.I0(n2551_adj_4859), .I1(n2618_adj_4855), 
            .I2(n2570), .I3(GND_net), .O(n2650));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1736_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_23 (.CI(n28772), .I0(n2838), .I1(VCC_net), 
            .CO(n28773));
    SB_LUT4 i13098_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position[21]), 
            .I2(n13302), .I3(GND_net), .O(n17837));   // verilog/coms.v(127[12] 295[6])
    defparam i13098_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1921_22_lut (.I0(GND_net), .I1(n2839), .I2(VCC_net), 
            .I3(n28771), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1222_add_4_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[17]), .I3(n28556), .O(n148)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1222_add_4_19 (.CI(n28556), .I0(GND_net), 
            .I1(communication_counter[17]), .CO(n28557));
    SB_LUT4 rem_4_add_1318_5_lut (.I0(GND_net), .I1(n1956), .I2(VCC_net), 
            .I3(n28989), .O(n2023)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1222_add_4_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[16]), .I3(n28555), .O(n149)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1723_3_lut (.I0(n2538_adj_4872), .I1(n2605), .I2(n2570), 
            .I3(GND_net), .O(n2637_adj_4846));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1739_rep_40_3_lut (.I0(n2554), .I1(n2621_adj_4852), .I2(n2570), 
            .I3(GND_net), .O(n2653));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1739_rep_40_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut_adj_1726 (.I0(n1846), .I1(n36006), .I2(n1847), .I3(n1848), 
            .O(n18));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i7_4_lut_adj_1726.LUT_INIT = 16'hfffe;
    SB_LUT4 i13099_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position[22]), 
            .I2(n13302), .I3(GND_net), .O(n17838));   // verilog/coms.v(127[12] 295[6])
    defparam i13099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_2_lut (.I0(n1853), .I1(n1852), .I2(GND_net), .I3(GND_net), 
            .O(n16));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY rem_4_add_1921_22 (.CI(n28771), .I0(n2839), .I1(VCC_net), 
            .CO(n28772));
    SB_CARRY rem_4_add_1318_5 (.CI(n28989), .I0(n1956), .I1(VCC_net), 
            .CO(n28990));
    SB_CARRY communication_counter_1222_add_4_18 (.CI(n28555), .I0(GND_net), 
            .I1(communication_counter[16]), .CO(n28556));
    SB_LUT4 rem_4_add_1921_21_lut (.I0(GND_net), .I1(n2840), .I2(VCC_net), 
            .I3(n28770), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1222_add_4_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[15]), .I3(n28554), .O(n150)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1222_add_4_17 (.CI(n28554), .I0(GND_net), 
            .I1(communication_counter[15]), .CO(n28555));
    SB_CARRY rem_4_add_1921_21 (.CI(n28770), .I0(n2840), .I1(VCC_net), 
            .CO(n28771));
    SB_LUT4 rem_4_add_1318_4_lut (.I0(GND_net), .I1(n1957), .I2(VCC_net), 
            .I3(n28988), .O(n2024)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1222_add_4_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[14]), .I3(n28553), .O(n151)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1318_4 (.CI(n28988), .I0(n1957), .I1(VCC_net), 
            .CO(n28989));
    SB_LUT4 rem_4_i1743_3_lut (.I0(n2558_adj_4856), .I1(n2625_adj_4848), 
            .I2(n2570), .I3(GND_net), .O(n2657));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1743_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1222_add_4_16 (.CI(n28553), .I0(GND_net), 
            .I1(communication_counter[14]), .CO(n28554));
    SB_LUT4 communication_counter_1222_add_4_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[13]), .I3(n28552), .O(n152)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1318_3_lut (.I0(GND_net), .I1(n1958), .I2(GND_net), 
            .I3(n28987), .O(n2025)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1318_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_20_lut (.I0(GND_net), .I1(n2841), .I2(VCC_net), 
            .I3(n28769), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_20 (.CI(n28769), .I0(n2841), .I1(VCC_net), 
            .CO(n28770));
    SB_CARRY rem_4_add_1318_3 (.CI(n28987), .I0(n1958), .I1(GND_net), 
            .CO(n28988));
    SB_LUT4 rem_4_add_1921_19_lut (.I0(GND_net), .I1(n2842), .I2(VCC_net), 
            .I3(n28768), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13100_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position[23]), 
            .I2(n13302), .I3(GND_net), .O(n17839));   // verilog/coms.v(127[12] 295[6])
    defparam i13100_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_4_lut (.I0(n1851), .I1(n18), .I2(n1845), .I3(n1844), 
            .O(n20));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY communication_counter_1222_add_4_15 (.CI(n28552), .I0(GND_net), 
            .I1(communication_counter[13]), .CO(n28553));
    SB_LUT4 communication_counter_1222_add_4_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[12]), .I3(n28551), .O(n153)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_19 (.CI(n28768), .I0(n2842), .I1(VCC_net), 
            .CO(n28769));
    SB_CARRY rem_4_add_1318_2 (.CI(VCC_net), .I0(n2058), .I1(VCC_net), 
            .CO(n28987));
    SB_LUT4 i13101_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position[8]), 
            .I2(n13302), .I3(GND_net), .O(n17840));   // verilog/coms.v(127[12] 295[6])
    defparam i13101_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1385_19_lut (.I0(n2075_adj_5028), .I1(n2042), .I2(VCC_net), 
            .I3(n28986), .O(n2141)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1921_18_lut (.I0(GND_net), .I1(n2843), .I2(VCC_net), 
            .I3(n28767), .O(n2910)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13102_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position[9]), 
            .I2(n13302), .I3(GND_net), .O(n17841));   // verilog/coms.v(127[12] 295[6])
    defparam i13102_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10_4_lut_adj_1727 (.I0(n1849), .I1(n20), .I2(n16), .I3(n1850), 
            .O(n1877));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i10_4_lut_adj_1727.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1921_18 (.CI(n28767), .I0(n2843), .I1(VCC_net), 
            .CO(n28768));
    SB_LUT4 rem_4_add_1921_17_lut (.I0(GND_net), .I1(n2844), .I2(VCC_net), 
            .I3(n28766), .O(n2911)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13103_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position[10]), 
            .I2(n13302), .I3(GND_net), .O(n17842));   // verilog/coms.v(127[12] 295[6])
    defparam i13103_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13104_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position[11]), 
            .I2(n13302), .I3(GND_net), .O(n17843));   // verilog/coms.v(127[12] 295[6])
    defparam i13104_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1222_add_4_14 (.CI(n28551), .I0(GND_net), 
            .I1(communication_counter[12]), .CO(n28552));
    SB_LUT4 rem_4_mux_3_i18_3_lut (.I0(communication_counter[17]), .I1(n16_adj_4793), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1858));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1222_add_4_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[11]), .I3(n28550), .O(n154)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13105_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position[12]), 
            .I2(n13302), .I3(GND_net), .O(n17844));   // verilog/coms.v(127[12] 295[6])
    defparam i13105_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1385_18_lut (.I0(GND_net), .I1(n2043), .I2(VCC_net), 
            .I3(n28985), .O(n2110)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1222_add_4_13 (.CI(n28550), .I0(GND_net), 
            .I1(communication_counter[11]), .CO(n28551));
    SB_LUT4 communication_counter_1222_add_4_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[10]), .I3(n28549), .O(n155)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13106_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position[13]), 
            .I2(n13302), .I3(GND_net), .O(n17845));   // verilog/coms.v(127[12] 295[6])
    defparam i13106_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1741_3_lut (.I0(n2556), .I1(n2623_adj_4850), .I2(n2570), 
            .I3(GND_net), .O(n2655));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1741_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF h1_55 (.Q(PIN_20_c), .C(clk32MHz), .D(hall1));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_LUT4 i13107_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position[14]), 
            .I2(n13302), .I3(GND_net), .O(n17846));   // verilog/coms.v(127[12] 295[6])
    defparam i13107_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1222_add_4_12 (.CI(n28549), .I0(GND_net), 
            .I1(communication_counter[10]), .CO(n28550));
    SB_CARRY rem_4_add_1921_17 (.CI(n28766), .I0(n2844), .I1(VCC_net), 
            .CO(n28767));
    SB_LUT4 communication_counter_1222_add_4_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[9]), .I3(n28548), .O(n156)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_18 (.CI(n28985), .I0(n2043), .I1(VCC_net), 
            .CO(n28986));
    SB_CARRY communication_counter_1222_add_4_11 (.CI(n28548), .I0(GND_net), 
            .I1(communication_counter[9]), .CO(n28549));
    SB_LUT4 i13108_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position[15]), 
            .I2(n13302), .I3(GND_net), .O(n17847));   // verilog/coms.v(127[12] 295[6])
    defparam i13108_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1921_16_lut (.I0(GND_net), .I1(n2845), .I2(VCC_net), 
            .I3(n28765), .O(n2912)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_16 (.CI(n28765), .I0(n2845), .I1(VCC_net), 
            .CO(n28766));
    SB_LUT4 rem_4_add_1921_15_lut (.I0(GND_net), .I1(n2846), .I2(VCC_net), 
            .I3(n28764), .O(n2913)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_17_lut (.I0(GND_net), .I1(n2044), .I2(VCC_net), 
            .I3(n28984), .O(n2111)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1222_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[8]), .I3(n28547), .O(n157)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1222_add_4_10 (.CI(n28547), .I0(GND_net), 
            .I1(communication_counter[8]), .CO(n28548));
    SB_LUT4 i13109_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position[0]), 
            .I2(n13302), .I3(GND_net), .O(n17848));   // verilog/coms.v(127[12] 295[6])
    defparam i13109_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13110_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position[1]), 
            .I2(n13302), .I3(GND_net), .O(n17849));   // verilog/coms.v(127[12] 295[6])
    defparam i13110_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_15 (.CI(n28764), .I0(n2846), .I1(VCC_net), 
            .CO(n28765));
    SB_LUT4 communication_counter_1222_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[7]), .I3(n28546), .O(n158)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1222_add_4_9 (.CI(n28546), .I0(GND_net), 
            .I1(communication_counter[7]), .CO(n28547));
    SB_LUT4 i13111_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position[2]), 
            .I2(n13302), .I3(GND_net), .O(n17850));   // verilog/coms.v(127[12] 295[6])
    defparam i13111_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1385_17 (.CI(n28984), .I0(n2044), .I1(VCC_net), 
            .CO(n28985));
    SB_LUT4 i13112_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position[3]), 
            .I2(n13302), .I3(GND_net), .O(n17851));   // verilog/coms.v(127[12] 295[6])
    defparam i13112_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1385_16_lut (.I0(GND_net), .I1(n2045), .I2(VCC_net), 
            .I3(n28983), .O(n2112)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1740_3_lut (.I0(n2555), .I1(n2622_adj_4851), .I2(n2570), 
            .I3(GND_net), .O(n2654));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1740_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1921_14_lut (.I0(GND_net), .I1(n2847), .I2(VCC_net), 
            .I3(n28763), .O(n2914)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i654_3_lut (.I0(n957), .I1(n1024), .I2(n986), .I3(GND_net), 
            .O(n1056));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1742_3_lut (.I0(n2557), .I1(n2624_adj_4849), .I2(n2570), 
            .I3(GND_net), .O(n2656));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1742_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1385_16 (.CI(n28983), .I0(n2045), .I1(VCC_net), 
            .CO(n28984));
    SB_LUT4 communication_counter_1222_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[6]), .I3(n28545), .O(n159)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13113_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position[4]), 
            .I2(n13302), .I3(GND_net), .O(n17852));   // verilog/coms.v(127[12] 295[6])
    defparam i13113_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13114_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position[5]), 
            .I2(n13302), .I3(GND_net), .O(n17853));   // verilog/coms.v(127[12] 295[6])
    defparam i13114_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13115_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position[6]), 
            .I2(n13302), .I3(GND_net), .O(n17854));   // verilog/coms.v(127[12] 295[6])
    defparam i13115_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13116_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position[7]), 
            .I2(n13302), .I3(GND_net), .O(n17855));   // verilog/coms.v(127[12] 295[6])
    defparam i13116_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13117_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n13302), .I3(GND_net), .O(n17856));   // verilog/coms.v(127[12] 295[6])
    defparam i13117_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_14 (.CI(n28763), .I0(n2847), .I1(VCC_net), 
            .CO(n28764));
    SB_CARRY communication_counter_1222_add_4_8 (.CI(n28545), .I0(GND_net), 
            .I1(communication_counter[6]), .CO(n28546));
    SB_LUT4 rem_4_i1662_3_lut (.I0(n2445), .I1(n2512), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2544_adj_4866));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1385_15_lut (.I0(GND_net), .I1(n2046), .I2(VCC_net), 
            .I3(n28982), .O(n2113)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13118_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n13302), .I3(GND_net), .O(n17857));   // verilog/coms.v(127[12] 295[6])
    defparam i13118_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1921_13_lut (.I0(GND_net), .I1(n2848), .I2(VCC_net), 
            .I3(n28762), .O(n2915)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_15 (.CI(n28982), .I0(n2046), .I1(VCC_net), 
            .CO(n28983));
    SB_LUT4 i13119_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n13302), .I3(GND_net), .O(n17858));   // verilog/coms.v(127[12] 295[6])
    defparam i13119_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_13 (.CI(n28762), .I0(n2848), .I1(VCC_net), 
            .CO(n28763));
    SB_LUT4 communication_counter_1222_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[5]), .I3(n28544), .O(n160)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1222_add_4_7 (.CI(n28544), .I0(GND_net), 
            .I1(communication_counter[5]), .CO(n28545));
    SB_LUT4 i13120_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n13302), .I3(GND_net), .O(n17859));   // verilog/coms.v(127[12] 295[6])
    defparam i13120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1222_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[4]), .I3(n28543), .O(n161)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_20_pad (.PACKAGE_PIN(PIN_20), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_20_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_20_pad.PIN_TYPE = 6'b011001;
    defparam PIN_20_pad.PULLUP = 1'b0;
    defparam PIN_20_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_20_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_19_pad (.PACKAGE_PIN(PIN_19), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_19_c_0)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_19_pad.PIN_TYPE = 6'b011001;
    defparam PIN_19_pad.PULLUP = 1'b0;
    defparam PIN_19_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_19_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 rem_4_add_1385_14_lut (.I0(GND_net), .I1(n2047), .I2(VCC_net), 
            .I3(n28981), .O(n2114)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_12_lut (.I0(GND_net), .I1(n2849), .I2(VCC_net), 
            .I3(n28761), .O(n2916)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_14 (.CI(n28981), .I0(n2047), .I1(VCC_net), 
            .CO(n28982));
    SB_CARRY communication_counter_1222_add_4_6 (.CI(n28543), .I0(GND_net), 
            .I1(communication_counter[4]), .CO(n28544));
    SB_CARRY rem_4_add_1921_12 (.CI(n28761), .I0(n2849), .I1(VCC_net), 
            .CO(n28762));
    SB_LUT4 rem_4_add_1385_13_lut (.I0(GND_net), .I1(n2048), .I2(VCC_net), 
            .I3(n28980), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_11_lut (.I0(GND_net), .I1(n2850), .I2(VCC_net), 
            .I3(n28760), .O(n2917)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1222_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[3]), .I3(n28542), .O(n162)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_11 (.CI(n28760), .I0(n2850), .I1(VCC_net), 
            .CO(n28761));
    SB_CARRY rem_4_add_1385_13 (.CI(n28980), .I0(n2048), .I1(VCC_net), 
            .CO(n28981));
    SB_LUT4 i13121_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n13302), .I3(GND_net), .O(n17860));   // verilog/coms.v(127[12] 295[6])
    defparam i13121_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY communication_counter_1222_add_4_5 (.CI(n28542), .I0(GND_net), 
            .I1(communication_counter[3]), .CO(n28543));
    SB_LUT4 rem_4_add_1385_12_lut (.I0(GND_net), .I1(n2049), .I2(VCC_net), 
            .I3(n28979), .O(n2116)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1661_3_lut (.I0(n2444), .I1(n2511), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2543_adj_4867));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1921_10_lut (.I0(GND_net), .I1(n2851), .I2(VCC_net), 
            .I3(n28759), .O(n2918)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_12 (.CI(n28979), .I0(n2049), .I1(VCC_net), 
            .CO(n28980));
    SB_LUT4 rem_4_i1659_3_lut (.I0(n2442), .I1(n2509), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2541_adj_4869));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1667_3_lut (.I0(n2450_adj_4884), .I1(n2517), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2549_adj_4861));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13122_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n13302), .I3(GND_net), .O(n17861));   // verilog/coms.v(127[12] 295[6])
    defparam i13122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13123_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n13302), .I3(GND_net), .O(n17862));   // verilog/coms.v(127[12] 295[6])
    defparam i13123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13124_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n13302), .I3(GND_net), .O(n17863));   // verilog/coms.v(127[12] 295[6])
    defparam i13124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1385_11_lut (.I0(GND_net), .I1(n2050), .I2(VCC_net), 
            .I3(n28978), .O(n2117)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 communication_counter_1222_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[2]), .I3(n28541), .O(n163)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_10 (.CI(n28759), .I0(n2851), .I1(VCC_net), 
            .CO(n28760));
    SB_CARRY communication_counter_1222_add_4_4 (.CI(n28541), .I0(GND_net), 
            .I1(communication_counter[2]), .CO(n28542));
    SB_LUT4 communication_counter_1222_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[1]), .I3(n28540), .O(n164)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_11 (.CI(n28978), .I0(n2050), .I1(VCC_net), 
            .CO(n28979));
    SB_LUT4 rem_4_add_1921_9_lut (.I0(GND_net), .I1(n2852), .I2(VCC_net), 
            .I3(n28758), .O(n2919)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1222_add_4_3 (.CI(n28540), .I0(GND_net), 
            .I1(communication_counter[1]), .CO(n28541));
    SB_LUT4 i13125_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n13302), .I3(GND_net), .O(n17864));   // verilog/coms.v(127[12] 295[6])
    defparam i13125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 communication_counter_1222_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(communication_counter[0]), .I3(VCC_net), .O(n165)) /* synthesis syn_instantiated=1 */ ;
    defparam communication_counter_1222_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY communication_counter_1222_add_4_2 (.CI(VCC_net), .I0(GND_net), 
            .I1(communication_counter[0]), .CO(n28540));
    SB_LUT4 add_5571_7_lut (.I0(GND_net), .I1(n3353), .I2(VCC_net), .I3(n28539), 
            .O(n10244)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5571_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5571_6_lut (.I0(GND_net), .I1(n3354), .I2(GND_net), .I3(n28538), 
            .O(n10245)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5571_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5571_6 (.CI(n28538), .I0(n3354), .I1(GND_net), .CO(n28539));
    SB_LUT4 i13126_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n13302), .I3(GND_net), .O(n17865));   // verilog/coms.v(127[12] 295[6])
    defparam i13126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5571_5_lut (.I0(GND_net), .I1(n3355), .I2(GND_net), .I3(n28537), 
            .O(n10246)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5571_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5571_5 (.CI(n28537), .I0(n3355), .I1(GND_net), .CO(n28538));
    SB_LUT4 add_5571_4_lut (.I0(GND_net), .I1(n3356), .I2(VCC_net), .I3(n28536), 
            .O(n10247)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5571_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1663_3_lut (.I0(n2446), .I1(n2513), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2545_adj_4865));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1663_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_9 (.CI(n28758), .I0(n2852), .I1(VCC_net), 
            .CO(n28759));
    SB_CARRY add_5571_4 (.CI(n28536), .I0(n3356), .I1(VCC_net), .CO(n28537));
    SB_LUT4 rem_4_add_1921_8_lut (.I0(GND_net), .I1(n2853), .I2(VCC_net), 
            .I3(n28757), .O(n2920)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5571_3_lut (.I0(GND_net), .I1(n3357), .I2(VCC_net), .I3(n28535), 
            .O(n10248)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5571_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5571_3 (.CI(n28535), .I0(n3357), .I1(VCC_net), .CO(n28536));
    SB_LUT4 i13127_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n13302), .I3(GND_net), .O(n17866));   // verilog/coms.v(127[12] 295[6])
    defparam i13127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1385_10_lut (.I0(GND_net), .I1(n2051), .I2(VCC_net), 
            .I3(n28977), .O(n2118)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_8 (.CI(n28757), .I0(n2853), .I1(VCC_net), 
            .CO(n28758));
    SB_LUT4 i13128_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n13302), .I3(GND_net), .O(n17867));   // verilog/coms.v(127[12] 295[6])
    defparam i13128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5571_2_lut (.I0(GND_net), .I1(n3358), .I2(GND_net), .I3(VCC_net), 
            .O(n10249)) /* synthesis syn_instantiated=1 */ ;
    defparam add_5571_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5571_2 (.CI(VCC_net), .I0(n3358), .I1(GND_net), .CO(n28535));
    SB_LUT4 i13129_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n13302), .I3(GND_net), .O(n17868));   // verilog/coms.v(127[12] 295[6])
    defparam i13129_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1385_10 (.CI(n28977), .I0(n2051), .I1(VCC_net), 
            .CO(n28978));
    SB_LUT4 rem_4_add_1385_9_lut (.I0(GND_net), .I1(n2052), .I2(VCC_net), 
            .I3(n28976), .O(n2119)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1921_7_lut (.I0(GND_net), .I1(n2854), .I2(GND_net), 
            .I3(n28756), .O(n2921)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13130_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n13302), .I3(GND_net), .O(n17869));   // verilog/coms.v(127[12] 295[6])
    defparam i13130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13131_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n13302), .I3(GND_net), .O(n17870));   // verilog/coms.v(127[12] 295[6])
    defparam i13131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1664_3_lut (.I0(n2447_adj_4887), .I1(n2514), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2546_adj_4864));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1671_3_lut (.I0(n2454_adj_4879), .I1(n2521), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2553_adj_4857));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2357_25_lut (.I0(n249), .I1(n43635), .I2(n248), .I3(n28534), 
            .O(displacement_23__N_229[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_25_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1385_9 (.CI(n28976), .I0(n2052), .I1(VCC_net), 
            .CO(n28977));
    SB_CARRY rem_4_add_1921_7 (.CI(n28756), .I0(n2854), .I1(GND_net), 
            .CO(n28757));
    SB_LUT4 rem_4_add_1385_8_lut (.I0(GND_net), .I1(n2053), .I2(VCC_net), 
            .I3(n28975), .O(n2120)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2357_24_lut (.I0(n393), .I1(n43635), .I2(n392), .I3(n28533), 
            .O(displacement_23__N_229[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1921_6_lut (.I0(GND_net), .I1(n2855), .I2(GND_net), 
            .I3(n28755), .O(n2922)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_8 (.CI(n28975), .I0(n2053), .I1(VCC_net), 
            .CO(n28976));
    SB_CARRY add_2357_24 (.CI(n28533), .I0(n43635), .I1(n392), .CO(n28534));
    SB_CARRY rem_4_add_1921_6 (.CI(n28755), .I0(n2855), .I1(GND_net), 
            .CO(n28756));
    SB_DFF communication_counter_1222__i0 (.Q(communication_counter[0]), .C(LED_c), 
           .D(n165));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_LUT4 add_2357_23_lut (.I0(n534), .I1(n43635), .I2(n533), .I3(n28532), 
            .O(displacement_23__N_229[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_23_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1385_7_lut (.I0(GND_net), .I1(n2054), .I2(GND_net), 
            .I3(n28974), .O(n2121)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_7 (.CI(n28974), .I0(n2054), .I1(GND_net), 
            .CO(n28975));
    SB_LUT4 rem_4_add_1921_5_lut (.I0(GND_net), .I1(n2856), .I2(VCC_net), 
            .I3(n28754), .O(n2923)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1385_6_lut (.I0(GND_net), .I1(n2055), .I2(GND_net), 
            .I3(n28973), .O(n2122)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_6 (.CI(n28973), .I0(n2055), .I1(GND_net), 
            .CO(n28974));
    SB_CARRY rem_4_add_1921_5 (.CI(n28754), .I0(n2856), .I1(VCC_net), 
            .CO(n28755));
    SB_LUT4 rem_4_add_1385_5_lut (.I0(GND_net), .I1(n2056), .I2(VCC_net), 
            .I3(n28972), .O(n2123)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_5 (.CI(n28972), .I0(n2056), .I1(VCC_net), 
            .CO(n28973));
    SB_LUT4 rem_4_add_1921_4_lut (.I0(GND_net), .I1(n2857), .I2(VCC_net), 
            .I3(n28753), .O(n2924)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_4 (.CI(n28753), .I0(n2857), .I1(VCC_net), 
            .CO(n28754));
    SB_LUT4 rem_4_add_1921_3_lut (.I0(GND_net), .I1(n2858), .I2(GND_net), 
            .I3(n28752), .O(n2925)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1921_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13132_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n13302), .I3(GND_net), .O(n17871));   // verilog/coms.v(127[12] 295[6])
    defparam i13132_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2357_23 (.CI(n28532), .I0(n43635), .I1(n533), .CO(n28533));
    SB_LUT4 i13133_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n13302), .I3(GND_net), .O(n17872));   // verilog/coms.v(127[12] 295[6])
    defparam i13133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1668_3_lut (.I0(n2451_adj_4883), .I1(n2518), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2550_adj_4860));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1385_4_lut (.I0(GND_net), .I1(n2057), .I2(VCC_net), 
            .I3(n28971), .O(n2124)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1921_3 (.CI(n28752), .I0(n2858), .I1(GND_net), 
            .CO(n28753));
    SB_CARRY rem_4_add_1385_4 (.CI(n28971), .I0(n2057), .I1(VCC_net), 
            .CO(n28972));
    SB_LUT4 i13134_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n13302), .I3(GND_net), .O(n17873));   // verilog/coms.v(127[12] 295[6])
    defparam i13134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13135_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n13302), .I3(GND_net), .O(n17874));   // verilog/coms.v(127[12] 295[6])
    defparam i13135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13136_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n13302), .I3(GND_net), .O(n17875));   // verilog/coms.v(127[12] 295[6])
    defparam i13136_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1921_2 (.CI(VCC_net), .I0(n2958_adj_4764), .I1(VCC_net), 
            .CO(n28752));
    SB_LUT4 rem_4_i1669_3_lut (.I0(n2452_adj_4882), .I1(n2519), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2551_adj_4859));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13137_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n13302), .I3(GND_net), .O(n17876));   // verilog/coms.v(127[12] 295[6])
    defparam i13137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13138_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n13302), .I3(GND_net), .O(n17877));   // verilog/coms.v(127[12] 295[6])
    defparam i13138_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1670_3_lut (.I0(n2453_adj_4881), .I1(n2520), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2552_adj_4858));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13139_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n13302), .I3(GND_net), .O(n17878));   // verilog/coms.v(127[12] 295[6])
    defparam i13139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1665_3_lut (.I0(n2448_adj_4886), .I1(n2515), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2547_adj_4863));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1666_3_lut (.I0(n2449_adj_4885), .I1(n2516), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2548_adj_4862));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2357_22_lut (.I0(n672), .I1(n43635), .I2(n671), .I3(n28531), 
            .O(displacement_23__N_229[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_i1675_3_lut (.I0(n2458_adj_4875), .I1(n2525), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2557));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1385_3_lut (.I0(GND_net), .I1(n2058), .I2(GND_net), 
            .I3(n28970), .O(n2125)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1385_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1385_3 (.CI(n28970), .I0(n2058), .I1(GND_net), 
            .CO(n28971));
    SB_LUT4 rem_4_add_1988_28_lut (.I0(n2966_adj_4763), .I1(n2933), .I2(VCC_net), 
            .I3(n28751), .O(n3032)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_i1673_3_lut (.I0(n2456_adj_4877), .I1(n2523), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2555));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13140_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n13302), .I3(GND_net), .O(n17879));   // verilog/coms.v(127[12] 295[6])
    defparam i13140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13141_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n13302), 
            .I3(GND_net), .O(n17880));   // verilog/coms.v(127[12] 295[6])
    defparam i13141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i41_4_lut (.I0(n2702), .I1(n80), .I2(n6220), 
            .I3(n2724), .O(n41_adj_5224));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i41_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 rem_4_i1672_3_lut (.I0(n2455_adj_4878), .I1(n2522), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2554));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i39_4_lut (.I0(n2703), .I1(n81), .I2(n6221), 
            .I3(n2724), .O(n39_adj_5223));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i39_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_mux_3_i1_3_lut (.I0(encoder0_position[0]), .I1(n25_adj_4711), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n1066));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i11_3_lut (.I0(communication_counter[10]), .I1(n23_adj_4786), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2558_adj_4856));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i45_4_lut (.I0(n2700), .I1(n78), .I2(n6218), 
            .I3(n2724), .O(n45_adj_5226));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i45_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i43_4_lut (.I0(n2701), .I1(n79), .I2(n6219), 
            .I3(n2724), .O(n43_adj_5225));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i43_4_lut.LUT_INIT = 16'hc399;
    SB_CARRY rem_4_add_1385_2 (.CI(VCC_net), .I0(n2158), .I1(VCC_net), 
            .CO(n28970));
    SB_LUT4 rem_4_add_1988_27_lut (.I0(GND_net), .I1(n2934), .I2(VCC_net), 
            .I3(n28750), .O(n3001_adj_4762)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_20_lut (.I0(n2174_adj_4984), .I1(n2141), .I2(VCC_net), 
            .I3(n28969), .O(n2240)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_46_LessThan_1830_i29_4_lut (.I0(n2708), .I1(n86), .I2(n6226), 
            .I3(n2724), .O(n29_adj_5217));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i29_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 rem_4_i1674_3_lut (.I0(n2457_adj_4876), .I1(n2524), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2556));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i31_4_lut (.I0(n2707), .I1(n85), .I2(n6225), 
            .I3(n2724), .O(n31_adj_5219));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i31_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 rem_4_i1593_3_lut (.I0(n2344), .I1(n2411), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2443));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i37_4_lut (.I0(n2704), .I1(n82), .I2(n6222), 
            .I3(n2724), .O(n37_adj_5222));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i37_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i21_4_lut (.I0(n2712), .I1(n90), .I2(n6230), 
            .I3(n2724), .O(n21_adj_5212));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i21_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 rem_4_i1592_3_lut (.I0(n2343), .I1(n2410), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2442));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i23_4_lut (.I0(n2711), .I1(n89), .I2(n6229), 
            .I3(n2724), .O(n23_adj_5213));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i23_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i25_4_lut (.I0(n2710), .I1(n88), .I2(n6228), 
            .I3(n2724), .O(n25_adj_5215));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i25_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 rem_4_add_1452_19_lut (.I0(GND_net), .I1(n2142), .I2(VCC_net), 
            .I3(n28968), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_27 (.CI(n28750), .I0(n2934), .I1(VCC_net), 
            .CO(n28751));
    SB_LUT4 rem_4_add_1988_26_lut (.I0(GND_net), .I1(n2935), .I2(VCC_net), 
            .I3(n28749), .O(n3002_adj_4761)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_26 (.CI(n28749), .I0(n2935), .I1(VCC_net), 
            .CO(n28750));
    SB_CARRY rem_4_add_1452_19 (.CI(n28968), .I0(n2142), .I1(VCC_net), 
            .CO(n28969));
    SB_LUT4 rem_4_add_1452_18_lut (.I0(GND_net), .I1(n2143), .I2(VCC_net), 
            .I3(n28967), .O(n2210)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_25_lut (.I0(GND_net), .I1(n2936), .I2(VCC_net), 
            .I3(n28748), .O(n3003_adj_4760)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1830_i17_4_lut (.I0(n2714), .I1(n92), .I2(n6232), 
            .I3(n2724), .O(n17_adj_5210));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i17_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 rem_4_i1590_3_lut (.I0(n2341), .I1(n2408), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2440));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1590_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1452_18 (.CI(n28967), .I0(n2143), .I1(VCC_net), 
            .CO(n28968));
    SB_CARRY rem_4_add_1988_25 (.CI(n28748), .I0(n2936), .I1(VCC_net), 
            .CO(n28749));
    SB_LUT4 div_46_LessThan_1830_i19_4_lut (.I0(n2713), .I1(n91), .I2(n6231), 
            .I3(n2724), .O(n19_adj_5211));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i19_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i9_4_lut (.I0(n2718), .I1(n96), .I2(n6236), 
            .I3(n2724), .O(n9_adj_5203));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i9_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4934));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1830_i7_4_lut (.I0(n2719), .I1(n97), .I2(n6237), 
            .I3(n2724), .O(n7_adj_5201));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i7_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i35_4_lut (.I0(n2705), .I1(n83), .I2(n6223), 
            .I3(n2724), .O(n35_adj_5221));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i35_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 rem_4_i1602_3_lut (.I0(n2353), .I1(n2420), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2452_adj_4882));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i11_4_lut (.I0(n2717), .I1(n95), .I2(n6235), 
            .I3(n2724), .O(n11_adj_5205));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i11_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i13_4_lut (.I0(n2716), .I1(n94), .I2(n6234), 
            .I3(n2724), .O(n13_adj_5207));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i13_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 rem_4_i1603_3_lut (.I0(n2354), .I1(n2421), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2453_adj_4881));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1452_17_lut (.I0(GND_net), .I1(n2144), .I2(VCC_net), 
            .I3(n28966), .O(n2211)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1830_i27_4_lut (.I0(n2709), .I1(n87), .I2(n6227), 
            .I3(n2724), .O(n27_adj_5216));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i27_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i15_4_lut (.I0(n2715), .I1(n93), .I2(n6233), 
            .I3(n2724), .O(n15_adj_5208));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i15_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_LessThan_1830_i33_4_lut (.I0(n2706), .I1(n84), .I2(n6224), 
            .I3(n2724), .O(n33_adj_5220));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i33_4_lut.LUT_INIT = 16'hc399;
    SB_LUT4 div_46_i1832_1_lut (.I0(n2801), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2802));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1832_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34449_4_lut (.I0(n27_adj_5216), .I1(n15_adj_5208), .I2(n13_adj_5207), 
            .I3(n11_adj_5205), .O(n41296));
    defparam i34449_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35732_3_lut (.I0(n2249), .I1(n2316), .I2(n2273_adj_4953), 
            .I3(GND_net), .O(n2348));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i35732_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i12_3_lut (.I0(n93), .I1(n84), .I2(n33_adj_5220), 
            .I3(GND_net), .O(n12_adj_5206));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_add_1988_24_lut (.I0(GND_net), .I1(n2937), .I2(VCC_net), 
            .I3(n28747), .O(n3004_adj_4759)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_24 (.CI(n28747), .I0(n2937), .I1(VCC_net), 
            .CO(n28748));
    SB_CARRY rem_4_add_1452_17 (.CI(n28966), .I0(n2144), .I1(VCC_net), 
            .CO(n28967));
    SB_LUT4 rem_4_add_1988_23_lut (.I0(GND_net), .I1(n2938), .I2(VCC_net), 
            .I3(n28746), .O(n3005_adj_4758)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35575_3_lut (.I0(n2348), .I1(n2415), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2447_adj_4887));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i35575_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34423_2_lut (.I0(n33_adj_5220), .I1(n15_adj_5208), .I2(GND_net), 
            .I3(GND_net), .O(n41270));
    defparam i34423_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_LessThan_1830_i10_3_lut (.I0(n95), .I1(n94), .I2(n13_adj_5207), 
            .I3(GND_net), .O(n10_adj_5204));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_add_1452_16_lut (.I0(GND_net), .I1(n2145), .I2(VCC_net), 
            .I3(n28965), .O(n2212)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_23 (.CI(n28746), .I0(n2938), .I1(VCC_net), 
            .CO(n28747));
    SB_CARRY rem_4_add_1452_16 (.CI(n28965), .I0(n2145), .I1(VCC_net), 
            .CO(n28966));
    SB_LUT4 div_46_LessThan_1830_i30_3_lut (.I0(n12_adj_5206), .I1(n83), 
            .I2(n35_adj_5221), .I3(GND_net), .O(n30_adj_5218));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_add_1452_15_lut (.I0(GND_net), .I1(n2146), .I2(VCC_net), 
            .I3(n28964), .O(n2213)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1828_3_lut (.I0(n2720), .I1(n6238), .I2(n2724), .I3(GND_net), 
            .O(n2798));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34516_3_lut (.I0(n7_adj_5201), .I1(n2798), .I2(n98), .I3(GND_net), 
            .O(n41363));
    defparam i34516_3_lut.LUT_INIT = 16'hebeb;
    SB_CARRY add_2357_22 (.CI(n28531), .I0(n43635), .I1(n671), .CO(n28532));
    SB_LUT4 i35132_4_lut (.I0(n13_adj_5207), .I1(n11_adj_5205), .I2(n9_adj_5203), 
            .I3(n41363), .O(n41979));
    defparam i35132_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35122_4_lut (.I0(n19_adj_5211), .I1(n17_adj_5210), .I2(n15_adj_5208), 
            .I3(n41979), .O(n41969));
    defparam i35122_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 rem_4_add_1988_22_lut (.I0(GND_net), .I1(n2939), .I2(VCC_net), 
            .I3(n28745), .O(n3006_adj_4757)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35834_4_lut (.I0(n25_adj_5215), .I1(n23_adj_5213), .I2(n21_adj_5212), 
            .I3(n41969), .O(n42681));
    defparam i35834_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_1988_22 (.CI(n28745), .I0(n2939), .I1(VCC_net), 
            .CO(n28746));
    SB_LUT4 i35402_4_lut (.I0(n31_adj_5219), .I1(n29_adj_5217), .I2(n27_adj_5216), 
            .I3(n42681), .O(n42249));
    defparam i35402_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35316_3_lut (.I0(n2250), .I1(n2317), .I2(n2273_adj_4953), 
            .I3(GND_net), .O(n2349));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i35316_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35317_3_lut (.I0(n2349), .I1(n2416), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2448_adj_4886));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i35317_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35920_4_lut (.I0(n37_adj_5222), .I1(n35_adj_5221), .I2(n33_adj_5220), 
            .I3(n42249), .O(n42767));
    defparam i35920_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1830_i16_3_lut (.I0(n91), .I1(n79), .I2(n43_adj_5225), 
            .I3(GND_net), .O(n16_adj_5209));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i16_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY rem_4_add_1452_15 (.CI(n28964), .I0(n2146), .I1(VCC_net), 
            .CO(n28965));
    SB_LUT4 rem_4_add_1988_21_lut (.I0(GND_net), .I1(n2940), .I2(VCC_net), 
            .I3(n28744), .O(n3007_adj_4756)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_14_lut (.I0(GND_net), .I1(n2147), .I2(VCC_net), 
            .I3(n28963), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_21 (.CI(n28744), .I0(n2940), .I1(VCC_net), 
            .CO(n28745));
    SB_LUT4 div_46_LessThan_1830_i6_3_lut (.I0(n98), .I1(n97), .I2(n7_adj_5201), 
            .I3(GND_net), .O(n6_adj_5200));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i6_3_lut.LUT_INIT = 16'h3535;
    SB_CARRY rem_4_add_1452_14 (.CI(n28963), .I0(n2147), .I1(VCC_net), 
            .CO(n28964));
    SB_LUT4 rem_4_add_1988_20_lut (.I0(GND_net), .I1(n2941), .I2(VCC_net), 
            .I3(n28743), .O(n3008_adj_4755)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35480_3_lut (.I0(n6_adj_5200), .I1(n90), .I2(n21_adj_5212), 
            .I3(GND_net), .O(n42327));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35480_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35481_3_lut (.I0(n42327), .I1(n89), .I2(n23_adj_5213), .I3(GND_net), 
            .O(n42328));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35481_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_2357_21_lut (.I0(n807), .I1(n43635), .I2(n806), .I3(n28530), 
            .O(displacement_23__N_229[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2357_21 (.CI(n28530), .I0(n43635), .I1(n806), .CO(n28531));
    SB_LUT4 add_2357_20_lut (.I0(n939), .I1(n43635), .I2(n938), .I3(n28529), 
            .O(displacement_23__N_229[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2357_20 (.CI(n28529), .I0(n43635), .I1(n938), .CO(n28530));
    SB_LUT4 i34479_4_lut (.I0(n21_adj_5212), .I1(n19_adj_5211), .I2(n17_adj_5210), 
            .I3(n9_adj_5203), .O(n41326));
    defparam i34479_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34391_2_lut (.I0(n43_adj_5225), .I1(n19_adj_5211), .I2(GND_net), 
            .I3(GND_net), .O(n41238));
    defparam i34391_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 rem_4_add_1452_13_lut (.I0(GND_net), .I1(n2148), .I2(VCC_net), 
            .I3(n28962), .O(n2215)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1596_3_lut (.I0(n2347), .I1(n2414), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2446));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i8_3_lut (.I0(n96), .I1(n92), .I2(n17_adj_5210), 
            .I3(GND_net), .O(n8_adj_5202));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_i1595_3_lut (.I0(n2346), .I1(n2413), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2445));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1594_3_lut (.I0(n2345), .I1(n2412), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2444));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35314_3_lut (.I0(n2253), .I1(n2320), .I2(n2273_adj_4953), 
            .I3(GND_net), .O(n2352));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i35314_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1452_13 (.CI(n28962), .I0(n2148), .I1(VCC_net), 
            .CO(n28963));
    SB_CARRY rem_4_add_1988_20 (.CI(n28743), .I0(n2941), .I1(VCC_net), 
            .CO(n28744));
    SB_LUT4 div_46_LessThan_1830_i24_3_lut (.I0(n16_adj_5209), .I1(n78), 
            .I2(n45_adj_5226), .I3(GND_net), .O(n24_adj_5214));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35315_3_lut (.I0(n2352), .I1(n2419), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2451_adj_4883));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i35315_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1600_3_lut (.I0(n2351), .I1(n2418), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2450_adj_4884));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34395_4_lut (.I0(n43_adj_5225), .I1(n25_adj_5215), .I2(n23_adj_5213), 
            .I3(n41326), .O(n41242));
    defparam i34395_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35617_4_lut (.I0(n24_adj_5214), .I1(n8_adj_5202), .I2(n45_adj_5226), 
            .I3(n41238), .O(n42464));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35617_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_2357_19_lut (.I0(n1068), .I1(n43635), .I2(n1067), .I3(n28528), 
            .O(displacement_23__N_229[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_19_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i34917_3_lut (.I0(n42328), .I1(n88), .I2(n25_adj_5215), .I3(GND_net), 
            .O(n41764));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34917_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i1829_3_lut (.I0(n1065), .I1(n6239), .I2(n2724), .I3(GND_net), 
            .O(n2799));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1829_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1830_i4_4_lut (.I0(n1066), .I1(n99), .I2(n2799), 
            .I3(n558), .O(n4_adj_5199));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1830_i4_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35478_3_lut (.I0(n4_adj_5199), .I1(n87), .I2(n27_adj_5216), 
            .I3(GND_net), .O(n42325));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35478_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_2357_19 (.CI(n28528), .I0(n43635), .I1(n1067), .CO(n28529));
    SB_LUT4 rem_4_add_1988_19_lut (.I0(GND_net), .I1(n2942), .I2(VCC_net), 
            .I3(n28742), .O(n3009_adj_4754)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_19 (.CI(n28742), .I0(n2942), .I1(VCC_net), 
            .CO(n28743));
    SB_LUT4 i35479_3_lut (.I0(n42325), .I1(n86), .I2(n29_adj_5217), .I3(GND_net), 
            .O(n42326));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35479_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35734_3_lut (.I0(n2251), .I1(n2318), .I2(n2273_adj_4953), 
            .I3(GND_net), .O(n2350));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i35734_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4933));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_1452_12_lut (.I0(GND_net), .I1(n2149), .I2(VCC_net), 
            .I3(n28961), .O(n2216)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35573_3_lut (.I0(n2350), .I1(n2417), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2449_adj_4885));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i35573_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1452_12 (.CI(n28961), .I0(n2149), .I1(VCC_net), 
            .CO(n28962));
    SB_LUT4 rem_4_add_1988_18_lut (.I0(GND_net), .I1(n2943_adj_4656), .I2(VCC_net), 
            .I3(n28741), .O(n3010_adj_4753)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34429_4_lut (.I0(n33_adj_5220), .I1(n31_adj_5219), .I2(n29_adj_5217), 
            .I3(n41296), .O(n41276));
    defparam i34429_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 rem_4_i1607_rep_52_3_lut (.I0(n2358_adj_4940), .I1(n2425), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2457_adj_4876));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1607_rep_52_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1605_3_lut (.I0(n2356), .I1(n2423), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2455_adj_4878));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2357_18_lut (.I0(n1194), .I1(n43635), .I2(n1193), .I3(n28527), 
            .O(displacement_23__N_229[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_18_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_i1604_3_lut (.I0(n2355), .I1(n2422), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2454_adj_4879));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35832_4_lut (.I0(n30_adj_5218), .I1(n10_adj_5204), .I2(n35_adj_5221), 
            .I3(n41270), .O(n42679));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35832_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34919_3_lut (.I0(n42326), .I1(n85), .I2(n31_adj_5219), .I3(GND_net), 
            .O(n41766));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34919_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_add_1452_11_lut (.I0(GND_net), .I1(n2150), .I2(VCC_net), 
            .I3(n28960), .O(n2217)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_18 (.CI(n28741), .I0(n2943_adj_4656), .I1(VCC_net), 
            .CO(n28742));
    SB_CARRY rem_4_add_1452_11 (.CI(n28960), .I0(n2150), .I1(VCC_net), 
            .CO(n28961));
    SB_LUT4 rem_4_i1524_3_lut (.I0(n2243), .I1(n2310), .I2(n2273_adj_4953), 
            .I3(GND_net), .O(n2342));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36006_4_lut (.I0(n41766), .I1(n42679), .I2(n35_adj_5221), 
            .I3(n41276), .O(n42853));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36006_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36007_3_lut (.I0(n42853), .I1(n82), .I2(n37_adj_5222), .I3(GND_net), 
            .O(n42854));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36007_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35952_3_lut (.I0(n42854), .I1(n81), .I2(n39_adj_5223), .I3(GND_net), 
            .O(n42799));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35952_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34397_4_lut (.I0(n43_adj_5225), .I1(n41_adj_5224), .I2(n39_adj_5223), 
            .I3(n42767), .O(n41244));
    defparam i34397_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35912_4_lut (.I0(n41764), .I1(n42464), .I2(n45_adj_5226), 
            .I3(n41242), .O(n42759));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35912_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 rem_4_i1523_3_lut (.I0(n2242), .I1(n2309), .I2(n2273_adj_4953), 
            .I3(GND_net), .O(n2341));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1523_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2357_18 (.CI(n28527), .I0(n43635), .I1(n1193), .CO(n28528));
    SB_LUT4 add_2357_17_lut (.I0(n1317), .I1(n43635), .I2(n1316), .I3(n28526), 
            .O(displacement_23__N_229[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1988_17_lut (.I0(GND_net), .I1(n2944_adj_4777), .I2(VCC_net), 
            .I3(n28740), .O(n3011_adj_4752)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34925_3_lut (.I0(n42799), .I1(n80), .I2(n41_adj_5224), .I3(GND_net), 
            .O(n41772));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34925_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i1807_3_lut (.I0(n2699), .I1(n6217), .I2(n2724), .I3(GND_net), 
            .O(n2777));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1807_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35914_4_lut (.I0(n41772), .I1(n42759), .I2(n45_adj_5226), 
            .I3(n41244), .O(n42761));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35914_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35915_3_lut (.I0(n42761), .I1(n77), .I2(n2777), .I3(GND_net), 
            .O(n2801));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35915_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 rem_4_i1522_3_lut (.I0(n2241), .I1(n2308), .I2(n2273_adj_4953), 
            .I3(GND_net), .O(n2340));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1522_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1988_17 (.CI(n28740), .I0(n2944_adj_4777), .I1(VCC_net), 
            .CO(n28741));
    SB_CARRY add_2357_17 (.CI(n28526), .I0(n43635), .I1(n1316), .CO(n28527));
    SB_LUT4 add_2357_16_lut (.I0(n1437), .I1(n43635), .I2(n1436), .I3(n28525), 
            .O(displacement_23__N_229[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i6_4_lut (.I0(n17011), .I1(\data_in_frame[14] [1]), .I2(n35626), 
            .I3(n35463), .O(n16_adj_5332));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1728 (.I0(\data_in_frame[9] [5]), .I1(n35562), 
            .I2(n35644), .I3(\data_in_frame[9] [6]), .O(n17_adj_5330));
    defparam i7_4_lut_adj_1728.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1729 (.I0(n17_adj_5330), .I1(\data_in_frame[6] [7]), 
            .I2(n16_adj_5332), .I3(n16086), .O(n37132));
    defparam i9_4_lut_adj_1729.LUT_INIT = 16'h6996;
    SB_LUT4 rem_4_add_1452_10_lut (.I0(GND_net), .I1(n2151), .I2(VCC_net), 
            .I3(n28959), .O(n2218)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1988_16_lut (.I0(GND_net), .I1(n2945_adj_4654), .I2(VCC_net), 
            .I3(n28739), .O(n3012_adj_4751)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_10 (.CI(n28959), .I0(n2151), .I1(VCC_net), 
            .CO(n28960));
    SB_CARRY rem_4_add_1988_16 (.CI(n28739), .I0(n2945_adj_4654), .I1(VCC_net), 
            .CO(n28740));
    SB_LUT4 rem_4_add_1452_9_lut (.I0(GND_net), .I1(n2152), .I2(VCC_net), 
            .I3(n28958), .O(n2219)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_9_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_11_pad (.PACKAGE_PIN(PIN_11), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_11_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_11_pad.PIN_TYPE = 6'b011001;
    defparam PIN_11_pad.PULLUP = 1'b0;
    defparam PIN_11_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_11_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 rem_4_add_1988_15_lut (.I0(GND_net), .I1(n2946_adj_4776), .I2(VCC_net), 
            .I3(n28738), .O(n3013_adj_4750)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1529_3_lut (.I0(n2248), .I1(n2315), .I2(n2273_adj_4953), 
            .I3(GND_net), .O(n2347));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1529_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1452_9 (.CI(n28958), .I0(n2152), .I1(VCC_net), 
            .CO(n28959));
    SB_CARRY rem_4_add_1988_15 (.CI(n28738), .I0(n2946_adj_4776), .I1(VCC_net), 
            .CO(n28739));
    SB_CARRY add_2357_16 (.CI(n28525), .I0(n43635), .I1(n1436), .CO(n28526));
    SB_LUT4 add_2357_15_lut (.I0(n1554_adj_4743), .I1(n43635), .I2(n1553_adj_4742), 
            .I3(n28524), .O(displacement_23__N_229[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1452_8_lut (.I0(GND_net), .I1(n2153), .I2(VCC_net), 
            .I3(n28957), .O(n2220)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2357_15 (.CI(n28524), .I0(n43635), .I1(n1553_adj_4742), 
            .CO(n28525));
    SB_CARRY rem_4_add_1452_8 (.CI(n28957), .I0(n2153), .I1(VCC_net), 
            .CO(n28958));
    SB_LUT4 add_2357_14_lut (.I0(n1668), .I1(n43635), .I2(n1667), .I3(n28523), 
            .O(displacement_23__N_229[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1988_14_lut (.I0(GND_net), .I1(n2947_adj_4655), .I2(VCC_net), 
            .I3(n28737), .O(n3014_adj_4749)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_7_lut (.I0(GND_net), .I1(n2154), .I2(GND_net), 
            .I3(n28956), .O(n2221)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_14 (.CI(n28737), .I0(n2947_adj_4655), .I1(VCC_net), 
            .CO(n28738));
    SB_CARRY rem_4_add_1452_7 (.CI(n28956), .I0(n2154), .I1(GND_net), 
            .CO(n28957));
    SB_CARRY add_2357_14 (.CI(n28523), .I0(n43635), .I1(n1667), .CO(n28524));
    SB_LUT4 rem_4_add_1452_6_lut (.I0(GND_net), .I1(n2155), .I2(GND_net), 
            .I3(n28955), .O(n2222)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1777_i31_2_lut (.I0(n2707), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5194));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1988_13_lut (.I0(GND_net), .I1(n2948_adj_4775), .I2(VCC_net), 
            .I3(n28736), .O(n3015_adj_4748)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2357_13_lut (.I0(n1779), .I1(n43635), .I2(n1778), .I3(n28522), 
            .O(displacement_23__N_229[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_13_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_i1533_rep_53_3_lut (.I0(n2252), .I1(n2319), .I2(n2273_adj_4953), 
            .I3(GND_net), .O(n2351));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1533_rep_53_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1528_3_lut (.I0(n2247), .I1(n2314), .I2(n2273_adj_4953), 
            .I3(GND_net), .O(n2346));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1528_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1452_6 (.CI(n28955), .I0(n2155), .I1(GND_net), 
            .CO(n28956));
    SB_LUT4 rem_4_i1526_3_lut (.I0(n2245), .I1(n2312), .I2(n2273_adj_4953), 
            .I3(GND_net), .O(n2344));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1526_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1988_13 (.CI(n28736), .I0(n2948_adj_4775), .I1(VCC_net), 
            .CO(n28737));
    SB_CARRY add_2357_13 (.CI(n28522), .I0(n43635), .I1(n1778), .CO(n28523));
    SB_LUT4 add_2357_12_lut (.I0(n1887), .I1(n43635), .I2(n1886), .I3(n28521), 
            .O(displacement_23__N_229[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2357_12 (.CI(n28521), .I0(n43635), .I1(n1886), .CO(n28522));
    SB_LUT4 div_46_LessThan_1777_i33_2_lut (.I0(n2706), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5196));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1988_12_lut (.I0(GND_net), .I1(n2949_adj_4774), .I2(VCC_net), 
            .I3(n28735), .O(n3016_adj_4747)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1452_5_lut (.I0(GND_net), .I1(n2156), .I2(VCC_net), 
            .I3(n28954), .O(n2223)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1452_5 (.CI(n28954), .I0(n2156), .I1(VCC_net), 
            .CO(n28955));
    SB_LUT4 rem_4_add_1452_4_lut (.I0(GND_net), .I1(n2157), .I2(VCC_net), 
            .I3(n28953), .O(n2224)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2357_11_lut (.I0(n1992), .I1(n43635), .I2(n1991), .I3(n28520), 
            .O(displacement_23__N_229[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1452_4 (.CI(n28953), .I0(n2157), .I1(VCC_net), 
            .CO(n28954));
    SB_LUT4 rem_4_add_1452_3_lut (.I0(GND_net), .I1(n2158), .I2(GND_net), 
            .I3(n28952), .O(n2225)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1452_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1527_3_lut (.I0(n2246), .I1(n2313), .I2(n2273_adj_4953), 
            .I3(GND_net), .O(n2345));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1777_i37_2_lut (.I0(n2704), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5198));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i37_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1452_3 (.CI(n28952), .I0(n2158), .I1(GND_net), 
            .CO(n28953));
    SB_CARRY add_2357_11 (.CI(n28520), .I0(n43635), .I1(n1991), .CO(n28521));
    SB_CARRY rem_4_add_1988_12 (.CI(n28735), .I0(n2949_adj_4774), .I1(VCC_net), 
            .CO(n28736));
    SB_CARRY rem_4_add_1452_2 (.CI(VCC_net), .I0(n2258), .I1(VCC_net), 
            .CO(n28952));
    SB_LUT4 div_46_LessThan_1777_i21_2_lut (.I0(n2712), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5188));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i23_2_lut (.I0(n2711), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5189));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1519_21_lut (.I0(n2273_adj_4953), .I1(n2240), .I2(VCC_net), 
            .I3(n28951), .O(n2339)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_46_LessThan_1777_i35_2_lut (.I0(n2705), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5197));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i2_3_lut (.I0(encoder0_position[1]), .I1(n24_adj_4712), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n1065));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1525_3_lut (.I0(n2244), .I1(n2311), .I2(n2273_adj_4953), 
            .I3(GND_net), .O(n2343));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1525_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2357_10_lut (.I0(n2094), .I1(n43635), .I2(n2093), .I3(n28519), 
            .O(displacement_23__N_229[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1988_11_lut (.I0(GND_net), .I1(n2950_adj_4773), .I2(VCC_net), 
            .I3(n28734), .O(n3017)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2357_10 (.CI(n28519), .I0(n43635), .I1(n2093), .CO(n28520));
    SB_LUT4 add_2357_9_lut (.I0(n2193), .I1(n43635), .I2(n2192), .I3(n28518), 
            .O(displacement_23__N_229[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_46_LessThan_1777_i25_2_lut (.I0(n2710), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5191));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i25_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2357_9 (.CI(n28518), .I0(n43635), .I1(n2192), .CO(n28519));
    SB_LUT4 add_2357_8_lut (.I0(n2289), .I1(n43635), .I2(n2288), .I3(n28517), 
            .O(displacement_23__N_229[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_8_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2357_8 (.CI(n28517), .I0(n43635), .I1(n2288), .CO(n28518));
    SB_LUT4 rem_4_add_1519_20_lut (.I0(GND_net), .I1(n2241), .I2(VCC_net), 
            .I3(n28950), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_11 (.CI(n28734), .I0(n2950_adj_4773), .I1(VCC_net), 
            .CO(n28735));
    SB_LUT4 div_46_LessThan_1777_i27_2_lut (.I0(n2709), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5192));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i27_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1519_20 (.CI(n28950), .I0(n2241), .I1(VCC_net), 
            .CO(n28951));
    SB_LUT4 add_2357_7_lut (.I0(n2382), .I1(n43635), .I2(n2381), .I3(n28516), 
            .O(displacement_23__N_229[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2357_7 (.CI(n28516), .I0(n43635), .I1(n2381), .CO(n28517));
    SB_LUT4 rem_4_add_1988_10_lut (.I0(GND_net), .I1(n2951_adj_4772), .I2(VCC_net), 
            .I3(n28733), .O(n3018)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_19_lut (.I0(GND_net), .I1(n2242), .I2(VCC_net), 
            .I3(n28949), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_10 (.CI(n28733), .I0(n2951_adj_4772), .I1(VCC_net), 
            .CO(n28734));
    SB_CARRY rem_4_add_1519_19 (.CI(n28949), .I0(n2242), .I1(VCC_net), 
            .CO(n28950));
    SB_LUT4 rem_4_add_1988_9_lut (.I0(GND_net), .I1(n2952_adj_4771), .I2(VCC_net), 
            .I3(n28732), .O(n3019)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1777_i9_2_lut (.I0(n2718), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_5179));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i9_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i1537_3_lut (.I0(n2256), .I1(n2323), .I2(n2273_adj_4953), 
            .I3(GND_net), .O(n2355));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1536_3_lut (.I0(n2255), .I1(n2322), .I2(n2273_adj_4953), 
            .I3(GND_net), .O(n2354));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1777_i13_2_lut (.I0(n2716), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5183));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i15_2_lut (.I0(n2715), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5185));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1519_18_lut (.I0(GND_net), .I1(n2243), .I2(VCC_net), 
            .I3(n28948), .O(n2310)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_18 (.CI(n28948), .I0(n2243), .I1(VCC_net), 
            .CO(n28949));
    SB_CARRY rem_4_add_1988_9 (.CI(n28732), .I0(n2952_adj_4771), .I1(VCC_net), 
            .CO(n28733));
    SB_LUT4 div_46_LessThan_1777_i17_2_lut (.I0(n2714), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5186));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1519_17_lut (.I0(GND_net), .I1(n2244), .I2(VCC_net), 
            .I3(n28947), .O(n2311)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_17 (.CI(n28947), .I0(n2244), .I1(VCC_net), 
            .CO(n28948));
    SB_LUT4 add_2357_6_lut (.I0(n2472), .I1(n43635), .I2(n2471), .I3(n28515), 
            .O(displacement_23__N_229[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1988_8_lut (.I0(GND_net), .I1(n2953_adj_4770), .I2(VCC_net), 
            .I3(n28731), .O(n3020)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_16_lut (.I0(GND_net), .I1(n2245), .I2(VCC_net), 
            .I3(n28946), .O(n2312)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_16 (.CI(n28946), .I0(n2245), .I1(VCC_net), 
            .CO(n28947));
    SB_CARRY rem_4_add_1988_8 (.CI(n28731), .I0(n2953_adj_4770), .I1(VCC_net), 
            .CO(n28732));
    SB_LUT4 div_46_LessThan_1777_i29_2_lut (.I0(n2708), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5193));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i1463_3_lut (.I0(n2150), .I1(n2217), .I2(n2174_adj_4984), 
            .I3(GND_net), .O(n2249));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1519_15_lut (.I0(GND_net), .I1(n2246), .I2(VCC_net), 
            .I3(n28945), .O(n2313)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_15 (.CI(n28945), .I0(n2246), .I1(VCC_net), 
            .CO(n28946));
    SB_LUT4 rem_4_add_1988_7_lut (.I0(GND_net), .I1(n2954_adj_4769), .I2(GND_net), 
            .I3(n28730), .O(n3021)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2357_6 (.CI(n28515), .I0(n43635), .I1(n2471), .CO(n28516));
    SB_CARRY rem_4_add_1988_7 (.CI(n28730), .I0(n2954_adj_4769), .I1(GND_net), 
            .CO(n28731));
    SB_LUT4 rem_4_add_1988_6_lut (.I0(GND_net), .I1(n2955_adj_4768), .I2(GND_net), 
            .I3(n28729), .O(n3022)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_6 (.CI(n28729), .I0(n2955_adj_4768), .I1(GND_net), 
            .CO(n28730));
    SB_LUT4 rem_4_add_1519_14_lut (.I0(GND_net), .I1(n2247), .I2(VCC_net), 
            .I3(n28944), .O(n2314)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2357_5_lut (.I0(n2559), .I1(n43635), .I2(n2558), .I3(n28514), 
            .O(displacement_23__N_229[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2357_5 (.CI(n28514), .I0(n43635), .I1(n2558), .CO(n28515));
    SB_LUT4 add_2357_4_lut (.I0(n2643), .I1(n43635), .I2(n2642), .I3(n28513), 
            .O(displacement_23__N_229[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2357_4 (.CI(n28513), .I0(n43635), .I1(n2642), .CO(n28514));
    SB_LUT4 div_46_LessThan_1777_i11_2_lut (.I0(n2717), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5181));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1777_i19_2_lut (.I0(n2713), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5187));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1779_1_lut (.I0(n2723), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1779_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34624_4_lut (.I0(n29_adj_5193), .I1(n17_adj_5186), .I2(n15_adj_5185), 
            .I3(n13_adj_5183), .O(n41471));
    defparam i34624_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY rem_4_add_1519_14 (.CI(n28944), .I0(n2247), .I1(VCC_net), 
            .CO(n28945));
    SB_LUT4 rem_4_add_1988_5_lut (.I0(GND_net), .I1(n2956_adj_4767), .I2(VCC_net), 
            .I3(n28728), .O(n3023)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1461_3_lut (.I0(n2148), .I1(n2215), .I2(n2174_adj_4984), 
            .I3(GND_net), .O(n2247));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34660_4_lut (.I0(n11_adj_5181), .I1(n9_adj_5179), .I2(n2719), 
            .I3(n98), .O(n41507));
    defparam i34660_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i35228_4_lut (.I0(n17_adj_5186), .I1(n15_adj_5185), .I2(n13_adj_5183), 
            .I3(n41507), .O(n42075));
    defparam i35228_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35220_4_lut (.I0(n23_adj_5189), .I1(n21_adj_5188), .I2(n19_adj_5187), 
            .I3(n42075), .O(n42067));
    defparam i35220_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33910_4_lut (.I0(n29_adj_5193), .I1(n27_adj_5192), .I2(n25_adj_5191), 
            .I3(n42067), .O(n40756));
    defparam i33910_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1777_i6_4_lut (.I0(n1065), .I1(n99), .I2(n2720), 
            .I3(n558), .O(n6_adj_5177));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i6_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 rem_4_add_1519_13_lut (.I0(GND_net), .I1(n2248), .I2(VCC_net), 
            .I3(n28943), .O(n2315)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_5 (.CI(n28728), .I0(n2956_adj_4767), .I1(VCC_net), 
            .CO(n28729));
    SB_LUT4 rem_4_i1459_3_lut (.I0(n2146), .I1(n2213), .I2(n2174_adj_4984), 
            .I3(GND_net), .O(n2245));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35488_3_lut (.I0(n6_adj_5177), .I1(n87), .I2(n29_adj_5193), 
            .I3(GND_net), .O(n42335));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35488_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_2357_3_lut (.I0(n2724), .I1(n43635), .I2(n2723), .I3(n28512), 
            .O(displacement_23__N_229[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2357_3 (.CI(n28512), .I0(n43635), .I1(n2723), .CO(n28513));
    SB_CARRY rem_4_add_1519_13 (.CI(n28943), .I0(n2248), .I1(VCC_net), 
            .CO(n28944));
    SB_LUT4 rem_4_add_1988_4_lut (.I0(GND_net), .I1(n2957_adj_4765), .I2(VCC_net), 
            .I3(n28727), .O(n3024)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2357_2_lut (.I0(n2802), .I1(n43635), .I2(n2801), .I3(VCC_net), 
            .O(displacement_23__N_229[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2357_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_2357_2 (.CI(VCC_net), .I0(n43635), .I1(n2801), .CO(n28512));
    SB_LUT4 div_46_LessThan_1777_i32_3_lut (.I0(n14_adj_5184), .I1(n83), 
            .I2(n37_adj_5198), .I3(GND_net), .O(n32_adj_5195));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35489_3_lut (.I0(n42335), .I1(n86), .I2(n31_adj_5194), .I3(GND_net), 
            .O(n42336));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35489_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_i1457_3_lut (.I0(n2144), .I1(n2211), .I2(n2174_adj_4984), 
            .I3(GND_net), .O(n2243));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1519_12_lut (.I0(GND_net), .I1(n2249), .I2(VCC_net), 
            .I3(n28942), .O(n2316)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2355_25_lut (.I0(GND_net), .I1(n2699), .I2(n78), .I3(n28511), 
            .O(n6217)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2355_24_lut (.I0(GND_net), .I1(n2700), .I2(n79), .I3(n28510), 
            .O(n6218)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2355_24 (.CI(n28510), .I0(n2700), .I1(n79), .CO(n28511));
    SB_CARRY rem_4_add_1988_4 (.CI(n28727), .I0(n2957_adj_4765), .I1(VCC_net), 
            .CO(n28728));
    SB_CARRY rem_4_add_1519_12 (.CI(n28942), .I0(n2249), .I1(VCC_net), 
            .CO(n28943));
    SB_LUT4 rem_4_add_1988_3_lut (.I0(GND_net), .I1(n2958_adj_4764), .I2(GND_net), 
            .I3(n28726), .O(n3025)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1988_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_11_lut (.I0(GND_net), .I1(n2250), .I2(VCC_net), 
            .I3(n28941), .O(n2317)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1988_3 (.CI(n28726), .I0(n2958_adj_4764), .I1(GND_net), 
            .CO(n28727));
    SB_LUT4 i34593_4_lut (.I0(n35_adj_5197), .I1(n33_adj_5196), .I2(n31_adj_5194), 
            .I3(n41471), .O(n41440));
    defparam i34593_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_2355_23_lut (.I0(GND_net), .I1(n2701), .I2(n80), .I3(n28509), 
            .O(n6219)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1458_3_lut (.I0(n2145), .I1(n2212), .I2(n2174_adj_4984), 
            .I3(GND_net), .O(n2244));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1458_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2355_23 (.CI(n28509), .I0(n2701), .I1(n80), .CO(n28510));
    SB_LUT4 add_2355_22_lut (.I0(GND_net), .I1(n2702), .I2(n81), .I3(n28508), 
            .O(n6220)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35818_4_lut (.I0(n32_adj_5195), .I1(n12_adj_5182), .I2(n37_adj_5198), 
            .I3(n41426), .O(n42665));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35818_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34905_3_lut (.I0(n42336), .I1(n85), .I2(n33_adj_5196), .I3(GND_net), 
            .O(n41752));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34905_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_1519_11 (.CI(n28941), .I0(n2250), .I1(VCC_net), 
            .CO(n28942));
    SB_CARRY rem_4_add_1988_2 (.CI(VCC_net), .I0(n3058), .I1(VCC_net), 
            .CO(n28726));
    SB_CARRY add_2355_22 (.CI(n28508), .I0(n2702), .I1(n81), .CO(n28509));
    SB_LUT4 i35705_3_lut (.I0(n8_adj_5178), .I1(n90), .I2(n23_adj_5189), 
            .I3(GND_net), .O(n42552));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35705_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_2355_21_lut (.I0(GND_net), .I1(n2703), .I2(n82), .I3(n28507), 
            .O(n6221)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2355_21 (.CI(n28507), .I0(n2703), .I1(n82), .CO(n28508));
    SB_LUT4 add_2355_20_lut (.I0(GND_net), .I1(n2704), .I2(n83), .I3(n28506), 
            .O(n6222)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2355_20 (.CI(n28506), .I0(n2704), .I1(n83), .CO(n28507));
    SB_LUT4 add_2355_19_lut (.I0(GND_net), .I1(n2705), .I2(n84), .I3(n28505), 
            .O(n6223)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2355_19 (.CI(n28505), .I0(n2705), .I1(n84), .CO(n28506));
    SB_LUT4 add_2355_18_lut (.I0(GND_net), .I1(n2706), .I2(n85), .I3(n28504), 
            .O(n6224)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1456_3_lut (.I0(n2143), .I1(n2210), .I2(n2174_adj_4984), 
            .I3(GND_net), .O(n2242));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35706_3_lut (.I0(n42552), .I1(n89), .I2(n25_adj_5191), .I3(GND_net), 
            .O(n42553));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35706_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34632_4_lut (.I0(n25_adj_5191), .I1(n23_adj_5189), .I2(n21_adj_5188), 
            .I3(n40770), .O(n41479));
    defparam i34632_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 rem_4_i1469_3_lut (.I0(n2156), .I1(n2223), .I2(n2174_adj_4984), 
            .I3(GND_net), .O(n2255));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35615_3_lut (.I0(n10_adj_5180), .I1(n91), .I2(n21_adj_5188), 
            .I3(GND_net), .O(n42462));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35615_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_i1460_3_lut (.I0(n2147), .I1(n2214), .I2(n2174_adj_4984), 
            .I3(GND_net), .O(n2246));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35614_3_lut (.I0(n42553), .I1(n88), .I2(n27_adj_5192), .I3(GND_net), 
            .O(n24_adj_5190));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35614_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_i1468_3_lut (.I0(n2155), .I1(n2222), .I2(n2174_adj_4984), 
            .I3(GND_net), .O(n2254));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35460_4_lut (.I0(n35_adj_5197), .I1(n33_adj_5196), .I2(n31_adj_5194), 
            .I3(n40756), .O(n42307));
    defparam i35460_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1466_3_lut (.I0(n2153), .I1(n2220), .I2(n2174_adj_4984), 
            .I3(GND_net), .O(n2252));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1466_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2355_18 (.CI(n28504), .I0(n2706), .I1(n85), .CO(n28505));
    SB_LUT4 rem_4_i1464_3_lut (.I0(n2151), .I1(n2218), .I2(n2174_adj_4984), 
            .I3(GND_net), .O(n2250));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36002_4_lut (.I0(n41752), .I1(n42665), .I2(n37_adj_5198), 
            .I3(n41440), .O(n42849));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36002_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35689_4_lut (.I0(n24_adj_5190), .I1(n42462), .I2(n27_adj_5192), 
            .I3(n41479), .O(n42536));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35689_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36034_4_lut (.I0(n42536), .I1(n42849), .I2(n37_adj_5198), 
            .I3(n42307), .O(n42881));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36034_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_2355_17_lut (.I0(GND_net), .I1(n2707), .I2(n86), .I3(n28503), 
            .O(n6225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1462_3_lut (.I0(n2149), .I1(n2216), .I2(n2174_adj_4984), 
            .I3(GND_net), .O(n2248));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2055_29_lut (.I0(n3065), .I1(n3032), .I2(VCC_net), 
            .I3(n28725), .O(n3131)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i36035_3_lut (.I0(n42881), .I1(n82), .I2(n2703), .I3(GND_net), 
            .O(n42882));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36035_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i36031_3_lut (.I0(n42882), .I1(n81), .I2(n2702), .I3(GND_net), 
            .O(n42878));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36031_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35874_3_lut (.I0(n42878), .I1(n80), .I2(n2701), .I3(GND_net), 
            .O(n42721));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35874_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35875_3_lut (.I0(n42721), .I1(n79), .I2(n2700), .I3(GND_net), 
            .O(n42722));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35875_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i2048_4_lut (.I0(n42722), .I1(n77), .I2(n78), .I3(n2699), 
            .O(n2723));
    defparam i2048_4_lut.LUT_INIT = 16'hceef;
    SB_LUT4 rem_4_i1455_3_lut (.I0(n2142), .I1(n2209), .I2(n2174_adj_4984), 
            .I3(GND_net), .O(n2241));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13142_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n13302), 
            .I3(GND_net), .O(n17881));   // verilog/coms.v(127[12] 295[6])
    defparam i13142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13143_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n13302), 
            .I3(GND_net), .O(n17882));   // verilog/coms.v(127[12] 295[6])
    defparam i13143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13144_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n13302), 
            .I3(GND_net), .O(n17883));   // verilog/coms.v(127[12] 295[6])
    defparam i13144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13145_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n13302), 
            .I3(GND_net), .O(n17884));   // verilog/coms.v(127[12] 295[6])
    defparam i13145_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2355_17 (.CI(n28503), .I0(n2707), .I1(n86), .CO(n28504));
    SB_LUT4 i13146_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n13302), 
            .I3(GND_net), .O(n17885));   // verilog/coms.v(127[12] 295[6])
    defparam i13146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1398_rep_71_3_lut (.I0(n2053), .I1(n2120), .I2(n2075_adj_5028), 
            .I3(GND_net), .O(n2152));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1398_rep_71_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(clk32MHz), .D(displacement_23__N_80[23]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_LUT4 i13147_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n13302), 
            .I3(GND_net), .O(n17886));   // verilog/coms.v(127[12] 295[6])
    defparam i13147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1730 (.I0(n1056), .I1(n1057), .I2(n1058), .I3(GND_net), 
            .O(n35946));
    defparam i1_3_lut_adj_1730.LUT_INIT = 16'hfefe;
    SB_LUT4 i13148_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n13302), 
            .I3(GND_net), .O(n17887));   // verilog/coms.v(127[12] 295[6])
    defparam i13148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1399_3_lut (.I0(n2054), .I1(n2121), .I2(n2075_adj_5028), 
            .I3(GND_net), .O(n2153));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2355_16_lut (.I0(GND_net), .I1(n2708), .I2(n87), .I3(n28502), 
            .O(n6226)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_10_lut (.I0(GND_net), .I1(n2251), .I2(VCC_net), 
            .I3(n28940), .O(n2318)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2355_16 (.CI(n28502), .I0(n2708), .I1(n87), .CO(n28503));
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(clk32MHz), .D(displacement_23__N_80[22]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_CARRY rem_4_add_1519_10 (.CI(n28940), .I0(n2251), .I1(VCC_net), 
            .CO(n28941));
    SB_LUT4 i13149_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n13302), 
            .I3(GND_net), .O(n17888));   // verilog/coms.v(127[12] 295[6])
    defparam i13149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13393_3_lut (.I0(\data_in_frame[24] [6]), .I1(rx_data[6]), 
            .I2(n36526), .I3(GND_net), .O(n18132));   // verilog/coms.v(127[12] 295[6])
    defparam i13393_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2355_15_lut (.I0(GND_net), .I1(n2709), .I2(n88), .I3(n28501), 
            .O(n6227)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2355_15 (.CI(n28501), .I0(n2709), .I1(n88), .CO(n28502));
    SB_LUT4 i13150_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n13302), 
            .I3(GND_net), .O(n17889));   // verilog/coms.v(127[12] 295[6])
    defparam i13150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13392_3_lut (.I0(\data_in_frame[24] [5]), .I1(rx_data[5]), 
            .I2(n36526), .I3(GND_net), .O(n18131));   // verilog/coms.v(127[12] 295[6])
    defparam i13392_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13391_3_lut (.I0(\data_in_frame[24] [4]), .I1(rx_data[4]), 
            .I2(n36526), .I3(GND_net), .O(n18130));   // verilog/coms.v(127[12] 295[6])
    defparam i13391_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1392_3_lut (.I0(n2047), .I1(n2114), .I2(n2075_adj_5028), 
            .I3(GND_net), .O(n2146));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1392_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2355_14_lut (.I0(GND_net), .I1(n2710), .I2(n89), .I3(n28500), 
            .O(n6228)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13151_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n13302), 
            .I3(GND_net), .O(n17890));   // verilog/coms.v(127[12] 295[6])
    defparam i13151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13390_3_lut (.I0(\data_in_frame[24] [3]), .I1(rx_data[3]), 
            .I2(n36526), .I3(GND_net), .O(n18129));   // verilog/coms.v(127[12] 295[6])
    defparam i13390_3_lut.LUT_INIT = 16'hacac;
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(clk32MHz), .D(displacement_23__N_80[21]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(clk32MHz), .D(displacement_23__N_80[20]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(clk32MHz), .D(displacement_23__N_80[19]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(clk32MHz), .D(displacement_23__N_80[18]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(clk32MHz), .D(displacement_23__N_80[17]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(clk32MHz), .D(displacement_23__N_80[16]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(clk32MHz), .D(displacement_23__N_80[15]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(clk32MHz), .D(displacement_23__N_80[14]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(clk32MHz), .D(displacement_23__N_80[13]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(clk32MHz), .D(displacement_23__N_80[12]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(clk32MHz), .D(displacement_23__N_80[11]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(clk32MHz), .D(displacement_23__N_80[10]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(clk32MHz), .D(displacement_23__N_80[9]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(clk32MHz), .D(displacement_23__N_80[8]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(clk32MHz), .D(displacement_23__N_80[7]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(clk32MHz), .D(displacement_23__N_80[6]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(clk32MHz), .D(displacement_23__N_80[5]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(clk32MHz), .D(displacement_23__N_80[4]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(clk32MHz), .D(displacement_23__N_80[3]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(clk32MHz), .D(displacement_23__N_80[2]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(clk32MHz), .D(displacement_23__N_80[1]));   // verilog/TinyFPGA_B.v(231[10] 233[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[22]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[21]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[20]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[19]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[18]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[17]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[16]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[15]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[14]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_CARRY add_2355_14 (.CI(n28500), .I0(n2710), .I1(n89), .CO(n28501));
    SB_LUT4 i13389_3_lut (.I0(\data_in_frame[24] [2]), .I1(rx_data[2]), 
            .I2(n36526), .I3(GND_net), .O(n18128));   // verilog/coms.v(127[12] 295[6])
    defparam i13389_3_lut.LUT_INIT = 16'hacac;
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[13]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[12]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[11]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[10]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[9]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[8]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[7]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_LUT4 i13152_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n13302), 
            .I3(GND_net), .O(n17891));   // verilog/coms.v(127[12] 295[6])
    defparam i13152_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[6]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[5]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_LUT4 rem_4_add_2055_28_lut (.I0(GND_net), .I1(n3033), .I2(VCC_net), 
            .I3(n28724), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_28_lut.LUT_INIT = 16'hC33C;
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[4]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[3]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[2]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(clk32MHz), .D(pwm_setpoint_22__N_57[1]));   // verilog/TinyFPGA_B.v(139[10] 152[6])
    SB_LUT4 i13388_3_lut (.I0(\data_in_frame[24] [1]), .I1(rx_data[1]), 
            .I2(n36526), .I3(GND_net), .O(n18127));   // verilog/coms.v(127[12] 295[6])
    defparam i13388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1391_3_lut (.I0(n2046), .I1(n2113), .I2(n2075_adj_5028), 
            .I3(GND_net), .O(n2145));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1391_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13153_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n13302), 
            .I3(GND_net), .O(n17892));   // verilog/coms.v(127[12] 295[6])
    defparam i13153_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13154_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n13302), 
            .I3(GND_net), .O(n17893));   // verilog/coms.v(127[12] 295[6])
    defparam i13154_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2055_28 (.CI(n28724), .I0(n3033), .I1(VCC_net), 
            .CO(n28725));
    SB_LUT4 i13512_3_lut (.I0(setpoint[22]), .I1(n4408), .I2(n37622), 
            .I3(GND_net), .O(n18251));   // verilog/coms.v(127[12] 295[6])
    defparam i13512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1722_i45_2_lut (.I0(n2619), .I1(n80), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_5176));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2355_13_lut (.I0(GND_net), .I1(n2711), .I2(n90), .I3(n28499), 
            .O(n6229)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2355_13 (.CI(n28499), .I0(n2711), .I1(n90), .CO(n28500));
    SB_LUT4 add_2355_12_lut (.I0(GND_net), .I1(n2712), .I2(n91), .I3(n28498), 
            .O(n6230)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1390_3_lut (.I0(n2045), .I1(n2112), .I2(n2075_adj_5028), 
            .I3(GND_net), .O(n2144));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1390_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2355_12 (.CI(n28498), .I0(n2712), .I1(n91), .CO(n28499));
    SB_LUT4 add_2355_11_lut (.I0(GND_net), .I1(n2713), .I2(n92), .I3(n28497), 
            .O(n6231)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2355_11 (.CI(n28497), .I0(n2713), .I1(n92), .CO(n28498));
    SB_LUT4 add_2355_10_lut (.I0(GND_net), .I1(n2714), .I2(n93), .I3(n28496), 
            .O(n6232)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1722_i43_2_lut (.I0(n2620), .I1(n81), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5174));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i43_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2355_10 (.CI(n28496), .I0(n2714), .I1(n93), .CO(n28497));
    SB_LUT4 div_46_LessThan_1722_i41_2_lut (.I0(n2621), .I1(n82), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5173));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1519_9_lut (.I0(GND_net), .I1(n2252), .I2(VCC_net), 
            .I3(n28939), .O(n2319)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_27_lut (.I0(GND_net), .I1(n3034), .I2(VCC_net), 
            .I3(n28723), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_9 (.CI(n28939), .I0(n2252), .I1(VCC_net), 
            .CO(n28940));
    SB_CARRY rem_4_add_2055_27 (.CI(n28723), .I0(n3034), .I1(VCC_net), 
            .CO(n28724));
    SB_LUT4 div_46_mux_3_i3_3_lut (.I0(encoder0_position[2]), .I1(n23_adj_4713), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n1064));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13387_3_lut (.I0(\data_in_frame[24] [0]), .I1(rx_data[0]), 
            .I2(n36526), .I3(GND_net), .O(n18126));   // verilog/coms.v(127[12] 295[6])
    defparam i13387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1722_i33_2_lut (.I0(n2625), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5168));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2355_9_lut (.I0(GND_net), .I1(n2715), .I2(n94), .I3(n28495), 
            .O(n6233)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1722_i35_2_lut (.I0(n2624), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5170));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_2055_26_lut (.I0(GND_net), .I1(n3035), .I2(VCC_net), 
            .I3(n28722), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1389_3_lut (.I0(n2044), .I1(n2111), .I2(n2075_adj_5028), 
            .I3(GND_net), .O(n2143));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1389_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2355_9 (.CI(n28495), .I0(n2715), .I1(n94), .CO(n28496));
    SB_LUT4 rem_4_add_648_7_lut (.I0(n986), .I1(n953), .I2(VCC_net), .I3(n27919), 
            .O(n1052)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_7_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_2355_8_lut (.I0(GND_net), .I1(n2716), .I2(n95), .I3(n28494), 
            .O(n6234)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1722_i27_2_lut (.I0(n2628), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5165));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i27_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2355_8 (.CI(n28494), .I0(n2716), .I1(n95), .CO(n28495));
    SB_LUT4 div_46_LessThan_1722_i29_2_lut (.I0(n2627), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5166));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13397_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n4593), .I3(GND_net), .O(n18136));   // verilog/coms.v(127[12] 295[6])
    defparam i13397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2355_7_lut (.I0(GND_net), .I1(n2717), .I2(n96), .I3(n28493), 
            .O(n6235)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1388_3_lut (.I0(n2043), .I1(n2110), .I2(n2075_adj_5028), 
            .I3(GND_net), .O(n2142));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1388_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13396_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n4593), .I3(GND_net), .O(n18135));   // verilog/coms.v(127[12] 295[6])
    defparam i13396_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_648_6_lut (.I0(GND_net), .I1(n954), .I2(GND_net), 
            .I3(n27918), .O(n1021)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1397_3_lut (.I0(n2052), .I1(n2119), .I2(n2075_adj_5028), 
            .I3(GND_net), .O(n2151));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1397_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13395_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n4593), .I3(GND_net), .O(n18134));   // verilog/coms.v(127[12] 295[6])
    defparam i13395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1722_i23_2_lut (.I0(n2630), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5163));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i25_2_lut (.I0(n2629), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5164));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i25_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2355_7 (.CI(n28493), .I0(n2717), .I1(n96), .CO(n28494));
    SB_LUT4 i13394_3_lut (.I0(\data_in_frame[24] [7]), .I1(rx_data[7]), 
            .I2(n36526), .I3(GND_net), .O(n18133));   // verilog/coms.v(127[12] 295[6])
    defparam i13394_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13405_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n4593), .I3(GND_net), .O(n18144));   // verilog/coms.v(127[12] 295[6])
    defparam i13405_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2355_6_lut (.I0(GND_net), .I1(n2718), .I2(n97), .I3(n28492), 
            .O(n6236)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13404_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n4593), .I3(GND_net), .O(n18143));   // verilog/coms.v(127[12] 295[6])
    defparam i13404_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_648_6 (.CI(n27918), .I0(n954), .I1(GND_net), .CO(n27919));
    SB_LUT4 i13415_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n4593), .I3(GND_net), .O(n18154));   // verilog/coms.v(127[12] 295[6])
    defparam i13415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13414_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n4593), .I3(GND_net), .O(n18153));   // verilog/coms.v(127[12] 295[6])
    defparam i13414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13413_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n4593), .I3(GND_net), .O(n18152));   // verilog/coms.v(127[12] 295[6])
    defparam i13413_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2355_6 (.CI(n28492), .I0(n2718), .I1(n97), .CO(n28493));
    SB_LUT4 rem_4_i1396_rep_68_3_lut (.I0(n2051), .I1(n2118), .I2(n2075_adj_5028), 
            .I3(GND_net), .O(n2150));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1396_rep_68_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2355_5_lut (.I0(GND_net), .I1(n2719), .I2(n98), .I3(n28491), 
            .O(n6237)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1722_i11_2_lut (.I0(n2636), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_5153));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i11_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i39_2_lut (.I0(n2622), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5172));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13417_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n4593), .I3(GND_net), .O(n18156));   // verilog/coms.v(127[12] 295[6])
    defparam i13417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13416_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n4593), .I3(GND_net), .O(n18155));   // verilog/coms.v(127[12] 295[6])
    defparam i13416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13419_3_lut (.I0(encoder0_position[2]), .I1(n3014), .I2(count_enable), 
            .I3(GND_net), .O(n18158));   // quad.v(35[10] 41[6])
    defparam i13419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1722_i37_2_lut (.I0(n2623), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5171));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13418_3_lut (.I0(encoder0_position[1]), .I1(n3015), .I2(count_enable), 
            .I3(GND_net), .O(n18157));   // quad.v(35[10] 41[6])
    defparam i13418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13421_3_lut (.I0(encoder0_position[4]), .I1(n3012), .I2(count_enable), 
            .I3(GND_net), .O(n18160));   // quad.v(35[10] 41[6])
    defparam i13421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13420_3_lut (.I0(encoder0_position[3]), .I1(n3013), .I2(count_enable), 
            .I3(GND_net), .O(n18159));   // quad.v(35[10] 41[6])
    defparam i13420_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2355_5 (.CI(n28491), .I0(n2719), .I1(n98), .CO(n28492));
    SB_LUT4 i13423_3_lut (.I0(encoder0_position[6]), .I1(n3010), .I2(count_enable), 
            .I3(GND_net), .O(n18162));   // quad.v(35[10] 41[6])
    defparam i13423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1395_3_lut (.I0(n2050), .I1(n2117), .I2(n2075_adj_5028), 
            .I3(GND_net), .O(n2149));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1395_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_1519_8_lut (.I0(GND_net), .I1(n2253), .I2(VCC_net), 
            .I3(n28938), .O(n2320)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_8 (.CI(n28938), .I0(n2253), .I1(VCC_net), 
            .CO(n28939));
    SB_LUT4 rem_4_i1394_3_lut (.I0(n2049), .I1(n2116), .I2(n2075_adj_5028), 
            .I3(GND_net), .O(n2148));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1394_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13422_3_lut (.I0(encoder0_position[5]), .I1(n3011), .I2(count_enable), 
            .I3(GND_net), .O(n18161));   // quad.v(35[10] 41[6])
    defparam i13422_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2055_26 (.CI(n28722), .I0(n3035), .I1(VCC_net), 
            .CO(n28723));
    SB_LUT4 rem_4_add_1519_7_lut (.I0(GND_net), .I1(n2254), .I2(GND_net), 
            .I3(n28937), .O(n2321)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13425_3_lut (.I0(encoder0_position[8]), .I1(n3008), .I2(count_enable), 
            .I3(GND_net), .O(n18164));   // quad.v(35[10] 41[6])
    defparam i13425_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13424_3_lut (.I0(encoder0_position[7]), .I1(n3009), .I2(count_enable), 
            .I3(GND_net), .O(n18163));   // quad.v(35[10] 41[6])
    defparam i13424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1722_i15_2_lut (.I0(n2634), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5157));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i17_2_lut (.I0(n2633), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5159));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1722_i19_2_lut (.I0(n2632), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5160));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_2055_25_lut (.I0(GND_net), .I1(n3036), .I2(VCC_net), 
            .I3(n28721), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_25_lut.LUT_INIT = 16'hC33C;
    SB_IO PIN_8_pad (.PACKAGE_PIN(PIN_8), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_8_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_8_pad.PIN_TYPE = 6'b011001;
    defparam PIN_8_pad.PULLUP = 1'b0;
    defparam PIN_8_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_8_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_7_pad (.PACKAGE_PIN(PIN_7), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_7_c_0)) /* synthesis IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_7_pad.PIN_TYPE = 6'b000001;
    defparam PIN_7_pad.PULLUP = 1'b0;
    defparam PIN_7_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_7_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 div_46_LessThan_1722_i31_2_lut (.I0(n2626), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5167));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2355_4_lut (.I0(GND_net), .I1(n2720), .I2(n99), .I3(n28490), 
            .O(n6238)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2355_4 (.CI(n28490), .I0(n2720), .I1(n99), .CO(n28491));
    SB_CARRY rem_4_add_1519_7 (.CI(n28937), .I0(n2254), .I1(GND_net), 
            .CO(n28938));
    SB_LUT4 rem_4_i1401_3_lut (.I0(n2056), .I1(n2123), .I2(n2075_adj_5028), 
            .I3(GND_net), .O(n2155));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1401_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_2055_25 (.CI(n28721), .I0(n3036), .I1(VCC_net), 
            .CO(n28722));
    SB_LUT4 rem_4_add_1519_6_lut (.I0(GND_net), .I1(n2255), .I2(GND_net), 
            .I3(n28936), .O(n2322)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_24_lut (.I0(GND_net), .I1(n3037), .I2(VCC_net), 
            .I3(n28720), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1722_i13_2_lut (.I0(n2635), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5155));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2355_3_lut (.I0(GND_net), .I1(n1065), .I2(n558), .I3(n28489), 
            .O(n6239)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2355_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2355_3 (.CI(n28489), .I0(n1065), .I1(n558), .CO(n28490));
    SB_CARRY add_2355_2 (.CI(VCC_net), .I0(n1066), .I1(VCC_net), .CO(n28489));
    SB_LUT4 div_46_LessThan_1722_i21_2_lut (.I0(n2631), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5162));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1724_1_lut (.I0(n2642), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2643));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1724_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1393_3_lut (.I0(n2048), .I1(n2115), .I2(n2075_adj_5028), 
            .I3(GND_net), .O(n2147));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1393_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2354_23_lut (.I0(GND_net), .I1(n2618), .I2(n79), .I3(n28488), 
            .O(n6193)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2354_22_lut (.I0(GND_net), .I1(n2619), .I2(n80), .I3(n28487), 
            .O(n6194)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1400_3_lut (.I0(n2055), .I1(n2122), .I2(n2075_adj_5028), 
            .I3(GND_net), .O(n2154));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33990_4_lut (.I0(n31_adj_5167), .I1(n19_adj_5160), .I2(n17_adj_5159), 
            .I3(n15_adj_5157), .O(n40836));
    defparam i33990_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 rem_4_i1331_3_lut (.I0(n1954), .I1(n2021), .I2(n1976_adj_4779), 
            .I3(GND_net), .O(n2053));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1331_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1329_3_lut (.I0(n1952), .I1(n2019), .I2(n1976_adj_4779), 
            .I3(GND_net), .O(n2051));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1329_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2354_22 (.CI(n28487), .I0(n2619), .I1(n80), .CO(n28488));
    SB_LUT4 add_2354_21_lut (.I0(GND_net), .I1(n2620), .I2(n81), .I3(n28486), 
            .O(n6195)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1722_i34_3_lut (.I0(n16_adj_5158), .I1(n83), 
            .I2(n39_adj_5172), .I3(GND_net), .O(n34_adj_5169));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34724_4_lut (.I0(n13_adj_5155), .I1(n11_adj_5153), .I2(n2637), 
            .I3(n98), .O(n41571));
    defparam i34724_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i35254_4_lut (.I0(n19_adj_5160), .I1(n17_adj_5159), .I2(n15_adj_5157), 
            .I3(n41571), .O(n42101));
    defparam i35254_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 rem_4_i1323_3_lut (.I0(n1946), .I1(n2013), .I2(n1976_adj_4779), 
            .I3(GND_net), .O(n2045));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1323_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13436_3_lut (.I0(encoder0_position[19]), .I1(n2997), .I2(count_enable), 
            .I3(GND_net), .O(n18175));   // quad.v(35[10] 41[6])
    defparam i13436_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35252_4_lut (.I0(n25_adj_5164), .I1(n23_adj_5163), .I2(n21_adj_5162), 
            .I3(n42101), .O(n42099));
    defparam i35252_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i33996_4_lut (.I0(n31_adj_5167), .I1(n29_adj_5166), .I2(n27_adj_5165), 
            .I3(n42099), .O(n40842));
    defparam i33996_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2354_21 (.CI(n28486), .I0(n2620), .I1(n81), .CO(n28487));
    SB_LUT4 i13435_3_lut (.I0(encoder0_position[18]), .I1(n2998), .I2(count_enable), 
            .I3(GND_net), .O(n18174));   // quad.v(35[10] 41[6])
    defparam i13435_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13434_3_lut (.I0(encoder0_position[17]), .I1(n2999), .I2(count_enable), 
            .I3(GND_net), .O(n18173));   // quad.v(35[10] 41[6])
    defparam i13434_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13433_3_lut (.I0(encoder0_position[16]), .I1(n3000), .I2(count_enable), 
            .I3(GND_net), .O(n18172));   // quad.v(35[10] 41[6])
    defparam i13433_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13432_3_lut (.I0(encoder0_position[15]), .I1(n3001), .I2(count_enable), 
            .I3(GND_net), .O(n18171));   // quad.v(35[10] 41[6])
    defparam i13432_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1519_6 (.CI(n28936), .I0(n2255), .I1(GND_net), 
            .CO(n28937));
    SB_CARRY rem_4_add_2055_24 (.CI(n28720), .I0(n3037), .I1(VCC_net), 
            .CO(n28721));
    SB_LUT4 add_2354_20_lut (.I0(GND_net), .I1(n2621), .I2(n82), .I3(n28485), 
            .O(n6196)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13431_3_lut (.I0(encoder0_position[14]), .I1(n3002), .I2(count_enable), 
            .I3(GND_net), .O(n18170));   // quad.v(35[10] 41[6])
    defparam i13431_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13430_3_lut (.I0(encoder0_position[13]), .I1(n3003), .I2(count_enable), 
            .I3(GND_net), .O(n18169));   // quad.v(35[10] 41[6])
    defparam i13430_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13429_3_lut (.I0(encoder0_position[12]), .I1(n3004), .I2(count_enable), 
            .I3(GND_net), .O(n18168));   // quad.v(35[10] 41[6])
    defparam i13429_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13428_3_lut (.I0(encoder0_position[11]), .I1(n3005), .I2(count_enable), 
            .I3(GND_net), .O(n18167));   // quad.v(35[10] 41[6])
    defparam i13428_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35470_4_lut (.I0(n37_adj_5171), .I1(n35_adj_5170), .I2(n33_adj_5168), 
            .I3(n40842), .O(n42317));
    defparam i35470_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13444_3_lut (.I0(encoder1_position[3]), .I1(n2963), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18183));   // quad.v(35[10] 41[6])
    defparam i13444_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2354_20 (.CI(n28485), .I0(n2621), .I1(n82), .CO(n28486));
    SB_LUT4 i13443_3_lut (.I0(encoder1_position[2]), .I1(n2964), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18182));   // quad.v(35[10] 41[6])
    defparam i13443_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13454_3_lut (.I0(encoder1_position[13]), .I1(n2953), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18193));   // quad.v(35[10] 41[6])
    defparam i13454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13453_3_lut (.I0(encoder1_position[12]), .I1(n2954), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18192));   // quad.v(35[10] 41[6])
    defparam i13453_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13452_3_lut (.I0(encoder1_position[11]), .I1(n2955), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18191));   // quad.v(35[10] 41[6])
    defparam i13452_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1324_3_lut (.I0(n1947), .I1(n2014), .I2(n1976_adj_4779), 
            .I3(GND_net), .O(n2046));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1324_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2354_19_lut (.I0(GND_net), .I1(n2622), .I2(n83), .I3(n28484), 
            .O(n6197)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13456_3_lut (.I0(encoder1_position[15]), .I1(n2951), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18195));   // quad.v(35[10] 41[6])
    defparam i13456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13455_3_lut (.I0(encoder1_position[14]), .I1(n2952), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18194));   // quad.v(35[10] 41[6])
    defparam i13455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13458_3_lut (.I0(encoder1_position[17]), .I1(n2949), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18197));   // quad.v(35[10] 41[6])
    defparam i13458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13457_3_lut (.I0(encoder1_position[16]), .I1(n2950), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18196));   // quad.v(35[10] 41[6])
    defparam i13457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35713_3_lut (.I0(n10_adj_5152), .I1(n90), .I2(n25_adj_5164), 
            .I3(GND_net), .O(n42560));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35713_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12_3_lut (.I0(bit_ctr[18]), .I1(n40713), .I2(n4483), .I3(GND_net), 
            .O(n33647));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 rem_4_i1321_3_lut (.I0(n1944), .I1(n2011), .I2(n1976_adj_4779), 
            .I3(GND_net), .O(n2043));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1321_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2354_19 (.CI(n28484), .I0(n2622), .I1(n83), .CO(n28485));
    SB_LUT4 i13460_3_lut (.I0(encoder1_position[19]), .I1(n2947), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18199));   // quad.v(35[10] 41[6])
    defparam i13460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13459_3_lut (.I0(encoder1_position[18]), .I1(n2948), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18198));   // quad.v(35[10] 41[6])
    defparam i13459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13462_3_lut (.I0(encoder1_position[21]), .I1(n2945), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18201));   // quad.v(35[10] 41[6])
    defparam i13462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13461_3_lut (.I0(encoder1_position[20]), .I1(n2946), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18200));   // quad.v(35[10] 41[6])
    defparam i13461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13464_3_lut (.I0(encoder1_position[23]), .I1(n2943), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18203));   // quad.v(35[10] 41[6])
    defparam i13464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2354_18_lut (.I0(GND_net), .I1(n2623), .I2(n84), .I3(n28483), 
            .O(n6198)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13463_3_lut (.I0(encoder1_position[22]), .I1(n2944), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18202));   // quad.v(35[10] 41[6])
    defparam i13463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13403_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n4593), .I3(GND_net), .O(n18142));   // verilog/coms.v(127[12] 295[6])
    defparam i13403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13402_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n4593), .I3(GND_net), .O(n18141));   // verilog/coms.v(127[12] 295[6])
    defparam i13402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13401_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n4593), .I3(GND_net), .O(n18140));   // verilog/coms.v(127[12] 295[6])
    defparam i13401_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13400_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n4593), .I3(GND_net), .O(n18139));   // verilog/coms.v(127[12] 295[6])
    defparam i13400_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13399_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n4593), .I3(GND_net), .O(n18138));   // verilog/coms.v(127[12] 295[6])
    defparam i13399_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13398_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n4593), .I3(GND_net), .O(n18137));   // verilog/coms.v(127[12] 295[6])
    defparam i13398_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35714_3_lut (.I0(n42560), .I1(n89), .I2(n27_adj_5165), .I3(GND_net), 
            .O(n42561));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35714_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_2354_18 (.CI(n28483), .I0(n2623), .I1(n84), .CO(n28484));
    SB_LUT4 i12_3_lut_adj_1731 (.I0(n40745), .I1(byte_transmit_counter[0]), 
            .I2(n24918), .I3(GND_net), .O(n34409));   // verilog/coms.v(127[12] 295[6])
    defparam i12_3_lut_adj_1731.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_3_lut_adj_1732 (.I0(n40703), .I1(bit_ctr[13]), .I2(n4483), 
            .I3(GND_net), .O(n33621));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1732.LUT_INIT = 16'hcaca;
    SB_LUT4 i34708_4_lut (.I0(n27_adj_5165), .I1(n25_adj_5164), .I2(n23_adj_5163), 
            .I3(n40856), .O(n41555));
    defparam i34708_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_46_LessThan_1722_i20_3_lut (.I0(n12_adj_5154), .I1(n91), 
            .I2(n23_adj_5163), .I3(GND_net), .O(n20_adj_5161));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i20_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_2354_17_lut (.I0(GND_net), .I1(n2624), .I2(n85), .I3(n28482), 
            .O(n6199)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13412_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n4593), .I3(GND_net), .O(n18151));   // verilog/coms.v(127[12] 295[6])
    defparam i13412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13411_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n4593), .I3(GND_net), .O(n18150));   // verilog/coms.v(127[12] 295[6])
    defparam i13411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13410_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n4593), .I3(GND_net), .O(n18149));   // verilog/coms.v(127[12] 295[6])
    defparam i13410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13409_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n4593), .I3(GND_net), .O(n18148));   // verilog/coms.v(127[12] 295[6])
    defparam i13409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13408_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n4593), .I3(GND_net), .O(n18147));   // verilog/coms.v(127[12] 295[6])
    defparam i13408_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35604_3_lut (.I0(n42561), .I1(n88), .I2(n29_adj_5166), .I3(GND_net), 
            .O(n42451));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35604_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13407_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n4593), .I3(GND_net), .O(n18146));   // verilog/coms.v(127[12] 295[6])
    defparam i13407_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2354_17 (.CI(n28482), .I0(n2624), .I1(n85), .CO(n28483));
    SB_LUT4 i13406_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n4593), .I3(GND_net), .O(n18145));   // verilog/coms.v(127[12] 295[6])
    defparam i13406_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_3_lut_adj_1733 (.I0(bit_ctr[11]), .I1(n40700), .I2(n4483), 
            .I3(GND_net), .O(n33601));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1733.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1722_i8_4_lut (.I0(n1064), .I1(n99), .I2(n2638), 
            .I3(n558), .O(n8_adj_5151));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i8_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 add_2354_16_lut (.I0(GND_net), .I1(n2625), .I2(n86), .I3(n28481), 
            .O(n6200)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1734 (.I0(color[9]), .I1(n25736), .I2(n25734), 
            .I3(GND_net), .O(n18215));
    defparam i1_3_lut_adj_1734.LUT_INIT = 16'hecec;
    SB_LUT4 i36743_4_lut (.I0(r_SM_Main[2]), .I1(n40689), .I2(n40690), 
            .I3(r_SM_Main[1]), .O(n24794));
    defparam i36743_4_lut.LUT_INIT = 16'h0511;
    SB_LUT4 rem_4_add_1519_5_lut (.I0(GND_net), .I1(n2256), .I2(VCC_net), 
            .I3(n28935), .O(n2323)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35711_3_lut (.I0(n8_adj_5151), .I1(n87), .I2(n31_adj_5167), 
            .I3(GND_net), .O(n42558));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35711_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_2354_16 (.CI(n28481), .I0(n2625), .I1(n86), .CO(n28482));
    SB_LUT4 i13474_3_lut (.I0(quadA_debounced), .I1(reg_B[1]), .I2(n36518), 
            .I3(GND_net), .O(n18213));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13474_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21117_3_lut (.I0(bit_ctr[0]), .I1(n40616), .I2(n4483), .I3(GND_net), 
            .O(n18212));
    defparam i21117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_2354_15_lut (.I0(GND_net), .I1(n2626), .I2(n87), .I3(n28480), 
            .O(n6201)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1735 (.I0(color[10]), .I1(n25736), .I2(n25734), 
            .I3(GND_net), .O(n18222));
    defparam i1_3_lut_adj_1735.LUT_INIT = 16'hecec;
    SB_LUT4 i12_3_lut_adj_1736 (.I0(bit_ctr[10]), .I1(n40699), .I2(n4483), 
            .I3(GND_net), .O(n33595));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1736.LUT_INIT = 16'hacac;
    SB_LUT4 i13491_3_lut (.I0(setpoint[1]), .I1(n4387), .I2(n37622), .I3(GND_net), 
            .O(n18230));   // verilog/coms.v(127[12] 295[6])
    defparam i13491_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_2354_15 (.CI(n28480), .I0(n2626), .I1(n87), .CO(n28481));
    SB_LUT4 i13490_3_lut (.I0(quadA_debounced_adj_4678), .I1(reg_B_adj_5411[1]), 
            .I2(n36342), .I3(GND_net), .O(n18229));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i13490_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13501_3_lut (.I0(setpoint[11]), .I1(n4397), .I2(n37622), 
            .I3(GND_net), .O(n18240));   // verilog/coms.v(127[12] 295[6])
    defparam i13501_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13500_3_lut (.I0(setpoint[10]), .I1(n4396), .I2(n37622), 
            .I3(GND_net), .O(n18239));   // verilog/coms.v(127[12] 295[6])
    defparam i13500_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35712_3_lut (.I0(n42558), .I1(n86), .I2(n33_adj_5168), .I3(GND_net), 
            .O(n42559));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35712_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33978_4_lut (.I0(n37_adj_5171), .I1(n35_adj_5170), .I2(n33_adj_5168), 
            .I3(n40836), .O(n40824));
    defparam i33978_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35928_4_lut (.I0(n34_adj_5169), .I1(n14_adj_5156), .I2(n39_adj_5172), 
            .I3(n40815), .O(n42775));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35928_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 rem_4_i1330_3_lut (.I0(n1953), .I1(n2020), .I2(n1976_adj_4779), 
            .I3(GND_net), .O(n2052));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1330_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35606_3_lut (.I0(n42559), .I1(n85), .I2(n35_adj_5170), .I3(GND_net), 
            .O(n42453));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35606_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13499_3_lut (.I0(setpoint[9]), .I1(n4395), .I2(n37622), .I3(GND_net), 
            .O(n18238));   // verilog/coms.v(127[12] 295[6])
    defparam i13499_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36024_4_lut (.I0(n42453), .I1(n42775), .I2(n39_adj_5172), 
            .I3(n40824), .O(n42871));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36024_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36025_3_lut (.I0(n42871), .I1(n82), .I2(n41_adj_5173), .I3(GND_net), 
            .O(n42872));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36025_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35993_3_lut (.I0(n42872), .I1(n81), .I2(n43_adj_5174), .I3(GND_net), 
            .O(n42840));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35993_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35936_4_lut (.I0(n43_adj_5174), .I1(n41_adj_5173), .I2(n39_adj_5172), 
            .I3(n42317), .O(n42783));
    defparam i35936_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13427_3_lut (.I0(encoder0_position[10]), .I1(n3006), .I2(count_enable), 
            .I3(GND_net), .O(n18166));   // quad.v(35[10] 41[6])
    defparam i13427_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35609_4_lut (.I0(n42451), .I1(n20_adj_5161), .I2(n29_adj_5166), 
            .I3(n41555), .O(n42456));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35609_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i13426_3_lut (.I0(encoder0_position[9]), .I1(n3007), .I2(count_enable), 
            .I3(GND_net), .O(n18165));   // quad.v(35[10] 41[6])
    defparam i13426_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35977_3_lut (.I0(n42840), .I1(n80), .I2(n45_adj_5176), .I3(GND_net), 
            .O(n44_adj_5175));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35977_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35611_4_lut (.I0(n44_adj_5175), .I1(n42456), .I2(n45_adj_5176), 
            .I3(n42783), .O(n42458));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35611_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1737 (.I0(n42458), .I1(n15910), .I2(n79), .I3(n2618), 
            .O(n2642));
    defparam i1_4_lut_adj_1737.LUT_INIT = 16'hceef;
    SB_LUT4 rem_4_i1327_3_lut (.I0(n1950), .I1(n2017), .I2(n1976_adj_4779), 
            .I3(GND_net), .O(n2049));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1327_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13155_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n13302), 
            .I3(GND_net), .O(n17894));   // verilog/coms.v(127[12] 295[6])
    defparam i13155_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13156_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n13302), 
            .I3(GND_net), .O(n17895));   // verilog/coms.v(127[12] 295[6])
    defparam i13156_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13157_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n13302), 
            .I3(GND_net), .O(n17896));   // verilog/coms.v(127[12] 295[6])
    defparam i13157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1665_i41_2_lut (.I0(n2537), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5150));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13503_3_lut (.I0(setpoint[13]), .I1(n4399), .I2(n37622), 
            .I3(GND_net), .O(n18242));   // verilog/coms.v(127[12] 295[6])
    defparam i13503_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1665_i37_2_lut (.I0(n2539), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5148));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i35_2_lut (.I0(n2540), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5146));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i4_3_lut (.I0(encoder0_position[3]), .I1(n22_adj_4714), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n1063));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1665_i39_2_lut (.I0(n2538), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5149));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i1326_3_lut (.I0(n1949), .I1(n2016), .I2(n1976_adj_4779), 
            .I3(GND_net), .O(n2048));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1326_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1328_3_lut (.I0(n1951), .I1(n2018), .I2(n1976_adj_4779), 
            .I3(GND_net), .O(n2050));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1328_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1665_i29_2_lut (.I0(n2543), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5143));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i31_2_lut (.I0(n2542), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5144));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i1325_3_lut (.I0(n1948), .I1(n2015), .I2(n1976_adj_4779), 
            .I3(GND_net), .O(n2047));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1325_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1665_i23_2_lut (.I0(n2546), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5140));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i25_2_lut (.I0(n2545), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5141));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i1333_3_lut (.I0(n1956), .I1(n2023), .I2(n1976_adj_4779), 
            .I3(GND_net), .O(n2055));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1333_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1665_i27_2_lut (.I0(n2544), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5142));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i27_2_lut.LUT_INIT = 16'h9999;
    SB_IO PIN_13_pad (.PACKAGE_PIN(PIN_13), .OUTPUT_ENABLE(VCC_net), .D_IN_0(PIN_13_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_13_pad.PIN_TYPE = 6'b000001;
    defparam PIN_13_pad.PULLUP = 1'b0;
    defparam PIN_13_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_13_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO PIN_21_pad (.PACKAGE_PIN(PIN_21), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(PIN_21_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam PIN_21_pad.PIN_TYPE = 6'b011001;
    defparam PIN_21_pad.PULLUP = 1'b0;
    defparam PIN_21_pad.NEG_TRIGGER = 1'b0;
    defparam PIN_21_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 rem_4_i1332_3_lut (.I0(n1955), .I1(n2022), .I2(n1976_adj_4779), 
            .I3(GND_net), .O(n2054));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1332_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1665_i17_2_lut (.I0(n2549), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5135));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i19_2_lut (.I0(n2548), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5137));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i21_2_lut (.I0(n2547), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5138));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i33_2_lut (.I0(n2541), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5145));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12_3_lut_adj_1738 (.I0(bit_ctr[17]), .I1(n40712), .I2(n4483), 
            .I3(GND_net), .O(n33645));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1738.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1739 (.I0(bit_ctr[5]), .I1(n40711), .I2(n4483), 
            .I3(GND_net), .O(n33643));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1739.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1740 (.I0(bit_ctr[4]), .I1(n40710), .I2(n4483), 
            .I3(GND_net), .O(n33641));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1740.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1741 (.I0(bit_ctr[16]), .I1(n40709), .I2(n4483), 
            .I3(GND_net), .O(n33639));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1741.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1742 (.I0(bit_ctr[15]), .I1(n40708), .I2(n4483), 
            .I3(GND_net), .O(n33635));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1742.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1743 (.I0(bit_ctr[27]), .I1(n40722), .I2(n4483), 
            .I3(GND_net), .O(n33665));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1743.LUT_INIT = 16'hacac;
    SB_LUT4 add_2354_14_lut (.I0(GND_net), .I1(n2627), .I2(n88), .I3(n28479), 
            .O(n6202)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1322_3_lut (.I0(n1945), .I1(n2012), .I2(n1976_adj_4779), 
            .I3(GND_net), .O(n2044));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1322_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1665_i13_2_lut (.I0(n2551), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_5131));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i13_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1665_i15_2_lut (.I0(n2550), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5133));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i1335_3_lut (.I0(n1958), .I1(n2025), .I2(n1976_adj_4779), 
            .I3(GND_net), .O(n2057));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1335_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1334_3_lut (.I0(n1957), .I1(n2024), .I2(n1976_adj_4779), 
            .I3(GND_net), .O(n2056));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1667_1_lut (.I0(n2558), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2559));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1667_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34055_4_lut (.I0(n33_adj_5145), .I1(n21_adj_5138), .I2(n19_adj_5137), 
            .I3(n17_adj_5135), .O(n40901));
    defparam i34055_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i12_3_lut_adj_1744 (.I0(bit_ctr[26]), .I1(n40721), .I2(n4483), 
            .I3(GND_net), .O(n33663));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1744.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1745 (.I0(bit_ctr[25]), .I1(n40720), .I2(n4483), 
            .I3(GND_net), .O(n33661));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1745.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1746 (.I0(bit_ctr[24]), .I1(n40719), .I2(n4483), 
            .I3(GND_net), .O(n33659));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1746.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1747 (.I0(bit_ctr[23]), .I1(n40718), .I2(n4483), 
            .I3(GND_net), .O(n33657));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1747.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1748 (.I0(bit_ctr[22]), .I1(n40717), .I2(n4483), 
            .I3(GND_net), .O(n33655));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1748.LUT_INIT = 16'hacac;
    SB_LUT4 i34766_4_lut (.I0(n15_adj_5133), .I1(n13_adj_5131), .I2(n2552), 
            .I3(n98), .O(n41613));
    defparam i34766_4_lut.LUT_INIT = 16'hfeef;
    SB_CARRY add_2354_14 (.CI(n28479), .I0(n2627), .I1(n88), .CO(n28480));
    SB_LUT4 i35270_4_lut (.I0(n21_adj_5138), .I1(n19_adj_5137), .I2(n17_adj_5135), 
            .I3(n41613), .O(n42117));
    defparam i35270_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35268_4_lut (.I0(n27_adj_5142), .I1(n25_adj_5141), .I2(n23_adj_5140), 
            .I3(n42117), .O(n42115));
    defparam i35268_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34059_4_lut (.I0(n33_adj_5145), .I1(n31_adj_5144), .I2(n29_adj_5143), 
            .I3(n42115), .O(n40905));
    defparam i34059_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1665_i10_4_lut (.I0(n1063), .I1(n99), .I2(n2553), 
            .I3(n558), .O(n10_adj_5129));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i10_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 add_2354_13_lut (.I0(GND_net), .I1(n2628), .I2(n89), .I3(n28478), 
            .O(n6203)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35717_3_lut (.I0(n10_adj_5129), .I1(n87), .I2(n33_adj_5145), 
            .I3(GND_net), .O(n42564));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35717_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35718_3_lut (.I0(n42564), .I1(n86), .I2(n35_adj_5146), .I3(GND_net), 
            .O(n42565));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35718_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i12_3_lut_adj_1749 (.I0(bit_ctr[21]), .I1(n40716), .I2(n4483), 
            .I3(GND_net), .O(n33653));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1749.LUT_INIT = 16'hacac;
    SB_LUT4 i12758_4_lut (.I0(n17505), .I1(r_Clock_Count_adj_5401[4]), .I2(n317), 
            .I3(r_SM_Main_adj_5400[2]), .O(n17497));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12758_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i12761_4_lut (.I0(n17505), .I1(r_Clock_Count_adj_5401[3]), .I2(n318), 
            .I3(r_SM_Main_adj_5400[2]), .O(n17500));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12761_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 div_46_LessThan_1665_i36_3_lut (.I0(n18_adj_5136), .I1(n83), 
            .I2(n41_adj_5150), .I3(GND_net), .O(n36_adj_5147));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34045_4_lut (.I0(n39_adj_5149), .I1(n37_adj_5148), .I2(n35_adj_5146), 
            .I3(n40901), .O(n40891));
    defparam i34045_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35947_4_lut (.I0(n36_adj_5147), .I1(n16_adj_5134), .I2(n41_adj_5150), 
            .I3(n40887), .O(n42794));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35947_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35600_3_lut (.I0(n42565), .I1(n85), .I2(n37_adj_5148), .I3(GND_net), 
            .O(n42447));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35600_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1665_i22_3_lut (.I0(n14_adj_5132), .I1(n91), 
            .I2(n25_adj_5141), .I3(GND_net), .O(n22_adj_5139));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i22_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4932));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4931));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4930));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35945_4_lut (.I0(n22_adj_5139), .I1(n12_adj_5130), .I2(n25_adj_5141), 
            .I3(n40928), .O(n42792));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35945_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35946_3_lut (.I0(n42792), .I1(n90), .I2(n27_adj_5142), .I3(GND_net), 
            .O(n42793));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35946_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35859_3_lut (.I0(n42793), .I1(n89), .I2(n29_adj_5143), .I3(GND_net), 
            .O(n42706));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35859_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35486_4_lut (.I0(n39_adj_5149), .I1(n37_adj_5148), .I2(n35_adj_5146), 
            .I3(n40905), .O(n42333));
    defparam i35486_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36022_4_lut (.I0(n42447), .I1(n42794), .I2(n41_adj_5150), 
            .I3(n40891), .O(n42869));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36022_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35789_3_lut (.I0(n42706), .I1(n88), .I2(n31_adj_5144), .I3(GND_net), 
            .O(n42636));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35789_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36036_4_lut (.I0(n42636), .I1(n42869), .I2(n41_adj_5150), 
            .I3(n42333), .O(n42883));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36036_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36037_3_lut (.I0(n42883), .I1(n82), .I2(n2536), .I3(GND_net), 
            .O(n42884));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36037_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i36033_3_lut (.I0(n42884), .I1(n81), .I2(n2535), .I3(GND_net), 
            .O(n42880));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36033_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1750 (.I0(n42880), .I1(n15904), .I2(n80), .I3(n2534), 
            .O(n2558));
    defparam i1_4_lut_adj_1750.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4929));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4928));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4927));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4926));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4925));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4924));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1751 (.I0(n2056), .I1(n2057), .I2(n2058), .I3(GND_net), 
            .O(n36038));
    defparam i1_3_lut_adj_1751.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1752 (.I0(n2044), .I1(n2054), .I2(n36038), .I3(n2055), 
            .O(n16_adj_5235));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i3_4_lut_adj_1752.LUT_INIT = 16'heaaa;
    SB_LUT4 i13158_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n13302), 
            .I3(GND_net), .O(n17897));   // verilog/coms.v(127[12] 295[6])
    defparam i13158_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13502_3_lut (.I0(setpoint[12]), .I1(n4398), .I2(n37622), 
            .I3(GND_net), .O(n18241));   // verilog/coms.v(127[12] 295[6])
    defparam i13502_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4923));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4922));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4921));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1124_3_lut (.I0(n1651_adj_4818), .I1(n1718), .I2(n1679), 
            .I3(GND_net), .O(n1750));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1124_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1126_3_lut (.I0(n1653_adj_4820), .I1(n1720), .I2(n1679), 
            .I3(GND_net), .O(n1752));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1129_3_lut (.I0(n1656), .I1(n1723), .I2(n1679), .I3(GND_net), 
            .O(n1755_adj_4808));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1123_3_lut (.I0(n1650_adj_4817), .I1(n1717), .I2(n1679), 
            .I3(GND_net), .O(n1749));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1123_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1128_3_lut (.I0(n1655), .I1(n1722), .I2(n1679), .I3(GND_net), 
            .O(n1754_adj_4807));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i19_3_lut (.I0(communication_counter[18]), .I1(n15_adj_4794), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1758_adj_4811));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1131_3_lut (.I0(n1658), .I1(n1725), .I2(n1679), .I3(GND_net), 
            .O(n1757_adj_4810));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1130_3_lut (.I0(n1657), .I1(n1724), .I2(n1679), .I3(GND_net), 
            .O(n1756_adj_4809));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1127_3_lut (.I0(n1654), .I1(n1721), .I2(n1679), .I3(GND_net), 
            .O(n1753));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1125_3_lut (.I0(n1652_adj_4819), .I1(n1719), .I2(n1679), 
            .I3(GND_net), .O(n1751));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1056_3_lut (.I0(n1551), .I1(n1618), .I2(n1580), .I3(GND_net), 
            .O(n1650_adj_4817));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1056_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i20_3_lut (.I0(communication_counter[19]), .I1(n14_adj_4795), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1658));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1063_3_lut (.I0(n1558), .I1(n1625), .I2(n1580), .I3(GND_net), 
            .O(n1657));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1606_i39_2_lut (.I0(n2451), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5126));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i9_4_lut_adj_1753 (.I0(n2047), .I1(n2050), .I2(n2048), .I3(n2049), 
            .O(n22_adj_5232));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i9_4_lut_adj_1753.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1754 (.I0(n1054), .I1(n1055), .I2(GND_net), .I3(GND_net), 
            .O(n38027));
    defparam i1_2_lut_adj_1754.LUT_INIT = 16'h8888;
    SB_LUT4 div_46_LessThan_1606_i37_2_lut (.I0(n2452), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5124));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i7_3_lut (.I0(n2052), .I1(n2043), .I2(n2042), .I3(GND_net), 
            .O(n20_adj_5233));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i7_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_i1062_3_lut (.I0(n1557), .I1(n1624), .I2(n1580), .I3(GND_net), 
            .O(n1656));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1061_3_lut (.I0(n1556), .I1(n1623), .I2(n1580), .I3(GND_net), 
            .O(n1655));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1060_3_lut (.I0(n1555), .I1(n1622), .I2(n1580), .I3(GND_net), 
            .O(n1654));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1054_3_lut (.I0(n1549), .I1(n1616), .I2(n1580), .I3(GND_net), 
            .O(n1648_adj_4815));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i988_3_lut (.I0(n1451), .I1(n1518), .I2(n1481), .I3(GND_net), 
            .O(n1550));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i987_3_lut (.I0(n1450), .I1(n1517), .I2(n1481), .I3(GND_net), 
            .O(n1549));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i986_3_lut (.I0(n1449), .I1(n1516), .I2(n1481), .I3(GND_net), 
            .O(n1548));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i991_3_lut (.I0(n1454), .I1(n1521), .I2(n1481), .I3(GND_net), 
            .O(n1553));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i993_3_lut (.I0(n1456), .I1(n1523), .I2(n1481), .I3(GND_net), 
            .O(n1555));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i989_3_lut (.I0(n1452), .I1(n1519), .I2(n1481), .I3(GND_net), 
            .O(n1551));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i992_3_lut (.I0(n1455), .I1(n1522), .I2(n1481), .I3(GND_net), 
            .O(n1554));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i919_3_lut (.I0(n1350), .I1(n1417), .I2(n1382), .I3(GND_net), 
            .O(n1449));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i919_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i923_3_lut (.I0(n1354), .I1(n1421), .I2(n1382), .I3(GND_net), 
            .O(n1453));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i922_3_lut (.I0(n1353), .I1(n1420_adj_4880), .I2(n1382), 
            .I3(GND_net), .O(n1452));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i920_3_lut (.I0(n1351), .I1(n1418), .I2(n1382), .I3(GND_net), 
            .O(n1450));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i920_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i921_3_lut (.I0(n1352), .I1(n1419), .I2(n1382), .I3(GND_net), 
            .O(n1451));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i921_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i926_3_lut (.I0(n1357), .I1(n1424), .I2(n1382), .I3(GND_net), 
            .O(n1456));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i855_3_lut (.I0(n1254), .I1(n1321), .I2(n1283), .I3(GND_net), 
            .O(n1353));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i854_3_lut (.I0(n1253), .I1(n1320), .I2(n1283), .I3(GND_net), 
            .O(n1352));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i852_3_lut (.I0(n1251), .I1(n1318), .I2(n1283), .I3(GND_net), 
            .O(n1350));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i857_3_lut (.I0(n1256), .I1(n1323), .I2(n1283), .I3(GND_net), 
            .O(n1355));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1606_i43_2_lut (.I0(n2449), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5128));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i41_2_lut (.I0(n2450), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5127));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i856_3_lut (.I0(n1255), .I1(n1322), .I2(n1283), .I3(GND_net), 
            .O(n1354));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i856_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i853_3_lut (.I0(n1252), .I1(n1319), .I2(n1283), .I3(GND_net), 
            .O(n1351));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i786_3_lut (.I0(n1153), .I1(n1220), .I2(n1184), .I3(GND_net), 
            .O(n1252));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i786_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i787_3_lut (.I0(n1154), .I1(n1221), .I2(n1184), .I3(GND_net), 
            .O(n1253));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i787_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i785_3_lut (.I0(n1152), .I1(n1219), .I2(n1184), .I3(GND_net), 
            .O(n1251));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i785_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i789_3_lut (.I0(n1156), .I1(n1223), .I2(n1184), .I3(GND_net), 
            .O(n1255));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i789_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i788_3_lut (.I0(n1155), .I1(n1222), .I2(n1184), .I3(GND_net), 
            .O(n1254));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i788_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i790_3_lut (.I0(n1157), .I1(n1224), .I2(n1184), .I3(GND_net), 
            .O(n1256));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i790_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1755 (.I0(n1256), .I1(n1257), .I2(n1258), .I3(GND_net), 
            .O(n35940));
    defparam i1_3_lut_adj_1755.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1756 (.I0(n1254), .I1(n1250), .I2(n35940), .I3(n1255), 
            .O(n6_adj_4746));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i1_4_lut_adj_1756.LUT_INIT = 16'heccc;
    SB_LUT4 i4_4_lut (.I0(n1251), .I1(n1253), .I2(n1252), .I3(n6_adj_4746), 
            .O(n1283));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i859_3_lut (.I0(n1258), .I1(n1325), .I2(n1283), .I3(GND_net), 
            .O(n1357));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i859_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i858_3_lut (.I0(n1257), .I1(n1324), .I2(n1283), .I3(GND_net), 
            .O(n1356));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i858_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1757 (.I0(n1356), .I1(n1357), .I2(n1358), .I3(GND_net), 
            .O(n35936));
    defparam i1_3_lut_adj_1757.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_4_lut (.I0(n1351), .I1(n1354), .I2(n35936), .I3(n1355), 
            .O(n8_adj_5270));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i2_4_lut.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_2_lut_adj_1758 (.I0(n1350), .I1(n1349), .I2(GND_net), .I3(GND_net), 
            .O(n7_adj_5271));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i1_2_lut_adj_1758.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(n1352), .I1(n7_adj_5271), .I2(n1353), .I3(n8_adj_5270), 
            .O(n1382));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i23_3_lut (.I0(communication_counter[22]), .I1(n11_adj_4798), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1358));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i927_3_lut (.I0(n1358), .I1(n1425), .I2(n1382), .I3(GND_net), 
            .O(n1457));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i925_3_lut (.I0(n1356), .I1(n1423), .I2(n1382), .I3(GND_net), 
            .O(n1455));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i924_3_lut (.I0(n1355), .I1(n1422), .I2(n1382), .I3(GND_net), 
            .O(n1454));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1759 (.I0(n1456), .I1(n1458), .I2(GND_net), .I3(GND_net), 
            .O(n38133));
    defparam i1_2_lut_adj_1759.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_mux_3_i5_3_lut (.I0(encoder0_position[4]), .I1(n21_adj_4666), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n1062));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1760 (.I0(n2046), .I1(n22_adj_5232), .I2(n16_adj_5235), 
            .I3(n2045), .O(n24_adj_5231));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i11_4_lut_adj_1760.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1606_i31_2_lut (.I0(n2455), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5121));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i33_2_lut (.I0(n2454), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5122));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1761 (.I0(n1454), .I1(n38133), .I2(n1455), .I3(n1457), 
            .O(n35969));
    defparam i1_4_lut_adj_1761.LUT_INIT = 16'ha080;
    SB_LUT4 i5_4_lut_adj_1762 (.I0(n35969), .I1(n1451), .I2(n1450), .I3(n1452), 
            .O(n12_adj_5234));
    defparam i5_4_lut_adj_1762.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1763 (.I0(n1453), .I1(n12_adj_5234), .I2(n1449), 
            .I3(n1448), .O(n1481));
    defparam i6_4_lut_adj_1763.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i22_3_lut (.I0(communication_counter[21]), .I1(n12_adj_4797), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1458));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i21_3_lut (.I0(communication_counter[20]), .I1(n13_adj_4796), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1558));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i995_3_lut (.I0(n1458), .I1(n1525), .I2(n1481), .I3(GND_net), 
            .O(n1557));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i994_3_lut (.I0(n1457), .I1(n1524), .I2(n1481), .I3(GND_net), 
            .O(n1556));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1764 (.I0(n1556), .I1(n1557), .I2(n1558), .I3(GND_net), 
            .O(n35966));
    defparam i1_3_lut_adj_1764.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1765 (.I0(n1554), .I1(n1551), .I2(n35966), .I3(n1555), 
            .O(n11_adj_5251));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i3_4_lut_adj_1765.LUT_INIT = 16'heccc;
    SB_LUT4 i5_4_lut_adj_1766 (.I0(n1548), .I1(n1549), .I2(n1547), .I3(n1550), 
            .O(n13_adj_5250));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i5_4_lut_adj_1766.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1767 (.I0(n13_adj_5250), .I1(n11_adj_5251), .I2(n1553), 
            .I3(n1552), .O(n1580));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i7_4_lut_adj_1767.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i990_3_lut (.I0(n1453), .I1(n1520), .I2(n1481), .I3(GND_net), 
            .O(n1552));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1057_3_lut (.I0(n1552), .I1(n1619), .I2(n1580), .I3(GND_net), 
            .O(n1651_adj_4818));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1057_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1058_3_lut (.I0(n1553), .I1(n1620), .I2(n1580), .I3(GND_net), 
            .O(n1652_adj_4819));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1059_3_lut (.I0(n1554), .I1(n1621), .I2(n1580), .I3(GND_net), 
            .O(n1653_adj_4820));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1053_3_lut (.I0(n1548), .I1(n1615), .I2(n1580), .I3(GND_net), 
            .O(n1647_adj_4814));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1053_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1768 (.I0(n1647_adj_4814), .I1(n1646_adj_4813), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5229));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i1_2_lut_adj_1768.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1769 (.I0(n1656), .I1(n1657), .I2(n1658), .I3(GND_net), 
            .O(n35983));
    defparam i1_3_lut_adj_1769.LUT_INIT = 16'hfefe;
    SB_LUT4 i7_4_lut_adj_1770 (.I0(n1653_adj_4820), .I1(n1652_adj_4819), 
            .I2(n1651_adj_4818), .I3(n10_adj_5229), .O(n16_adj_5227));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i7_4_lut_adj_1770.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut_adj_1771 (.I0(n1648_adj_4815), .I1(n1654), .I2(n35983), 
            .I3(n1655), .O(n11_adj_5228));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i2_4_lut_adj_1771.LUT_INIT = 16'heaaa;
    SB_LUT4 i8_4_lut (.I0(n11_adj_5228), .I1(n16_adj_5227), .I2(n1649_adj_4816), 
            .I3(n1650_adj_4817), .O(n1679));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i1055_3_lut (.I0(n1550), .I1(n1617), .I2(n1580), .I3(GND_net), 
            .O(n1649_adj_4816));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1055_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1122_3_lut (.I0(n1649_adj_4816), .I1(n1716), .I2(n1679), 
            .I3(GND_net), .O(n1748));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1122_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13505_3_lut (.I0(setpoint[15]), .I1(n4401), .I2(n37622), 
            .I3(GND_net), .O(n18244));   // verilog/coms.v(127[12] 295[6])
    defparam i13505_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1606_i25_2_lut (.I0(n2458), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5118));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13504_3_lut (.I0(setpoint[14]), .I1(n4400), .I2(n37622), 
            .I3(GND_net), .O(n18243));   // verilog/coms.v(127[12] 295[6])
    defparam i13504_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1606_i27_2_lut (.I0(n2457), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5119));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i29_2_lut (.I0(n2456), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5120));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_i1121_3_lut (.I0(n1648_adj_4815), .I1(n1715), .I2(n1679), 
            .I3(GND_net), .O(n1747));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1121_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1120_3_lut (.I0(n1647_adj_4814), .I1(n1714), .I2(n1679), 
            .I3(GND_net), .O(n1746));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1120_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1772 (.I0(n1746), .I1(n1747), .I2(n1745), .I3(n1748), 
            .O(n16_adj_5358));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i6_4_lut_adj_1772.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1773 (.I0(n1756_adj_4809), .I1(n1757_adj_4810), 
            .I2(n1758_adj_4811), .I3(GND_net), .O(n35975));
    defparam i1_3_lut_adj_1773.LUT_INIT = 16'hfefe;
    SB_LUT4 i8_3_lut (.I0(n1751), .I1(n16_adj_5358), .I2(n1753), .I3(GND_net), 
            .O(n18_adj_5274));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i8_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_adj_1774 (.I0(n1754_adj_4807), .I1(n1749), .I2(n35975), 
            .I3(n1755_adj_4808), .O(n13_adj_4938));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i3_4_lut_adj_1774.LUT_INIT = 16'heccc;
    SB_LUT4 i9_4_lut_adj_1775 (.I0(n13_adj_4938), .I1(n18_adj_5274), .I2(n1752), 
            .I3(n1750), .O(n1778_adj_4812));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i9_4_lut_adj_1775.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1606_i15_2_lut (.I0(n2463), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_5109));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i15_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i17_2_lut (.I0(n2462), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5111));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_4_lut_adj_1776 (.I0(n1052), .I1(n38027), .I2(n1053), .I3(n35946), 
            .O(n1085));
    defparam i1_4_lut_adj_1776.LUT_INIT = 16'hfefa;
    SB_LUT4 rem_4_i655_3_lut (.I0(n958), .I1(n1025), .I2(n986), .I3(GND_net), 
            .O(n1057));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4920));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1606_i19_2_lut (.I0(n2461), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5113));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i21_2_lut (.I0(n2460), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5115));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1606_i23_2_lut (.I0(n2459), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5116));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12_4_lut (.I0(n2051), .I1(n24_adj_5231), .I2(n20_adj_5233), 
            .I3(n2053), .O(n2075_adj_5028));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1606_i35_2_lut (.I0(n2453), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5123));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1608_1_lut (.I0(n2471), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2472));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1608_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4919));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1777 (.I0(one_wire_N_513[9]), .I1(start), .I2(GND_net), 
            .I3(GND_net), .O(n10));
    defparam i1_2_lut_adj_1777.LUT_INIT = 16'heeee;
    SB_LUT4 i7_4_lut_adj_1778 (.I0(one_wire_N_513[8]), .I1(state[1]), .I2(one_wire_N_513[11]), 
            .I3(n10), .O(n16_adj_5359));
    defparam i7_4_lut_adj_1778.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1779 (.I0(one_wire_N_513[6]), .I1(n16_adj_5359), 
            .I2(n11_adj_5254), .I3(one_wire_N_513[10]), .O(n35873));
    defparam i8_4_lut_adj_1779.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i16_3_lut (.I0(communication_counter[15]), .I1(n18_adj_4791), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2058));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34125_4_lut (.I0(n35_adj_5123), .I1(n23_adj_5116), .I2(n21_adj_5115), 
            .I3(n19_adj_5113), .O(n40971));
    defparam i34125_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34862_4_lut (.I0(n17_adj_5111), .I1(n15_adj_5109), .I2(n2464), 
            .I3(n98), .O(n41709));
    defparam i34862_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 rem_4_i1403_3_lut (.I0(n2058), .I1(n2125), .I2(n2075_adj_5028), 
            .I3(GND_net), .O(n2157));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1403_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1402_3_lut (.I0(n2057), .I1(n2124), .I2(n2075_adj_5028), 
            .I3(GND_net), .O(n2156));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1402_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35300_4_lut (.I0(n23_adj_5116), .I1(n21_adj_5115), .I2(n19_adj_5113), 
            .I3(n41709), .O(n42147));
    defparam i35300_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_3_lut_adj_1780 (.I0(n2156), .I1(n2157), .I2(n2158), .I3(GND_net), 
            .O(n35996));
    defparam i1_3_lut_adj_1780.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_mux_3_i24_3_lut (.I0(communication_counter[23]), .I1(n10_adj_4799), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1258));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i719_3_lut (.I0(n1054), .I1(n1121), .I2(n1085), .I3(GND_net), 
            .O(n1153));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i719_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i718_3_lut (.I0(n1053), .I1(n1120), .I2(n1085), .I3(GND_net), 
            .O(n1152));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i718_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i723_3_lut (.I0(n1058), .I1(n1125), .I2(n1085), .I3(GND_net), 
            .O(n1157));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i723_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35288_4_lut (.I0(n29_adj_5120), .I1(n27_adj_5119), .I2(n25_adj_5118), 
            .I3(n42147), .O(n42135));
    defparam i35288_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34129_4_lut (.I0(n35_adj_5123), .I1(n33_adj_5122), .I2(n31_adj_5121), 
            .I3(n42135), .O(n40975));
    defparam i34129_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1606_i12_4_lut (.I0(n1062), .I1(n99), .I2(n2465), 
            .I3(n558), .O(n12_adj_5107));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i12_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i13507_3_lut (.I0(setpoint[17]), .I1(n4403), .I2(n37622), 
            .I3(GND_net), .O(n18246));   // verilog/coms.v(127[12] 295[6])
    defparam i13507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35725_3_lut (.I0(n12_adj_5107), .I1(n87), .I2(n35_adj_5123), 
            .I3(GND_net), .O(n42572));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35725_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_i721_3_lut (.I0(n1056), .I1(n1123), .I2(n1085), .I3(GND_net), 
            .O(n1155));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i721_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i720_3_lut (.I0(n1055), .I1(n1122), .I2(n1085), .I3(GND_net), 
            .O(n1154));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i720_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i651_3_lut (.I0(n954), .I1(n1021), .I2(n986), .I3(GND_net), 
            .O(n1053));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i584_3_lut (.I0(n852), .I1(n6_adj_4668), .I2(n884), 
            .I3(GND_net), .O(n954));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i584_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_mux_3_i30_3_lut (.I0(communication_counter[29]), .I1(n4_adj_4805), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n748));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i31_3_lut (.I0(communication_counter[30]), .I1(n3_adj_4806), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n852));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i28_3_lut (.I0(communication_counter[27]), .I1(n6_adj_4803), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n855));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i29_3_lut (.I0(communication_counter[28]), .I1(n5_adj_4804), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n749));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i27_3_lut (.I0(communication_counter[26]), .I1(n7_adj_4802), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n958));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i586_3_lut (.I0(n749), .I1(n855), .I2(n884), .I3(GND_net), 
            .O(n956));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i586_3_lut.LUT_INIT = 16'h9a9a;
    SB_LUT4 i23146_2_lut (.I0(n855), .I1(n884), .I2(GND_net), .I3(GND_net), 
            .O(n957));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i23146_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 rem_4_i722_3_lut (.I0(n1057), .I1(n1124), .I2(n1085), .I3(GND_net), 
            .O(n1156));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i722_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1781 (.I0(n1156), .I1(n1158), .I2(GND_net), .I3(GND_net), 
            .O(n38031));
    defparam i1_2_lut_adj_1781.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1782 (.I0(n1154), .I1(n38031), .I2(n1155), .I3(n1157), 
            .O(n35942));
    defparam i1_4_lut_adj_1782.LUT_INIT = 16'ha080;
    SB_LUT4 div_46_LessThan_1606_i38_3_lut (.I0(n20_adj_5114), .I1(n83), 
            .I2(n43_adj_5128), .I3(GND_net), .O(n38_adj_5125));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_1519_5 (.CI(n28935), .I0(n2256), .I1(VCC_net), 
            .CO(n28936));
    SB_LUT4 rem_4_add_2055_23_lut (.I0(GND_net), .I1(n3038), .I2(VCC_net), 
            .I3(n28719), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1519_4_lut (.I0(GND_net), .I1(n2257), .I2(VCC_net), 
            .I3(n28934), .O(n2324)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35726_3_lut (.I0(n42572), .I1(n86), .I2(n37_adj_5124), .I3(GND_net), 
            .O(n42573));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35726_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34117_4_lut (.I0(n41_adj_5127), .I1(n39_adj_5126), .I2(n37_adj_5124), 
            .I3(n40971), .O(n40963));
    defparam i34117_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY rem_4_add_1519_4 (.CI(n28934), .I0(n2257), .I1(VCC_net), 
            .CO(n28935));
    SB_CARRY rem_4_add_2055_23 (.CI(n28719), .I0(n3038), .I1(VCC_net), 
            .CO(n28720));
    SB_LUT4 rem_4_add_2055_22_lut (.I0(GND_net), .I1(n3039), .I2(VCC_net), 
            .I3(n28718), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i13506_3_lut (.I0(setpoint[16]), .I1(n4402), .I2(n37622), 
            .I3(GND_net), .O(n18245));   // verilog/coms.v(127[12] 295[6])
    defparam i13506_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35723_4_lut (.I0(n38_adj_5125), .I1(n18_adj_5112), .I2(n43_adj_5128), 
            .I3(n40957), .O(n42570));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35723_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35594_3_lut (.I0(n42573), .I1(n85), .I2(n39_adj_5126), .I3(GND_net), 
            .O(n42441));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35594_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_2055_22 (.CI(n28718), .I0(n3039), .I1(VCC_net), 
            .CO(n28719));
    SB_CARRY add_2354_13 (.CI(n28478), .I0(n2628), .I1(n89), .CO(n28479));
    SB_LUT4 rem_4_add_1519_3_lut (.I0(GND_net), .I1(n2258), .I2(GND_net), 
            .I3(n28933), .O(n2325)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1519_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_21_lut (.I0(GND_net), .I1(n3040), .I2(VCC_net), 
            .I3(n28717), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1519_3 (.CI(n28933), .I0(n2258), .I1(GND_net), 
            .CO(n28934));
    SB_CARRY rem_4_add_2055_21 (.CI(n28717), .I0(n3040), .I1(VCC_net), 
            .CO(n28718));
    SB_CARRY rem_4_add_1519_2 (.CI(VCC_net), .I0(n2358_adj_4940), .I1(VCC_net), 
            .CO(n28933));
    SB_LUT4 rem_4_add_2055_20_lut (.I0(GND_net), .I1(n3041), .I2(VCC_net), 
            .I3(n28716), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_22_lut (.I0(n2372_adj_4939), .I1(n2339), .I2(VCC_net), 
            .I3(n28932), .O(n2438)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_2055_20 (.CI(n28716), .I0(n3041), .I1(VCC_net), 
            .CO(n28717));
    SB_LUT4 rem_4_add_648_5_lut (.I0(GND_net), .I1(n955), .I2(GND_net), 
            .I3(n27917), .O(n1022)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_21_lut (.I0(GND_net), .I1(n2340), .I2(VCC_net), 
            .I3(n28931), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_19_lut (.I0(GND_net), .I1(n3042), .I2(VCC_net), 
            .I3(n28715), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1606_i24_3_lut (.I0(n16_adj_5110), .I1(n91), 
            .I2(n27_adj_5119), .I3(GND_net), .O(n24_adj_5117));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i24_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35943_4_lut (.I0(n24_adj_5117), .I1(n14_adj_5108), .I2(n27_adj_5119), 
            .I3(n41018), .O(n42790));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35943_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35944_3_lut (.I0(n42790), .I1(n90), .I2(n29_adj_5120), .I3(GND_net), 
            .O(n42791));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35944_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35861_3_lut (.I0(n42791), .I1(n89), .I2(n31_adj_5121), .I3(GND_net), 
            .O(n42708));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35861_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35522_4_lut (.I0(n41_adj_5127), .I1(n39_adj_5126), .I2(n37_adj_5124), 
            .I3(n40975), .O(n42369));
    defparam i35522_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35930_4_lut (.I0(n42441), .I1(n42570), .I2(n43_adj_5128), 
            .I3(n40963), .O(n42777));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35930_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35787_3_lut (.I0(n42708), .I1(n88), .I2(n33_adj_5122), .I3(GND_net), 
            .O(n42634));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35787_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i36028_4_lut (.I0(n42634), .I1(n42777), .I2(n43_adj_5128), 
            .I3(n42369), .O(n42875));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36028_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36029_3_lut (.I0(n42875), .I1(n82), .I2(n2448), .I3(GND_net), 
            .O(n42876));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36029_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 add_2354_12_lut (.I0(GND_net), .I1(n2629), .I2(n90), .I3(n28477), 
            .O(n6204)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1783 (.I0(n42876), .I1(n15987), .I2(n81), .I3(n2447), 
            .O(n2471));
    defparam i1_4_lut_adj_1783.LUT_INIT = 16'hceef;
    SB_LUT4 i3_4_lut_adj_1784 (.I0(n35942), .I1(n1152), .I2(n1151), .I3(n1153), 
            .O(n1184));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i3_4_lut_adj_1784.LUT_INIT = 16'hfffe;
    SB_CARRY add_2354_12 (.CI(n28477), .I0(n2629), .I1(n90), .CO(n28478));
    SB_LUT4 add_2354_11_lut (.I0(GND_net), .I1(n2630), .I2(n91), .I3(n28476), 
            .O(n6205)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_19 (.CI(n28715), .I0(n3042), .I1(VCC_net), 
            .CO(n28716));
    SB_CARRY add_2354_11 (.CI(n28476), .I0(n2630), .I1(n91), .CO(n28477));
    SB_CARRY rem_4_add_1586_21 (.CI(n28931), .I0(n2340), .I1(VCC_net), 
            .CO(n28932));
    SB_LUT4 rem_4_add_2055_18_lut (.I0(GND_net), .I1(n3043), .I2(VCC_net), 
            .I3(n28714), .O(n3110)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2354_10_lut (.I0(GND_net), .I1(n2631), .I2(n92), .I3(n28475), 
            .O(n6206)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_20_lut (.I0(GND_net), .I1(n2341), .I2(VCC_net), 
            .I3(n28930), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_18 (.CI(n28714), .I0(n3043), .I1(VCC_net), 
            .CO(n28715));
    SB_CARRY add_2354_10 (.CI(n28475), .I0(n2631), .I1(n92), .CO(n28476));
    SB_LUT4 add_2354_9_lut (.I0(GND_net), .I1(n2632), .I2(n93), .I3(n28474), 
            .O(n6207)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2354_9 (.CI(n28474), .I0(n2632), .I1(n93), .CO(n28475));
    SB_LUT4 add_2354_8_lut (.I0(GND_net), .I1(n2633), .I2(n94), .I3(n28473), 
            .O(n6208)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2354_8 (.CI(n28473), .I0(n2633), .I1(n94), .CO(n28474));
    SB_LUT4 add_2354_7_lut (.I0(GND_net), .I1(n2634), .I2(n95), .I3(n28472), 
            .O(n6209)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_20 (.CI(n28930), .I0(n2341), .I1(VCC_net), 
            .CO(n28931));
    SB_LUT4 rem_4_add_2055_17_lut (.I0(GND_net), .I1(n3044), .I2(VCC_net), 
            .I3(n28713), .O(n3111)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2354_7 (.CI(n28472), .I0(n2634), .I1(n95), .CO(n28473));
    SB_CARRY rem_4_add_2055_17 (.CI(n28713), .I0(n3044), .I1(VCC_net), 
            .CO(n28714));
    SB_LUT4 rem_4_add_1586_19_lut (.I0(GND_net), .I1(n2342), .I2(VCC_net), 
            .I3(n28929), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_19 (.CI(n28929), .I0(n2342), .I1(VCC_net), 
            .CO(n28930));
    SB_LUT4 rem_4_add_2055_16_lut (.I0(GND_net), .I1(n3045), .I2(VCC_net), 
            .I3(n28712), .O(n3112)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2354_6_lut (.I0(GND_net), .I1(n2635), .I2(n96), .I3(n28471), 
            .O(n6210)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2354_6 (.CI(n28471), .I0(n2635), .I1(n96), .CO(n28472));
    SB_LUT4 add_2354_5_lut (.I0(GND_net), .I1(n2636), .I2(n97), .I3(n28470), 
            .O(n6211)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2354_5 (.CI(n28470), .I0(n2636), .I1(n97), .CO(n28471));
    SB_LUT4 add_2354_4_lut (.I0(GND_net), .I1(n2637), .I2(n98), .I3(n28469), 
            .O(n6212)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2354_4 (.CI(n28469), .I0(n2637), .I1(n98), .CO(n28470));
    SB_LUT4 add_2354_3_lut (.I0(GND_net), .I1(n2638), .I2(n99), .I3(n28468), 
            .O(n6213)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2354_3 (.CI(n28468), .I0(n2638), .I1(n99), .CO(n28469));
    SB_LUT4 add_2354_2_lut (.I0(GND_net), .I1(n1064), .I2(n558), .I3(VCC_net), 
            .O(n6214)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2354_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2354_2 (.CI(VCC_net), .I0(n1064), .I1(n558), .CO(n28468));
    SB_LUT4 add_2353_22_lut (.I0(GND_net), .I1(n2534), .I2(n80), .I3(n28467), 
            .O(n6170)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2353_21_lut (.I0(GND_net), .I1(n2535), .I2(n81), .I3(n28466), 
            .O(n6171)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2353_21 (.CI(n28466), .I0(n2535), .I1(n81), .CO(n28467));
    SB_LUT4 add_2353_20_lut (.I0(GND_net), .I1(n2536), .I2(n82), .I3(n28465), 
            .O(n6172)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_18_lut (.I0(GND_net), .I1(n2343), .I2(VCC_net), 
            .I3(n28928), .O(n2410)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_16 (.CI(n28712), .I0(n3045), .I1(VCC_net), 
            .CO(n28713));
    SB_CARRY rem_4_add_1586_18 (.CI(n28928), .I0(n2343), .I1(VCC_net), 
            .CO(n28929));
    SB_LUT4 rem_4_add_1586_17_lut (.I0(GND_net), .I1(n2344), .I2(VCC_net), 
            .I3(n28927), .O(n2411)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_15_lut (.I0(GND_net), .I1(n3046), .I2(VCC_net), 
            .I3(n28711), .O(n3113)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2353_20 (.CI(n28465), .I0(n2536), .I1(n82), .CO(n28466));
    SB_LUT4 add_2353_19_lut (.I0(GND_net), .I1(n2537), .I2(n83), .I3(n28464), 
            .O(n6173)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_15 (.CI(n28711), .I0(n3046), .I1(VCC_net), 
            .CO(n28712));
    SB_CARRY rem_4_add_1586_17 (.CI(n28927), .I0(n2344), .I1(VCC_net), 
            .CO(n28928));
    SB_LUT4 rem_4_add_2055_14_lut (.I0(GND_net), .I1(n3047), .I2(VCC_net), 
            .I3(n28710), .O(n3114)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_14 (.CI(n28710), .I0(n3047), .I1(VCC_net), 
            .CO(n28711));
    SB_LUT4 rem_4_add_1586_16_lut (.I0(GND_net), .I1(n2345), .I2(VCC_net), 
            .I3(n28926), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_16 (.CI(n28926), .I0(n2345), .I1(VCC_net), 
            .CO(n28927));
    SB_LUT4 rem_4_add_2055_13_lut (.I0(GND_net), .I1(n3048), .I2(VCC_net), 
            .I3(n28709), .O(n3115)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_13 (.CI(n28709), .I0(n3048), .I1(VCC_net), 
            .CO(n28710));
    SB_LUT4 rem_4_add_1586_15_lut (.I0(GND_net), .I1(n2346), .I2(VCC_net), 
            .I3(n28925), .O(n2413)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_12_lut (.I0(GND_net), .I1(n3049), .I2(VCC_net), 
            .I3(n28708), .O(n3116)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_15 (.CI(n28925), .I0(n2346), .I1(VCC_net), 
            .CO(n28926));
    SB_CARRY rem_4_add_2055_12 (.CI(n28708), .I0(n3049), .I1(VCC_net), 
            .CO(n28709));
    SB_CARRY add_2353_19 (.CI(n28464), .I0(n2537), .I1(n83), .CO(n28465));
    SB_LUT4 rem_4_add_1586_14_lut (.I0(GND_net), .I1(n2347), .I2(VCC_net), 
            .I3(n28924), .O(n2414)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_11_lut (.I0(GND_net), .I1(n3050), .I2(VCC_net), 
            .I3(n28707), .O(n3117)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2353_18_lut (.I0(GND_net), .I1(n2538), .I2(n84), .I3(n28463), 
            .O(n6174)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_14 (.CI(n28924), .I0(n2347), .I1(VCC_net), 
            .CO(n28925));
    SB_CARRY rem_4_add_2055_11 (.CI(n28707), .I0(n3050), .I1(VCC_net), 
            .CO(n28708));
    SB_CARRY add_2353_18 (.CI(n28463), .I0(n2538), .I1(n84), .CO(n28464));
    SB_LUT4 rem_4_add_2055_10_lut (.I0(GND_net), .I1(n3051), .I2(VCC_net), 
            .I3(n28706), .O(n3118)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2353_17_lut (.I0(GND_net), .I1(n2539), .I2(n85), .I3(n28462), 
            .O(n6175)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2353_17 (.CI(n28462), .I0(n2539), .I1(n85), .CO(n28463));
    SB_LUT4 add_2353_16_lut (.I0(GND_net), .I1(n2540), .I2(n86), .I3(n28461), 
            .O(n6176)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2353_16 (.CI(n28461), .I0(n2540), .I1(n86), .CO(n28462));
    SB_LUT4 add_2353_15_lut (.I0(GND_net), .I1(n2541), .I2(n87), .I3(n28460), 
            .O(n6177)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_13_lut (.I0(GND_net), .I1(n2348), .I2(VCC_net), 
            .I3(n28923), .O(n2415)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_10 (.CI(n28706), .I0(n3051), .I1(VCC_net), 
            .CO(n28707));
    SB_CARRY add_2353_15 (.CI(n28460), .I0(n2541), .I1(n87), .CO(n28461));
    SB_CARRY rem_4_add_1586_13 (.CI(n28923), .I0(n2348), .I1(VCC_net), 
            .CO(n28924));
    SB_LUT4 rem_4_add_2055_9_lut (.I0(GND_net), .I1(n3052), .I2(VCC_net), 
            .I3(n28705), .O(n3119)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_12_lut (.I0(GND_net), .I1(n2349), .I2(VCC_net), 
            .I3(n28922), .O(n2416)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_9 (.CI(n28705), .I0(n3052), .I1(VCC_net), 
            .CO(n28706));
    SB_LUT4 add_2353_14_lut (.I0(GND_net), .I1(n2542), .I2(n88), .I3(n28459), 
            .O(n6178)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2353_14 (.CI(n28459), .I0(n2542), .I1(n88), .CO(n28460));
    SB_LUT4 add_2353_13_lut (.I0(GND_net), .I1(n2543), .I2(n89), .I3(n28458), 
            .O(n6179)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2353_13 (.CI(n28458), .I0(n2543), .I1(n89), .CO(n28459));
    SB_LUT4 add_2353_12_lut (.I0(GND_net), .I1(n2544), .I2(n90), .I3(n28457), 
            .O(n6180)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_12 (.CI(n28922), .I0(n2349), .I1(VCC_net), 
            .CO(n28923));
    SB_LUT4 rem_4_add_2055_8_lut (.I0(GND_net), .I1(n3053), .I2(VCC_net), 
            .I3(n28704), .O(n3120)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2353_12 (.CI(n28457), .I0(n2544), .I1(n90), .CO(n28458));
    SB_CARRY rem_4_add_2055_8 (.CI(n28704), .I0(n3053), .I1(VCC_net), 
            .CO(n28705));
    SB_LUT4 rem_4_add_1586_11_lut (.I0(GND_net), .I1(n2350), .I2(VCC_net), 
            .I3(n28921), .O(n2417)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_11 (.CI(n28921), .I0(n2350), .I1(VCC_net), 
            .CO(n28922));
    SB_LUT4 rem_4_add_2055_7_lut (.I0(GND_net), .I1(n3054), .I2(GND_net), 
            .I3(n28703), .O(n3121)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2353_11_lut (.I0(GND_net), .I1(n2545), .I2(n91), .I3(n28456), 
            .O(n6181)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2353_11 (.CI(n28456), .I0(n2545), .I1(n91), .CO(n28457));
    SB_LUT4 rem_4_add_1586_10_lut (.I0(GND_net), .I1(n2351), .I2(VCC_net), 
            .I3(n28920), .O(n2418)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_7 (.CI(n28703), .I0(n3054), .I1(GND_net), 
            .CO(n28704));
    SB_LUT4 add_2353_10_lut (.I0(GND_net), .I1(n2546), .I2(n92), .I3(n28455), 
            .O(n6182)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_5 (.CI(n27917), .I0(n955), .I1(GND_net), .CO(n27918));
    SB_LUT4 rem_4_add_2055_6_lut (.I0(GND_net), .I1(n3055), .I2(GND_net), 
            .I3(n28702), .O(n3122)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_10 (.CI(n28920), .I0(n2351), .I1(VCC_net), 
            .CO(n28921));
    SB_CARRY rem_4_add_2055_6 (.CI(n28702), .I0(n3055), .I1(GND_net), 
            .CO(n28703));
    SB_LUT4 rem_4_add_1586_9_lut (.I0(GND_net), .I1(n2352), .I2(VCC_net), 
            .I3(n28919), .O(n2419)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_5_lut (.I0(GND_net), .I1(n3056), .I2(VCC_net), 
            .I3(n28701), .O(n3123)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_9 (.CI(n28919), .I0(n2352), .I1(VCC_net), 
            .CO(n28920));
    SB_CARRY rem_4_add_2055_5 (.CI(n28701), .I0(n3056), .I1(VCC_net), 
            .CO(n28702));
    SB_LUT4 rem_4_add_1586_8_lut (.I0(GND_net), .I1(n2353), .I2(VCC_net), 
            .I3(n28918), .O(n2420)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_4_lut (.I0(GND_net), .I1(n3057), .I2(VCC_net), 
            .I3(n28700), .O(n3124)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2353_10 (.CI(n28455), .I0(n2546), .I1(n92), .CO(n28456));
    SB_LUT4 add_2353_9_lut (.I0(GND_net), .I1(n2547), .I2(n93), .I3(n28454), 
            .O(n6183)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2353_9 (.CI(n28454), .I0(n2547), .I1(n93), .CO(n28455));
    SB_LUT4 add_2353_8_lut (.I0(GND_net), .I1(n2548), .I2(n94), .I3(n28453), 
            .O(n6184)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2353_8 (.CI(n28453), .I0(n2548), .I1(n94), .CO(n28454));
    SB_LUT4 rem_4_add_648_4_lut (.I0(GND_net), .I1(n956), .I2(VCC_net), 
            .I3(n27916), .O(n1023)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2353_7_lut (.I0(GND_net), .I1(n2549), .I2(n95), .I3(n28452), 
            .O(n6185)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2353_7 (.CI(n28452), .I0(n2549), .I1(n95), .CO(n28453));
    SB_LUT4 div_46_LessThan_1545_i45_2_lut (.I0(n2358), .I1(n83), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_5106));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i45_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1586_8 (.CI(n28918), .I0(n2353), .I1(VCC_net), 
            .CO(n28919));
    SB_CARRY rem_4_add_2055_4 (.CI(n28700), .I0(n3057), .I1(VCC_net), 
            .CO(n28701));
    SB_LUT4 rem_4_add_1586_7_lut (.I0(GND_net), .I1(n2354), .I2(GND_net), 
            .I3(n28917), .O(n2421)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2055_3_lut (.I0(GND_net), .I1(n3058), .I2(GND_net), 
            .I3(n28699), .O(n3125)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2055_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2353_6_lut (.I0(GND_net), .I1(n2550), .I2(n96), .I3(n28451), 
            .O(n6186)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_7 (.CI(n28917), .I0(n2354), .I1(GND_net), 
            .CO(n28918));
    SB_LUT4 rem_4_add_1586_6_lut (.I0(GND_net), .I1(n2355), .I2(GND_net), 
            .I3(n28916), .O(n2422)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_3 (.CI(n28699), .I0(n3058), .I1(GND_net), 
            .CO(n28700));
    SB_CARRY add_2353_6 (.CI(n28451), .I0(n2550), .I1(n96), .CO(n28452));
    SB_LUT4 div_46_LessThan_1545_i41_2_lut (.I0(n2360), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5104));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i39_2_lut (.I0(n2361), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5102));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2353_5_lut (.I0(GND_net), .I1(n2551), .I2(n97), .I3(n28450), 
            .O(n6187)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2055_2 (.CI(VCC_net), .I0(n3158), .I1(VCC_net), 
            .CO(n28699));
    SB_LUT4 div_46_mux_3_i6_3_lut (.I0(encoder0_position[5]), .I1(n20_adj_4699), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n1061));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1545_i43_2_lut (.I0(n2359), .I1(n84), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5105));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i33_2_lut (.I0(n2364), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5099));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i35_2_lut (.I0(n2363), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5100));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i35_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2353_5 (.CI(n28450), .I0(n2551), .I1(n97), .CO(n28451));
    SB_LUT4 rem_4_add_2122_30_lut (.I0(n3164), .I1(n3131), .I2(VCC_net), 
            .I3(n28698), .O(n3230)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_1586_6 (.CI(n28916), .I0(n2355), .I1(GND_net), 
            .CO(n28917));
    SB_LUT4 i4_4_lut_adj_1785 (.I0(n2154), .I1(n2147), .I2(n35996), .I3(n2155), 
            .O(n18_adj_5336));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i4_4_lut_adj_1785.LUT_INIT = 16'heccc;
    SB_LUT4 div_46_LessThan_1545_i27_2_lut (.I0(n2367), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5096));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2353_4_lut (.I0(GND_net), .I1(n2552), .I2(n98), .I3(n28449), 
            .O(n6188)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_29_lut (.I0(GND_net), .I1(n3132), .I2(VCC_net), 
            .I3(n28697), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1545_i29_2_lut (.I0(n2366), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5097));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i31_2_lut (.I0(n2365), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5098));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_mux_3_i25_3_lut (.I0(communication_counter[24]), .I1(n9_adj_4800), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n1158));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1545_i17_2_lut (.I0(n2372), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5087));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i19_2_lut (.I0(n2371), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5089));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i21_2_lut (.I0(n2370), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5091));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i23_2_lut (.I0(n2369), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5093));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1586_5_lut (.I0(GND_net), .I1(n2356), .I2(VCC_net), 
            .I3(n28915), .O(n2423)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1545_i25_2_lut (.I0(n2368), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5094));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1545_i37_2_lut (.I0(n2362), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5101));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1547_1_lut (.I0(n2381), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2382));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1547_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut_adj_1786 (.I0(n2148), .I1(n2149), .I2(n2150), .I3(n2151), 
            .O(n24_adj_5334));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i10_4_lut_adj_1786.LUT_INIT = 16'hfffe;
    SB_LUT4 i34230_4_lut (.I0(n37_adj_5101), .I1(n25_adj_5094), .I2(n23_adj_5093), 
            .I3(n21_adj_5091), .O(n41076));
    defparam i34230_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34972_4_lut (.I0(n19_adj_5089), .I1(n17_adj_5087), .I2(n2373), 
            .I3(n98), .O(n41819));
    defparam i34972_4_lut.LUT_INIT = 16'hfeef;
    SB_LUT4 i13509_3_lut (.I0(setpoint[19]), .I1(n4405), .I2(n37622), 
            .I3(GND_net), .O(n18248));   // verilog/coms.v(127[12] 295[6])
    defparam i13509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35344_4_lut (.I0(n25_adj_5094), .I1(n23_adj_5093), .I2(n21_adj_5091), 
            .I3(n41819), .O(n42191));
    defparam i35344_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35342_4_lut (.I0(n31_adj_5098), .I1(n29_adj_5097), .I2(n27_adj_5096), 
            .I3(n42191), .O(n42189));
    defparam i35342_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i34232_4_lut (.I0(n37_adj_5101), .I1(n35_adj_5100), .I2(n33_adj_5099), 
            .I3(n42189), .O(n41078));
    defparam i34232_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1545_i14_4_lut (.I0(n1061), .I1(n99), .I2(n2374), 
            .I3(n558), .O(n14_adj_5085));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i14_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i8_4_lut_adj_1787 (.I0(n2142), .I1(n2143), .I2(n2141), .I3(n2144), 
            .O(n22_adj_5335));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i8_4_lut_adj_1787.LUT_INIT = 16'hfffe;
    SB_LUT4 i35490_3_lut (.I0(n14_adj_5085), .I1(n87), .I2(n37_adj_5101), 
            .I3(GND_net), .O(n42337));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35490_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35491_3_lut (.I0(n42337), .I1(n86), .I2(n39_adj_5102), .I3(GND_net), 
            .O(n42338));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35491_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1545_i40_3_lut (.I0(n22_adj_5092), .I1(n83), 
            .I2(n45_adj_5106), .I3(GND_net), .O(n40_adj_5103));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34215_4_lut (.I0(n43_adj_5105), .I1(n41_adj_5104), .I2(n39_adj_5102), 
            .I3(n41076), .O(n41061));
    defparam i34215_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i13508_3_lut (.I0(setpoint[18]), .I1(n4404), .I2(n37622), 
            .I3(GND_net), .O(n18247));   // verilog/coms.v(127[12] 295[6])
    defparam i13508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35587_4_lut (.I0(n40_adj_5103), .I1(n20_adj_5090), .I2(n45_adj_5106), 
            .I3(n41053), .O(n42434));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35587_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34903_3_lut (.I0(n42338), .I1(n85), .I2(n41_adj_5104), .I3(GND_net), 
            .O(n41750));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34903_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_i791_3_lut (.I0(n1158), .I1(n1225), .I2(n1184), .I3(GND_net), 
            .O(n1257));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i791_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1545_i26_3_lut (.I0(n18_adj_5088), .I1(n91), 
            .I2(n29_adj_5097), .I3(GND_net), .O(n26_adj_5095));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35814_4_lut (.I0(n26_adj_5095), .I1(n16_adj_5086), .I2(n29_adj_5097), 
            .I3(n41122), .O(n42661));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35814_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35815_3_lut (.I0(n42661), .I1(n90), .I2(n31_adj_5098), .I3(GND_net), 
            .O(n42662));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35815_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35694_3_lut (.I0(n42662), .I1(n89), .I2(n33_adj_5099), .I3(GND_net), 
            .O(n42541));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35694_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35625_4_lut (.I0(n43_adj_5105), .I1(n41_adj_5104), .I2(n39_adj_5102), 
            .I3(n41078), .O(n42472));
    defparam i35625_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35906_4_lut (.I0(n41750), .I1(n42434), .I2(n45_adj_5106), 
            .I3(n41061), .O(n42753));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35906_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34901_3_lut (.I0(n42541), .I1(n88), .I2(n35_adj_5100), .I3(GND_net), 
            .O(n41748));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34901_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35908_4_lut (.I0(n41748), .I1(n42753), .I2(n45_adj_5106), 
            .I3(n42472), .O(n42755));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35908_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i13511_3_lut (.I0(setpoint[21]), .I1(n4407), .I2(n37622), 
            .I3(GND_net), .O(n18250));   // verilog/coms.v(127[12] 295[6])
    defparam i13511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1788 (.I0(n42755), .I1(n15983), .I2(n82), .I3(n2357), 
            .O(n2381));
    defparam i1_4_lut_adj_1788.LUT_INIT = 16'hceef;
    SB_CARRY add_2353_4 (.CI(n28449), .I0(n2552), .I1(n98), .CO(n28450));
    SB_LUT4 add_2353_3_lut (.I0(GND_net), .I1(n2553), .I2(n99), .I3(n28448), 
            .O(n6189)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_29 (.CI(n28697), .I0(n3132), .I1(VCC_net), 
            .CO(n28698));
    SB_CARRY add_2353_3 (.CI(n28448), .I0(n2553), .I1(n99), .CO(n28449));
    SB_LUT4 add_2353_2_lut (.I0(GND_net), .I1(n1063), .I2(n558), .I3(VCC_net), 
            .O(n6190)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2353_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2353_2 (.CI(VCC_net), .I0(n1063), .I1(n558), .CO(n28448));
    SB_LUT4 div_46_LessThan_1482_i37_2_lut (.I0(n2269), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5081));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i43_2_lut (.I0(n2266), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5084));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i41_2_lut (.I0(n2267), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5083));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i39_2_lut (.I0(n2268), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5082));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i7_3_lut (.I0(encoder0_position[6]), .I1(n19_adj_4700), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n1060));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1482_i19_2_lut (.I0(n2278), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5069));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i19_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i21_2_lut (.I0(n2277), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5071));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i31_2_lut (.I0(n2272), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5078));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i12_4_lut_adj_1789 (.I0(n2145), .I1(n24_adj_5334), .I2(n18_adj_5336), 
            .I3(n2146), .O(n26_adj_5333));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i12_4_lut_adj_1789.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1482_i33_2_lut (.I0(n2271), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5079));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i35_2_lut (.I0(n2270), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5080));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1482_i23_2_lut (.I0(n2276), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5073));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13510_3_lut (.I0(setpoint[20]), .I1(n4406), .I2(n37622), 
            .I3(GND_net), .O(n18249));   // verilog/coms.v(127[12] 295[6])
    defparam i13510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1482_i25_2_lut (.I0(n2275), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5074));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13442_3_lut (.I0(encoder1_position[1]), .I1(n2965), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18181));   // quad.v(35[10] 41[6])
    defparam i13442_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2352_21_lut (.I0(GND_net), .I1(n2447), .I2(n81), .I3(n28447), 
            .O(n6148)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1482_i27_2_lut (.I0(n2274), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5075));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i27_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1586_5 (.CI(n28915), .I0(n2356), .I1(VCC_net), 
            .CO(n28916));
    SB_LUT4 div_46_LessThan_1482_i29_2_lut (.I0(n2273), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5077));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1484_1_lut (.I0(n2288), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2289));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1484_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_add_2122_28_lut (.I0(GND_net), .I1(n3133), .I2(VCC_net), 
            .I3(n28696), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2352_20_lut (.I0(GND_net), .I1(n2448), .I2(n82), .I3(n28446), 
            .O(n6149)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_4_lut (.I0(GND_net), .I1(n2357_adj_4941), .I2(VCC_net), 
            .I3(n28914), .O(n2424)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2352_20 (.CI(n28446), .I0(n2448), .I1(n82), .CO(n28447));
    SB_LUT4 div_46_LessThan_1482_i17_2_lut (.I0(n2279), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_5067));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i17_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i34379_4_lut (.I0(n23_adj_5073), .I1(n21_adj_5071), .I2(n19_adj_5069), 
            .I3(n17_adj_5067), .O(n41226));
    defparam i34379_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY rem_4_add_1586_4 (.CI(n28914), .I0(n2357_adj_4941), .I1(VCC_net), 
            .CO(n28915));
    SB_LUT4 add_2352_19_lut (.I0(GND_net), .I1(n2449), .I2(n83), .I3(n28445), 
            .O(n6150)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34369_4_lut (.I0(n29_adj_5077), .I1(n27_adj_5075), .I2(n25_adj_5074), 
            .I3(n41226), .O(n41216));
    defparam i34369_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY add_2352_19 (.CI(n28445), .I0(n2449), .I1(n83), .CO(n28446));
    SB_LUT4 add_2352_18_lut (.I0(GND_net), .I1(n2450), .I2(n84), .I3(n28444), 
            .O(n6151)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35637_4_lut (.I0(n35_adj_5080), .I1(n33_adj_5079), .I2(n31_adj_5078), 
            .I3(n41216), .O(n42484));
    defparam i35637_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1482_i16_4_lut (.I0(n1060), .I1(n99), .I2(n2280), 
            .I3(n558), .O(n16_adj_5066));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i16_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35494_3_lut (.I0(n16_adj_5066), .I1(n87), .I2(n39_adj_5082), 
            .I3(GND_net), .O(n42341));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35494_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_2122_28 (.CI(n28696), .I0(n3133), .I1(VCC_net), 
            .CO(n28697));
    SB_CARRY add_2352_18 (.CI(n28444), .I0(n2450), .I1(n84), .CO(n28445));
    SB_LUT4 add_2352_17_lut (.I0(GND_net), .I1(n2451), .I2(n85), .I3(n28443), 
            .O(n6152)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2352_17 (.CI(n28443), .I0(n2451), .I1(n85), .CO(n28444));
    SB_LUT4 add_2352_16_lut (.I0(GND_net), .I1(n2452), .I2(n86), .I3(n28442), 
            .O(n6153)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2352_16 (.CI(n28442), .I0(n2452), .I1(n86), .CO(n28443));
    SB_LUT4 add_2352_15_lut (.I0(GND_net), .I1(n2453), .I2(n87), .I3(n28441), 
            .O(n6154)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2352_15 (.CI(n28441), .I0(n2453), .I1(n87), .CO(n28442));
    SB_LUT4 add_2352_14_lut (.I0(GND_net), .I1(n2454), .I2(n88), .I3(n28440), 
            .O(n6155)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2352_14 (.CI(n28440), .I0(n2454), .I1(n88), .CO(n28441));
    SB_LUT4 add_2352_13_lut (.I0(GND_net), .I1(n2455), .I2(n89), .I3(n28439), 
            .O(n6156)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2352_13 (.CI(n28439), .I0(n2455), .I1(n89), .CO(n28440));
    SB_LUT4 add_2352_12_lut (.I0(GND_net), .I1(n2456), .I2(n90), .I3(n28438), 
            .O(n6157)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1586_3_lut (.I0(GND_net), .I1(n2358_adj_4940), .I2(GND_net), 
            .I3(n28913), .O(n2425)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1586_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_27_lut (.I0(GND_net), .I1(n3134), .I2(VCC_net), 
            .I3(n28695), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2352_12 (.CI(n28438), .I0(n2456), .I1(n90), .CO(n28439));
    SB_LUT4 add_2352_11_lut (.I0(GND_net), .I1(n2457), .I2(n91), .I3(n28437), 
            .O(n6158)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2352_11 (.CI(n28437), .I0(n2457), .I1(n91), .CO(n28438));
    SB_LUT4 i35495_3_lut (.I0(n42341), .I1(n86), .I2(n41_adj_5083), .I3(GND_net), 
            .O(n42342));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35495_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_2352_10_lut (.I0(GND_net), .I1(n2458), .I2(n92), .I3(n28436), 
            .O(n6159)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34988_4_lut (.I0(n41_adj_5083), .I1(n39_adj_5082), .I2(n27_adj_5075), 
            .I3(n41222), .O(n41835));
    defparam i34988_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35583_3_lut (.I0(n22_adj_5072), .I1(n93), .I2(n27_adj_5075), 
            .I3(GND_net), .O(n42430));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35583_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34893_3_lut (.I0(n42342), .I1(n85), .I2(n43_adj_5084), .I3(GND_net), 
            .O(n41740));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34893_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i13_4_lut (.I0(n2153), .I1(n26_adj_5333), .I2(n22_adj_5335), 
            .I3(n2152), .O(n2174_adj_4984));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_2352_10 (.CI(n28436), .I0(n2458), .I1(n92), .CO(n28437));
    SB_LUT4 add_2352_9_lut (.I0(GND_net), .I1(n2459), .I2(n93), .I3(n28435), 
            .O(n6160)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1586_3 (.CI(n28913), .I0(n2358_adj_4940), .I1(GND_net), 
            .CO(n28914));
    SB_CARRY add_2352_9 (.CI(n28435), .I0(n2459), .I1(n93), .CO(n28436));
    SB_LUT4 div_46_LessThan_1482_i28_3_lut (.I0(n20_adj_5070), .I1(n91), 
            .I2(n31_adj_5078), .I3(GND_net), .O(n28_adj_5076));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35804_4_lut (.I0(n28_adj_5076), .I1(n18_adj_5068), .I2(n31_adj_5078), 
            .I3(n41212), .O(n42651));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35804_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35805_3_lut (.I0(n42651), .I1(n90), .I2(n33_adj_5079), .I3(GND_net), 
            .O(n42652));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35805_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35700_3_lut (.I0(n42652), .I1(n89), .I2(n35_adj_5080), .I3(GND_net), 
            .O(n42547));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35700_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_2352_8_lut (.I0(GND_net), .I1(n2460), .I2(n94), .I3(n28434), 
            .O(n6161)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2352_8 (.CI(n28434), .I0(n2460), .I1(n94), .CO(n28435));
    SB_CARRY rem_4_add_1586_2 (.CI(VCC_net), .I0(n2458_adj_4875), .I1(VCC_net), 
            .CO(n28913));
    SB_CARRY rem_4_add_2122_27 (.CI(n28695), .I0(n3134), .I1(VCC_net), 
            .CO(n28696));
    SB_LUT4 i34992_4_lut (.I0(n41_adj_5083), .I1(n39_adj_5082), .I2(n37_adj_5081), 
            .I3(n42484), .O(n41839));
    defparam i34992_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 add_2352_7_lut (.I0(GND_net), .I1(n2461), .I2(n95), .I3(n28433), 
            .O(n6162)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35697_4_lut (.I0(n41740), .I1(n42430), .I2(n43_adj_5084), 
            .I3(n41835), .O(n42544));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35697_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 rem_4_add_2122_26_lut (.I0(GND_net), .I1(n3135), .I2(VCC_net), 
            .I3(n28694), .O(n3202)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2352_7 (.CI(n28433), .I0(n2461), .I1(n95), .CO(n28434));
    SB_LUT4 rem_4_add_1653_23_lut (.I0(n2471_adj_4874), .I1(n2438), .I2(VCC_net), 
            .I3(n28912), .O(n2537_adj_4873)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_2122_26 (.CI(n28694), .I0(n3135), .I1(VCC_net), 
            .CO(n28695));
    SB_LUT4 add_2352_6_lut (.I0(GND_net), .I1(n2462), .I2(n96), .I3(n28432), 
            .O(n6163)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_25_lut (.I0(GND_net), .I1(n3136), .I2(VCC_net), 
            .I3(n28693), .O(n3203)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_4 (.CI(n27916), .I0(n956), .I1(VCC_net), .CO(n27917));
    SB_CARRY add_2352_6 (.CI(n28432), .I0(n2462), .I1(n96), .CO(n28433));
    SB_LUT4 add_2352_5_lut (.I0(GND_net), .I1(n2463), .I2(n97), .I3(n28431), 
            .O(n6164)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_22_lut (.I0(GND_net), .I1(n2439), .I2(VCC_net), 
            .I3(n28911), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_25 (.CI(n28693), .I0(n3136), .I1(VCC_net), 
            .CO(n28694));
    SB_CARRY rem_4_add_1653_22 (.CI(n28911), .I0(n2439), .I1(VCC_net), 
            .CO(n28912));
    SB_LUT4 rem_4_add_2122_24_lut (.I0(GND_net), .I1(n3137), .I2(VCC_net), 
            .I3(n28692), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_21_lut (.I0(GND_net), .I1(n2440), .I2(VCC_net), 
            .I3(n28910), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_24 (.CI(n28692), .I0(n3137), .I1(VCC_net), 
            .CO(n28693));
    SB_LUT4 i34891_3_lut (.I0(n42547), .I1(n88), .I2(n37_adj_5081), .I3(GND_net), 
            .O(n41738));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34891_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35959_4_lut (.I0(n41738), .I1(n42544), .I2(n43_adj_5084), 
            .I3(n41839), .O(n42806));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35959_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35960_3_lut (.I0(n42806), .I1(n84), .I2(n2265), .I3(GND_net), 
            .O(n42807));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35960_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1790 (.I0(n42807), .I1(n16000), .I2(n83), .I3(n2264), 
            .O(n2288));
    defparam i1_4_lut_adj_1790.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_1417_i39_2_lut (.I0(n2172), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5062));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i45_2_lut (.I0(n2169), .I1(n85), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_5065));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i43_2_lut (.I0(n2170), .I1(n86), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5064));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i41_2_lut (.I0(n2171), .I1(n87), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5063));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i8_3_lut (.I0(encoder0_position[7]), .I1(n18_adj_4701), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n1059));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1417_i21_2_lut (.I0(n2181), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5049));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i23_2_lut (.I0(n2180), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5051));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_mux_3_i15_3_lut (.I0(communication_counter[14]), .I1(n19_adj_4790), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2158));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34071_3_lut_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(n24782), .I3(start), .O(n40728));
    defparam i34071_3_lut_4_lut.LUT_INIT = 16'hff10;
    SB_LUT4 div_46_LessThan_1417_i33_2_lut (.I0(n2175), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5059));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i33_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1653_21 (.CI(n28910), .I0(n2440), .I1(VCC_net), 
            .CO(n28911));
    SB_LUT4 rem_4_add_2122_23_lut (.I0(GND_net), .I1(n3138), .I2(VCC_net), 
            .I3(n28691), .O(n3205)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_23 (.CI(n28691), .I0(n3138), .I1(VCC_net), 
            .CO(n28692));
    SB_LUT4 rem_4_add_1653_20_lut (.I0(GND_net), .I1(n2441), .I2(VCC_net), 
            .I3(n28909), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_20 (.CI(n28909), .I0(n2441), .I1(VCC_net), 
            .CO(n28910));
    SB_LUT4 rem_4_add_2122_22_lut (.I0(GND_net), .I1(n3139), .I2(VCC_net), 
            .I3(n28690), .O(n3206)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2352_5 (.CI(n28431), .I0(n2463), .I1(n97), .CO(n28432));
    SB_LUT4 rem_4_add_1653_19_lut (.I0(GND_net), .I1(n2442), .I2(VCC_net), 
            .I3(n28908), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2352_4_lut (.I0(GND_net), .I1(n2464), .I2(n98), .I3(n28430), 
            .O(n6165)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2352_4 (.CI(n28430), .I0(n2464), .I1(n98), .CO(n28431));
    SB_LUT4 add_2352_3_lut (.I0(GND_net), .I1(n2465), .I2(n99), .I3(n28429), 
            .O(n6166)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2352_3 (.CI(n28429), .I0(n2465), .I1(n99), .CO(n28430));
    SB_LUT4 add_2352_2_lut (.I0(GND_net), .I1(n1062), .I2(n558), .I3(VCC_net), 
            .O(n6167)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2352_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2352_2 (.CI(VCC_net), .I0(n1062), .I1(n558), .CO(n28429));
    SB_LUT4 add_2351_20_lut (.I0(GND_net), .I1(n2357), .I2(n82), .I3(n28428), 
            .O(n6127)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2351_19_lut (.I0(GND_net), .I1(n2358), .I2(n83), .I3(n28427), 
            .O(n6128)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2351_19 (.CI(n28427), .I0(n2358), .I1(n83), .CO(n28428));
    SB_LUT4 add_2351_18_lut (.I0(GND_net), .I1(n2359), .I2(n84), .I3(n28426), 
            .O(n6129)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2351_18 (.CI(n28426), .I0(n2359), .I1(n84), .CO(n28427));
    SB_LUT4 add_2351_17_lut (.I0(GND_net), .I1(n2360), .I2(n85), .I3(n28425), 
            .O(n6130)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2351_17 (.CI(n28425), .I0(n2360), .I1(n85), .CO(n28426));
    SB_LUT4 add_2351_16_lut (.I0(GND_net), .I1(n2361), .I2(n86), .I3(n28424), 
            .O(n6131)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2351_16 (.CI(n28424), .I0(n2361), .I1(n86), .CO(n28425));
    SB_LUT4 add_2351_15_lut (.I0(GND_net), .I1(n2362), .I2(n87), .I3(n28423), 
            .O(n6132)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2351_15 (.CI(n28423), .I0(n2362), .I1(n87), .CO(n28424));
    SB_LUT4 add_2351_14_lut (.I0(GND_net), .I1(n2363), .I2(n88), .I3(n28422), 
            .O(n6133)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2351_14 (.CI(n28422), .I0(n2363), .I1(n88), .CO(n28423));
    SB_LUT4 add_2351_13_lut (.I0(GND_net), .I1(n2364), .I2(n89), .I3(n28421), 
            .O(n6134)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2351_13 (.CI(n28421), .I0(n2364), .I1(n89), .CO(n28422));
    SB_LUT4 add_2351_12_lut (.I0(GND_net), .I1(n2365), .I2(n90), .I3(n28420), 
            .O(n6135)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2351_12 (.CI(n28420), .I0(n2365), .I1(n90), .CO(n28421));
    SB_LUT4 add_2351_11_lut (.I0(GND_net), .I1(n2366), .I2(n91), .I3(n28419), 
            .O(n6136)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2351_11 (.CI(n28419), .I0(n2366), .I1(n91), .CO(n28420));
    SB_LUT4 add_2351_10_lut (.I0(GND_net), .I1(n2367), .I2(n92), .I3(n28418), 
            .O(n6137)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2351_10 (.CI(n28418), .I0(n2367), .I1(n92), .CO(n28419));
    SB_LUT4 add_2351_9_lut (.I0(GND_net), .I1(n2368), .I2(n93), .I3(n28417), 
            .O(n6138)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2351_9 (.CI(n28417), .I0(n2368), .I1(n93), .CO(n28418));
    SB_LUT4 add_2351_8_lut (.I0(GND_net), .I1(n2369), .I2(n94), .I3(n28416), 
            .O(n6139)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_3_lut_4_lut (.I0(\neo_pixel_transmitter.done ), .I1(state[0]), 
            .I2(n24782), .I3(state[1]), .O(n37483));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 div_46_LessThan_1417_i35_2_lut (.I0(n2174), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5060));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i37_2_lut (.I0(n2173), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5061));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i37_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2351_8 (.CI(n28416), .I0(n2369), .I1(n94), .CO(n28417));
    SB_LUT4 add_2351_7_lut (.I0(GND_net), .I1(n2370), .I2(n95), .I3(n28415), 
            .O(n6140)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2351_7 (.CI(n28415), .I0(n2370), .I1(n95), .CO(n28416));
    SB_LUT4 div_46_LessThan_1417_i29_2_lut (.I0(n2177), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5056));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i31_2_lut (.I0(n2176), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5058));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 add_2351_6_lut (.I0(GND_net), .I1(n2371), .I2(n96), .I3(n28414), 
            .O(n6141)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_22 (.CI(n28690), .I0(n3139), .I1(VCC_net), 
            .CO(n28691));
    SB_CARRY add_2351_6 (.CI(n28414), .I0(n2371), .I1(n96), .CO(n28415));
    SB_LUT4 div_46_LessThan_1417_i25_2_lut (.I0(n2179), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5053));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1417_i27_2_lut (.I0(n2178), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5055));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1419_1_lut (.I0(n2192), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2193));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1419_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1417_i19_2_lut (.I0(n2182), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_5047));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i19_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1653_19 (.CI(n28908), .I0(n2442), .I1(VCC_net), 
            .CO(n28909));
    SB_LUT4 rem_4_add_2122_21_lut (.I0(GND_net), .I1(n3140), .I2(VCC_net), 
            .I3(n28689), .O(n3207)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2351_5_lut (.I0(GND_net), .I1(n2372), .I2(n97), .I3(n28413), 
            .O(n6142)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34427_4_lut (.I0(n25_adj_5053), .I1(n23_adj_5051), .I2(n21_adj_5049), 
            .I3(n19_adj_5047), .O(n41274));
    defparam i34427_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34421_4_lut (.I0(n31_adj_5058), .I1(n29_adj_5056), .I2(n27_adj_5055), 
            .I3(n41274), .O(n41268));
    defparam i34421_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35643_4_lut (.I0(n37_adj_5061), .I1(n35_adj_5060), .I2(n33_adj_5059), 
            .I3(n41268), .O(n42490));
    defparam i35643_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1417_i18_4_lut (.I0(n1059), .I1(n99), .I2(n2183), 
            .I3(n558), .O(n18_adj_5046));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i18_4_lut.LUT_INIT = 16'h0317;
    SB_CARRY add_2351_5 (.CI(n28413), .I0(n2372), .I1(n97), .CO(n28414));
    SB_LUT4 add_2351_4_lut (.I0(GND_net), .I1(n2373), .I2(n98), .I3(n28412), 
            .O(n6143)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35500_3_lut (.I0(n18_adj_5046), .I1(n87), .I2(n41_adj_5063), 
            .I3(GND_net), .O(n42347));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35500_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35501_3_lut (.I0(n42347), .I1(n86), .I2(n43_adj_5064), .I3(GND_net), 
            .O(n42348));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35501_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35030_4_lut (.I0(n43_adj_5064), .I1(n41_adj_5063), .I2(n29_adj_5056), 
            .I3(n41272), .O(n41877));
    defparam i35030_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_46_LessThan_1417_i26_3_lut (.I0(n24_adj_5052), .I1(n93), 
            .I2(n29_adj_5056), .I3(GND_net), .O(n26_adj_5054));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i26_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34887_3_lut (.I0(n42348), .I1(n85), .I2(n45_adj_5065), .I3(GND_net), 
            .O(n41734));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34887_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1417_i30_3_lut (.I0(n22_adj_5050), .I1(n91), 
            .I2(n33_adj_5059), .I3(GND_net), .O(n30_adj_5057));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35796_4_lut (.I0(n30_adj_5057), .I1(n20_adj_5048), .I2(n33_adj_5059), 
            .I3(n41258), .O(n42643));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35796_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35797_3_lut (.I0(n42643), .I1(n90), .I2(n35_adj_5060), .I3(GND_net), 
            .O(n42644));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35797_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_2351_4 (.CI(n28412), .I0(n2373), .I1(n98), .CO(n28413));
    SB_LUT4 add_2351_3_lut (.I0(GND_net), .I1(n2374), .I2(n99), .I3(n28411), 
            .O(n6144)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_18_lut (.I0(GND_net), .I1(n2443), .I2(VCC_net), 
            .I3(n28907), .O(n2510)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35702_3_lut (.I0(n42644), .I1(n89), .I2(n37_adj_5061), .I3(GND_net), 
            .O(n42549));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35702_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_2122_21 (.CI(n28689), .I0(n3140), .I1(VCC_net), 
            .CO(n28690));
    SB_LUT4 i35036_4_lut (.I0(n43_adj_5064), .I1(n41_adj_5063), .I2(n39_adj_5062), 
            .I3(n42490), .O(n41883));
    defparam i35036_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35578_4_lut (.I0(n41734), .I1(n26_adj_5054), .I2(n45_adj_5065), 
            .I3(n41877), .O(n42425));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35578_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34885_3_lut (.I0(n42549), .I1(n88), .I2(n39_adj_5062), .I3(GND_net), 
            .O(n41732));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34885_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35580_4_lut (.I0(n41732), .I1(n42425), .I2(n45_adj_5065), 
            .I3(n41883), .O(n42427));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35580_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1791 (.I0(n42427), .I1(n15901), .I2(n84), .I3(n2168), 
            .O(n2192));
    defparam i1_4_lut_adj_1791.LUT_INIT = 16'hceef;
    SB_LUT4 i13159_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n13302), 
            .I3(GND_net), .O(n17898));   // verilog/coms.v(127[12] 295[6])
    defparam i13159_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2351_3 (.CI(n28411), .I0(n2374), .I1(n99), .CO(n28412));
    SB_LUT4 add_2351_2_lut (.I0(GND_net), .I1(n1061), .I2(n558), .I3(VCC_net), 
            .O(n6145)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2351_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_648_3_lut (.I0(GND_net), .I1(n957), .I2(VCC_net), 
            .I3(n27915), .O(n1024)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1350_i41_2_lut (.I0(n2072), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5045));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1350_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i37_2_lut (.I0(n2074), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5043));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1350_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i39_2_lut (.I0(n2073), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5044));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1350_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i35_2_lut (.I0(n2075), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5042));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1350_i35_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2351_2 (.CI(VCC_net), .I0(n1061), .I1(n558), .CO(n28411));
    SB_LUT4 add_2350_19_lut (.I0(GND_net), .I1(n2264), .I2(n83), .I3(n28410), 
            .O(n6107)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2350_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_20_lut (.I0(GND_net), .I1(n3141), .I2(VCC_net), 
            .I3(n28688), .O(n3208)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_mux_3_i9_3_lut (.I0(encoder0_position[8]), .I1(n17_adj_4702), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n1058_adj_4737));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_2350_18_lut (.I0(GND_net), .I1(n2265), .I2(n84), .I3(n28409), 
            .O(n6108)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2350_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2350_18 (.CI(n28409), .I0(n2265), .I1(n84), .CO(n28410));
    SB_LUT4 add_2350_17_lut (.I0(GND_net), .I1(n2266), .I2(n85), .I3(n28408), 
            .O(n6109)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2350_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2350_17 (.CI(n28408), .I0(n2266), .I1(n85), .CO(n28409));
    SB_LUT4 add_2350_16_lut (.I0(GND_net), .I1(n2267), .I2(n86), .I3(n28407), 
            .O(n6110)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2350_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2350_16 (.CI(n28407), .I0(n2267), .I1(n86), .CO(n28408));
    SB_LUT4 add_2350_15_lut (.I0(GND_net), .I1(n2268), .I2(n87), .I3(n28406), 
            .O(n6111)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2350_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2350_15 (.CI(n28406), .I0(n2268), .I1(n87), .CO(n28407));
    SB_LUT4 add_2350_14_lut (.I0(GND_net), .I1(n2269), .I2(n88), .I3(n28405), 
            .O(n6112)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2350_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2350_14 (.CI(n28405), .I0(n2269), .I1(n88), .CO(n28406));
    SB_LUT4 add_2350_13_lut (.I0(GND_net), .I1(n2270), .I2(n89), .I3(n28404), 
            .O(n6113)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2350_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2350_13 (.CI(n28404), .I0(n2270), .I1(n89), .CO(n28405));
    SB_LUT4 add_2350_12_lut (.I0(GND_net), .I1(n2271), .I2(n90), .I3(n28403), 
            .O(n6114)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2350_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2350_12 (.CI(n28403), .I0(n2271), .I1(n90), .CO(n28404));
    SB_LUT4 add_2350_11_lut (.I0(GND_net), .I1(n2272), .I2(n91), .I3(n28402), 
            .O(n6115)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2350_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2350_11 (.CI(n28402), .I0(n2272), .I1(n91), .CO(n28403));
    SB_LUT4 add_2350_10_lut (.I0(GND_net), .I1(n2273), .I2(n92), .I3(n28401), 
            .O(n6116)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2350_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2350_10 (.CI(n28401), .I0(n2273), .I1(n92), .CO(n28402));
    SB_LUT4 add_2350_9_lut (.I0(GND_net), .I1(n2274), .I2(n93), .I3(n28400), 
            .O(n6117)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2350_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2350_9 (.CI(n28400), .I0(n2274), .I1(n93), .CO(n28401));
    SB_LUT4 add_2350_8_lut (.I0(GND_net), .I1(n2275), .I2(n94), .I3(n28399), 
            .O(n6118)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2350_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2350_8 (.CI(n28399), .I0(n2275), .I1(n94), .CO(n28400));
    SB_LUT4 add_2350_7_lut (.I0(GND_net), .I1(n2276), .I2(n95), .I3(n28398), 
            .O(n6119)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2350_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_18 (.CI(n28907), .I0(n2443), .I1(VCC_net), 
            .CO(n28908));
    SB_LUT4 rem_4_add_1653_17_lut (.I0(GND_net), .I1(n2444), .I2(VCC_net), 
            .I3(n28906), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_20 (.CI(n28688), .I0(n3141), .I1(VCC_net), 
            .CO(n28689));
    SB_CARRY add_2350_7 (.CI(n28398), .I0(n2276), .I1(n95), .CO(n28399));
    SB_LUT4 add_2350_6_lut (.I0(GND_net), .I1(n2277), .I2(n96), .I3(n28397), 
            .O(n6120)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2350_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2350_6 (.CI(n28397), .I0(n2277), .I1(n96), .CO(n28398));
    SB_LUT4 add_2350_5_lut (.I0(GND_net), .I1(n2278), .I2(n97), .I3(n28396), 
            .O(n6121)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2350_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2350_5 (.CI(n28396), .I0(n2278), .I1(n97), .CO(n28397));
    SB_LUT4 add_2350_4_lut (.I0(GND_net), .I1(n2279), .I2(n98), .I3(n28395), 
            .O(n6122)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2350_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2350_4 (.CI(n28395), .I0(n2279), .I1(n98), .CO(n28396));
    SB_LUT4 add_2350_3_lut (.I0(GND_net), .I1(n2280), .I2(n99), .I3(n28394), 
            .O(n6123)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2350_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2350_3 (.CI(n28394), .I0(n2280), .I1(n99), .CO(n28395));
    SB_LUT4 add_2350_2_lut (.I0(GND_net), .I1(n1060), .I2(n558), .I3(VCC_net), 
            .O(n6124)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2350_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2350_2 (.CI(VCC_net), .I0(n1060), .I1(n558), .CO(n28394));
    SB_LUT4 add_2349_18_lut (.I0(GND_net), .I1(n2168), .I2(n84), .I3(n28393), 
            .O(n6088)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2349_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2349_17_lut (.I0(GND_net), .I1(n2169), .I2(n85), .I3(n28392), 
            .O(n6089)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2349_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2349_17 (.CI(n28392), .I0(n2169), .I1(n85), .CO(n28393));
    SB_LUT4 add_2349_16_lut (.I0(GND_net), .I1(n2170), .I2(n86), .I3(n28391), 
            .O(n6090)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2349_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2349_16 (.CI(n28391), .I0(n2170), .I1(n86), .CO(n28392));
    SB_LUT4 add_2349_15_lut (.I0(GND_net), .I1(n2171), .I2(n87), .I3(n28390), 
            .O(n6091)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2349_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2349_15 (.CI(n28390), .I0(n2171), .I1(n87), .CO(n28391));
    SB_LUT4 add_2349_14_lut (.I0(GND_net), .I1(n2172), .I2(n88), .I3(n28389), 
            .O(n6092)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2349_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_3 (.CI(n27915), .I0(n957), .I1(VCC_net), .CO(n27916));
    SB_LUT4 rem_4_mux_3_i14_3_lut (.I0(communication_counter[13]), .I1(n20_adj_4789), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2258));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1350_i23_2_lut (.I0(n2081), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5032));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1350_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i25_2_lut (.I0(n2080), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5034));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1350_i25_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2349_14 (.CI(n28389), .I0(n2172), .I1(n88), .CO(n28390));
    SB_LUT4 add_2349_13_lut (.I0(GND_net), .I1(n2173), .I2(n89), .I3(n28388), 
            .O(n6093)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2349_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1350_i27_2_lut (.I0(n2079), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5036));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1350_i27_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1653_17 (.CI(n28906), .I0(n2444), .I1(VCC_net), 
            .CO(n28907));
    SB_LUT4 div_46_LessThan_1350_i29_2_lut (.I0(n2078), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5038));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1350_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i31_2_lut (.I0(n2077), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5039));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1350_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1350_i33_2_lut (.I0(n2076), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5041));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1350_i33_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_2349_13 (.CI(n28388), .I0(n2173), .I1(n89), .CO(n28389));
    SB_LUT4 add_2349_12_lut (.I0(GND_net), .I1(n2174), .I2(n90), .I3(n28387), 
            .O(n6094)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2349_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_19_lut (.I0(GND_net), .I1(n3142), .I2(VCC_net), 
            .I3(n28687), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i1352_1_lut (.I0(n2093), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n2094));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1352_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1471_3_lut (.I0(n2158), .I1(n2225), .I2(n2174_adj_4984), 
            .I3(GND_net), .O(n2257));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1350_i21_2_lut (.I0(n2082), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_5030));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1350_i21_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i34482_4_lut (.I0(n27_adj_5036), .I1(n25_adj_5034), .I2(n23_adj_5032), 
            .I3(n21_adj_5030), .O(n41329));
    defparam i34482_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34474_4_lut (.I0(n33_adj_5041), .I1(n31_adj_5039), .I2(n29_adj_5038), 
            .I3(n41329), .O(n41321));
    defparam i34474_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 rem_4_i1470_3_lut (.I0(n2157), .I1(n2224), .I2(n2174_adj_4984), 
            .I3(GND_net), .O(n2256));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1470_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_2349_12 (.CI(n28387), .I0(n2174), .I1(n90), .CO(n28388));
    SB_LUT4 add_2349_11_lut (.I0(GND_net), .I1(n2175), .I2(n91), .I3(n28386), 
            .O(n6095)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2349_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1350_i20_4_lut (.I0(n1058_adj_4737), .I1(n99), 
            .I2(n2083), .I3(n558), .O(n20_adj_5029));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1350_i20_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_1350_i28_3_lut (.I0(n26_adj_5035), .I1(n93), 
            .I2(n31_adj_5039), .I3(GND_net), .O(n28_adj_5037));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1350_i28_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY add_2349_11 (.CI(n28386), .I0(n2175), .I1(n91), .CO(n28387));
    SB_DFF communication_counter_1222__i1 (.Q(communication_counter[1]), .C(LED_c), 
           .D(n164));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_LUT4 add_2349_10_lut (.I0(GND_net), .I1(n2176), .I2(n92), .I3(n28385), 
            .O(n6096)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2349_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2349_10 (.CI(n28385), .I0(n2176), .I1(n92), .CO(n28386));
    SB_LUT4 div_46_LessThan_1350_i32_3_lut (.I0(n24_adj_5033), .I1(n91), 
            .I2(n35_adj_5042), .I3(GND_net), .O(n32_adj_5040));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1350_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35878_4_lut (.I0(n32_adj_5040), .I1(n22_adj_5031), .I2(n35_adj_5042), 
            .I3(n41314), .O(n42725));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35878_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35879_3_lut (.I0(n42725), .I1(n90), .I2(n37_adj_5043), .I3(GND_net), 
            .O(n42726));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35879_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35710_3_lut (.I0(n42726), .I1(n89), .I2(n39_adj_5044), .I3(GND_net), 
            .O(n42557));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35710_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 add_2349_9_lut (.I0(GND_net), .I1(n2177), .I2(n93), .I3(n28384), 
            .O(n6097)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2349_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2349_9 (.CI(n28384), .I0(n2177), .I1(n93), .CO(n28385));
    SB_LUT4 add_2349_8_lut (.I0(GND_net), .I1(n2178), .I2(n94), .I3(n28383), 
            .O(n6098)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2349_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2349_8 (.CI(n28383), .I0(n2178), .I1(n94), .CO(n28384));
    SB_LUT4 add_2349_7_lut (.I0(GND_net), .I1(n2179), .I2(n95), .I3(n28382), 
            .O(n6099)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2349_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2349_7 (.CI(n28382), .I0(n2179), .I1(n95), .CO(n28383));
    SB_LUT4 add_2349_6_lut (.I0(GND_net), .I1(n2180), .I2(n96), .I3(n28381), 
            .O(n6100)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2349_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2349_6 (.CI(n28381), .I0(n2180), .I1(n96), .CO(n28382));
    SB_LUT4 add_2349_5_lut (.I0(GND_net), .I1(n2181), .I2(n97), .I3(n28380), 
            .O(n6101)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2349_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2349_5 (.CI(n28380), .I0(n2181), .I1(n97), .CO(n28381));
    SB_LUT4 add_2349_4_lut (.I0(GND_net), .I1(n2182), .I2(n98), .I3(n28379), 
            .O(n6102)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2349_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2349_4 (.CI(n28379), .I0(n2182), .I1(n98), .CO(n28380));
    SB_LUT4 add_2349_3_lut (.I0(GND_net), .I1(n2183), .I2(n99), .I3(n28378), 
            .O(n6103)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2349_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2349_3 (.CI(n28378), .I0(n2183), .I1(n99), .CO(n28379));
    SB_LUT4 add_2349_2_lut (.I0(GND_net), .I1(n1059), .I2(n558), .I3(VCC_net), 
            .O(n6104)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2349_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2349_2 (.CI(VCC_net), .I0(n1059), .I1(n558), .CO(n28378));
    SB_LUT4 add_2348_17_lut (.I0(GND_net), .I1(n2069), .I2(n85), .I3(n28377), 
            .O(n6070)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2348_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2348_16_lut (.I0(GND_net), .I1(n2070), .I2(n86), .I3(n28376), 
            .O(n6071)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2348_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2348_16 (.CI(n28376), .I0(n2070), .I1(n86), .CO(n28377));
    SB_LUT4 add_2348_15_lut (.I0(GND_net), .I1(n2071), .I2(n87), .I3(n28375), 
            .O(n6072)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2348_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2348_15 (.CI(n28375), .I0(n2071), .I1(n87), .CO(n28376));
    SB_LUT4 add_2348_14_lut (.I0(GND_net), .I1(n2072), .I2(n88), .I3(n28374), 
            .O(n6073)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2348_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2348_14 (.CI(n28374), .I0(n2072), .I1(n88), .CO(n28375));
    SB_LUT4 add_2348_13_lut (.I0(GND_net), .I1(n2073), .I2(n89), .I3(n28373), 
            .O(n6074)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2348_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2348_13 (.CI(n28373), .I0(n2073), .I1(n89), .CO(n28374));
    SB_LUT4 add_2348_12_lut (.I0(GND_net), .I1(n2074), .I2(n90), .I3(n28372), 
            .O(n6075)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2348_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2348_12 (.CI(n28372), .I0(n2074), .I1(n90), .CO(n28373));
    SB_LUT4 add_2348_11_lut (.I0(GND_net), .I1(n2075), .I2(n91), .I3(n28371), 
            .O(n6076)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2348_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2348_11 (.CI(n28371), .I0(n2075), .I1(n91), .CO(n28372));
    SB_LUT4 add_2348_10_lut (.I0(GND_net), .I1(n2076), .I2(n92), .I3(n28370), 
            .O(n6077)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2348_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2348_10 (.CI(n28370), .I0(n2076), .I1(n92), .CO(n28371));
    SB_LUT4 add_2348_9_lut (.I0(GND_net), .I1(n2077), .I2(n93), .I3(n28369), 
            .O(n6078)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2348_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2348_9 (.CI(n28369), .I0(n2077), .I1(n93), .CO(n28370));
    SB_LUT4 add_2348_8_lut (.I0(GND_net), .I1(n2078), .I2(n94), .I3(n28368), 
            .O(n6079)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2348_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2348_8 (.CI(n28368), .I0(n2078), .I1(n94), .CO(n28369));
    SB_LUT4 add_2348_7_lut (.I0(GND_net), .I1(n2079), .I2(n95), .I3(n28367), 
            .O(n6080)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2348_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2348_7 (.CI(n28367), .I0(n2079), .I1(n95), .CO(n28368));
    SB_LUT4 add_2348_6_lut (.I0(GND_net), .I1(n2080), .I2(n96), .I3(n28366), 
            .O(n6081)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2348_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2348_6 (.CI(n28366), .I0(n2080), .I1(n96), .CO(n28367));
    SB_LUT4 add_2348_5_lut (.I0(GND_net), .I1(n2081), .I2(n97), .I3(n28365), 
            .O(n6082)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2348_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2348_5 (.CI(n28365), .I0(n2081), .I1(n97), .CO(n28366));
    SB_LUT4 add_2348_4_lut (.I0(GND_net), .I1(n2082), .I2(n98), .I3(n28364), 
            .O(n6083)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2348_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2348_4 (.CI(n28364), .I0(n2082), .I1(n98), .CO(n28365));
    SB_LUT4 add_2348_3_lut (.I0(GND_net), .I1(n2083), .I2(n99), .I3(n28363), 
            .O(n6084)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2348_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2348_3 (.CI(n28363), .I0(n2083), .I1(n99), .CO(n28364));
    SB_LUT4 add_2348_2_lut (.I0(GND_net), .I1(n1058_adj_4737), .I2(n558), 
            .I3(VCC_net), .O(n6085)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2348_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2348_2 (.CI(VCC_net), .I0(n1058_adj_4737), .I1(n558), 
            .CO(n28363));
    SB_LUT4 add_2347_16_lut (.I0(GND_net), .I1(n1967), .I2(n86), .I3(n28362), 
            .O(n6053)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2347_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2347_15_lut (.I0(GND_net), .I1(n1968), .I2(n87), .I3(n28361), 
            .O(n6054)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2347_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2347_15 (.CI(n28361), .I0(n1968), .I1(n87), .CO(n28362));
    SB_LUT4 add_2347_14_lut (.I0(GND_net), .I1(n1969), .I2(n88), .I3(n28360), 
            .O(n6055)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2347_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2347_14 (.CI(n28360), .I0(n1969), .I1(n88), .CO(n28361));
    SB_LUT4 add_2347_13_lut (.I0(GND_net), .I1(n1970), .I2(n89), .I3(n28359), 
            .O(n6056)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2347_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2347_13 (.CI(n28359), .I0(n1970), .I1(n89), .CO(n28360));
    SB_LUT4 add_2347_12_lut (.I0(GND_net), .I1(n1971), .I2(n90), .I3(n28358), 
            .O(n6057)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2347_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2347_12 (.CI(n28358), .I0(n1971), .I1(n90), .CO(n28359));
    SB_LUT4 add_2347_11_lut (.I0(GND_net), .I1(n1972), .I2(n91), .I3(n28357), 
            .O(n6058)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2347_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2347_11 (.CI(n28357), .I0(n1972), .I1(n91), .CO(n28358));
    SB_LUT4 add_2347_10_lut (.I0(GND_net), .I1(n1973), .I2(n92), .I3(n28356), 
            .O(n6059)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2347_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2347_10 (.CI(n28356), .I0(n1973), .I1(n92), .CO(n28357));
    SB_LUT4 add_2347_9_lut (.I0(GND_net), .I1(n1974), .I2(n93), .I3(n28355), 
            .O(n6060)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2347_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2347_9 (.CI(n28355), .I0(n1974), .I1(n93), .CO(n28356));
    SB_LUT4 add_2347_8_lut (.I0(GND_net), .I1(n1975), .I2(n94), .I3(n28354), 
            .O(n6061)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2347_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2347_8 (.CI(n28354), .I0(n1975), .I1(n94), .CO(n28355));
    SB_LUT4 add_2347_7_lut (.I0(GND_net), .I1(n1976), .I2(n95), .I3(n28353), 
            .O(n6062)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2347_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2347_7 (.CI(n28353), .I0(n1976), .I1(n95), .CO(n28354));
    SB_LUT4 add_2347_6_lut (.I0(GND_net), .I1(n1977), .I2(n96), .I3(n28352), 
            .O(n6063)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2347_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2347_6 (.CI(n28352), .I0(n1977), .I1(n96), .CO(n28353));
    SB_LUT4 add_2347_5_lut (.I0(GND_net), .I1(n1978), .I2(n97), .I3(n28351), 
            .O(n6064)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2347_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2347_5 (.CI(n28351), .I0(n1978), .I1(n97), .CO(n28352));
    SB_LUT4 add_2347_4_lut (.I0(GND_net), .I1(n1979), .I2(n98), .I3(n28350), 
            .O(n6065)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2347_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2347_4 (.CI(n28350), .I0(n1979), .I1(n98), .CO(n28351));
    SB_LUT4 add_2347_3_lut (.I0(GND_net), .I1(n1980), .I2(n99), .I3(n28349), 
            .O(n6066)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2347_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2347_3 (.CI(n28349), .I0(n1980), .I1(n99), .CO(n28350));
    SB_LUT4 add_2347_2_lut (.I0(GND_net), .I1(n1057_adj_4736), .I2(n558), 
            .I3(VCC_net), .O(n6067)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2347_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2347_2 (.CI(VCC_net), .I0(n1057_adj_4736), .I1(n558), 
            .CO(n28349));
    SB_LUT4 add_2346_15_lut (.I0(GND_net), .I1(n1862), .I2(n87), .I3(n28348), 
            .O(n6037)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2346_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2346_14_lut (.I0(GND_net), .I1(n1863), .I2(n88), .I3(n28347), 
            .O(n6038)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2346_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2346_14 (.CI(n28347), .I0(n1863), .I1(n88), .CO(n28348));
    SB_LUT4 add_2346_13_lut (.I0(GND_net), .I1(n1864), .I2(n89), .I3(n28346), 
            .O(n6039)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2346_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2346_13 (.CI(n28346), .I0(n1864), .I1(n89), .CO(n28347));
    SB_LUT4 add_2346_12_lut (.I0(GND_net), .I1(n1865), .I2(n90), .I3(n28345), 
            .O(n6040)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2346_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2346_12 (.CI(n28345), .I0(n1865), .I1(n90), .CO(n28346));
    SB_LUT4 add_2346_11_lut (.I0(GND_net), .I1(n1866), .I2(n91), .I3(n28344), 
            .O(n6041)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2346_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2346_11 (.CI(n28344), .I0(n1866), .I1(n91), .CO(n28345));
    SB_LUT4 add_2346_10_lut (.I0(GND_net), .I1(n1867), .I2(n92), .I3(n28343), 
            .O(n6042)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2346_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2346_10 (.CI(n28343), .I0(n1867), .I1(n92), .CO(n28344));
    SB_LUT4 add_2346_9_lut (.I0(GND_net), .I1(n1868), .I2(n93), .I3(n28342), 
            .O(n6043)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2346_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2346_9 (.CI(n28342), .I0(n1868), .I1(n93), .CO(n28343));
    SB_LUT4 add_2346_8_lut (.I0(GND_net), .I1(n1869), .I2(n94), .I3(n28341), 
            .O(n6044)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2346_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2346_8 (.CI(n28341), .I0(n1869), .I1(n94), .CO(n28342));
    SB_LUT4 add_2346_7_lut (.I0(GND_net), .I1(n1870), .I2(n95), .I3(n28340), 
            .O(n6045)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2346_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2346_7 (.CI(n28340), .I0(n1870), .I1(n95), .CO(n28341));
    SB_LUT4 add_2346_6_lut (.I0(GND_net), .I1(n1871), .I2(n96), .I3(n28339), 
            .O(n6046)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2346_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2346_6 (.CI(n28339), .I0(n1871), .I1(n96), .CO(n28340));
    SB_LUT4 i35653_4_lut (.I0(n39_adj_5044), .I1(n37_adj_5043), .I2(n35_adj_5042), 
            .I3(n41321), .O(n42500));
    defparam i35653_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_2122_19 (.CI(n28687), .I0(n3142), .I1(VCC_net), 
            .CO(n28688));
    SB_LUT4 rem_4_add_648_2_lut (.I0(GND_net), .I1(n958), .I2(GND_net), 
            .I3(VCC_net), .O(n1025)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_648_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_18_lut (.I0(GND_net), .I1(n3143), .I2(VCC_net), 
            .I3(n28686), .O(n3210)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2346_5_lut (.I0(GND_net), .I1(n1872), .I2(n97), .I3(n28338), 
            .O(n6047)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2346_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_648_2 (.CI(VCC_net), .I0(n958), .I1(GND_net), .CO(n27915));
    SB_LUT4 rem_4_add_1653_16_lut (.I0(GND_net), .I1(n2445), .I2(VCC_net), 
            .I3(n28905), .O(n2512)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2346_5 (.CI(n28338), .I0(n1872), .I1(n97), .CO(n28339));
    SB_CARRY rem_4_add_1653_16 (.CI(n28905), .I0(n2445), .I1(VCC_net), 
            .CO(n28906));
    SB_CARRY rem_4_add_2122_18 (.CI(n28686), .I0(n3143), .I1(VCC_net), 
            .CO(n28687));
    SB_LUT4 rem_4_add_2122_17_lut (.I0(GND_net), .I1(n3144), .I2(VCC_net), 
            .I3(n28685), .O(n3211)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_17 (.CI(n28685), .I0(n3144), .I1(VCC_net), 
            .CO(n28686));
    SB_LUT4 add_2346_4_lut (.I0(GND_net), .I1(n1873), .I2(n98), .I3(n28337), 
            .O(n6048)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2346_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_16_lut (.I0(GND_net), .I1(n3145), .I2(VCC_net), 
            .I3(n28684), .O(n3212)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2346_4 (.CI(n28337), .I0(n1873), .I1(n98), .CO(n28338));
    SB_LUT4 rem_4_add_1653_15_lut (.I0(GND_net), .I1(n2446), .I2(VCC_net), 
            .I3(n28904), .O(n2513)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_16 (.CI(n28684), .I0(n3145), .I1(VCC_net), 
            .CO(n28685));
    SB_CARRY rem_4_add_1653_15 (.CI(n28904), .I0(n2446), .I1(VCC_net), 
            .CO(n28905));
    SB_LUT4 rem_4_add_1653_14_lut (.I0(GND_net), .I1(n2447_adj_4887), .I2(VCC_net), 
            .I3(n28903), .O(n2514)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2346_3_lut (.I0(GND_net), .I1(n1874), .I2(n99), .I3(n28336), 
            .O(n6049)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2346_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2346_3 (.CI(n28336), .I0(n1874), .I1(n99), .CO(n28337));
    SB_LUT4 i35880_4_lut (.I0(n28_adj_5037), .I1(n20_adj_5029), .I2(n31_adj_5039), 
            .I3(n41324), .O(n42727));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35880_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34875_3_lut (.I0(n42557), .I1(n88), .I2(n41_adj_5045), .I3(GND_net), 
            .O(n41722));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34875_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_1653_14 (.CI(n28903), .I0(n2447_adj_4887), .I1(VCC_net), 
            .CO(n28904));
    SB_LUT4 rem_4_add_1653_13_lut (.I0(GND_net), .I1(n2448_adj_4886), .I2(VCC_net), 
            .I3(n28902), .O(n2515)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_13 (.CI(n28902), .I0(n2448_adj_4886), .I1(VCC_net), 
            .CO(n28903));
    SB_LUT4 rem_4_add_2122_15_lut (.I0(GND_net), .I1(n3146), .I2(VCC_net), 
            .I3(n28683), .O(n3213)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_12_lut (.I0(GND_net), .I1(n2449_adj_4885), .I2(VCC_net), 
            .I3(n28901), .O(n2516)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_15 (.CI(n28683), .I0(n3146), .I1(VCC_net), 
            .CO(n28684));
    SB_CARRY rem_4_add_1653_12 (.CI(n28901), .I0(n2449_adj_4885), .I1(VCC_net), 
            .CO(n28902));
    SB_LUT4 rem_4_add_2122_14_lut (.I0(GND_net), .I1(n3147), .I2(VCC_net), 
            .I3(n28682), .O(n3214)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_14 (.CI(n28682), .I0(n3147), .I1(VCC_net), 
            .CO(n28683));
    SB_LUT4 rem_4_add_1653_11_lut (.I0(GND_net), .I1(n2450_adj_4884), .I2(VCC_net), 
            .I3(n28900), .O(n2517)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_13_lut (.I0(GND_net), .I1(n3148), .I2(VCC_net), 
            .I3(n28681), .O(n3215)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_13 (.CI(n28681), .I0(n3148), .I1(VCC_net), 
            .CO(n28682));
    SB_LUT4 add_2346_2_lut (.I0(GND_net), .I1(n1056_adj_4735), .I2(n558), 
            .I3(VCC_net), .O(n6050)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2346_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_12_lut (.I0(GND_net), .I1(n3149), .I2(VCC_net), 
            .I3(n28680), .O(n3216)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_11 (.CI(n28900), .I0(n2450_adj_4884), .I1(VCC_net), 
            .CO(n28901));
    SB_LUT4 rem_4_add_1653_10_lut (.I0(GND_net), .I1(n2451_adj_4883), .I2(VCC_net), 
            .I3(n28899), .O(n2518)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35934_4_lut (.I0(n41722), .I1(n42727), .I2(n41_adj_5045), 
            .I3(n42500), .O(n42781));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35934_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_2346_2 (.CI(VCC_net), .I0(n1056_adj_4735), .I1(n558), 
            .CO(n28336));
    SB_CARRY rem_4_add_1653_10 (.CI(n28899), .I0(n2451_adj_4883), .I1(VCC_net), 
            .CO(n28900));
    SB_CARRY rem_4_add_2122_12 (.CI(n28680), .I0(n3149), .I1(VCC_net), 
            .CO(n28681));
    SB_LUT4 add_2345_14_lut (.I0(GND_net), .I1(n1754), .I2(n88), .I3(n28335), 
            .O(n6022)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2345_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2345_13_lut (.I0(GND_net), .I1(n1755), .I2(n89), .I3(n28334), 
            .O(n6023)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2345_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_11_lut (.I0(GND_net), .I1(n3150), .I2(VCC_net), 
            .I3(n28679), .O(n3217)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35935_3_lut (.I0(n42781), .I1(n87), .I2(n2071), .I3(GND_net), 
            .O(n42782));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35935_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35883_3_lut (.I0(n42782), .I1(n86), .I2(n2070), .I3(GND_net), 
            .O(n42730));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35883_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 rem_4_add_1653_9_lut (.I0(GND_net), .I1(n2452_adj_4882), .I2(VCC_net), 
            .I3(n28898), .O(n2519)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2345_13 (.CI(n28334), .I0(n1755), .I1(n89), .CO(n28335));
    SB_LUT4 add_2345_12_lut (.I0(GND_net), .I1(n1756), .I2(n90), .I3(n28333), 
            .O(n6024)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2345_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2345_12 (.CI(n28333), .I0(n1756), .I1(n90), .CO(n28334));
    SB_CARRY rem_4_add_2122_11 (.CI(n28679), .I0(n3150), .I1(VCC_net), 
            .CO(n28680));
    SB_CARRY rem_4_add_1653_9 (.CI(n28898), .I0(n2452_adj_4882), .I1(VCC_net), 
            .CO(n28899));
    SB_LUT4 add_2345_11_lut (.I0(GND_net), .I1(n1757), .I2(n91), .I3(n28332), 
            .O(n6025)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2345_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1792 (.I0(n42730), .I1(n15897), .I2(n85), .I3(n2069), 
            .O(n2093));
    defparam i1_4_lut_adj_1792.LUT_INIT = 16'hceef;
    SB_CARRY add_2345_11 (.CI(n28332), .I0(n1757), .I1(n91), .CO(n28333));
    SB_LUT4 add_2345_10_lut (.I0(GND_net), .I1(n1758), .I2(n92), .I3(n28331), 
            .O(n6026)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2345_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2345_10 (.CI(n28331), .I0(n1758), .I1(n92), .CO(n28332));
    SB_LUT4 add_2345_9_lut (.I0(GND_net), .I1(n1759), .I2(n93), .I3(n28330), 
            .O(n6027)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2345_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2345_9 (.CI(n28330), .I0(n1759), .I1(n93), .CO(n28331));
    SB_LUT4 add_2345_8_lut (.I0(GND_net), .I1(n1760), .I2(n94), .I3(n28329), 
            .O(n6028)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2345_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2345_8 (.CI(n28329), .I0(n1760), .I1(n94), .CO(n28330));
    SB_LUT4 add_2345_7_lut (.I0(GND_net), .I1(n1761), .I2(n95), .I3(n28328), 
            .O(n6029)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2345_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2345_7 (.CI(n28328), .I0(n1761), .I1(n95), .CO(n28329));
    SB_LUT4 add_2345_6_lut (.I0(GND_net), .I1(n1762), .I2(n96), .I3(n28327), 
            .O(n6030)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2345_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2345_6 (.CI(n28327), .I0(n1762), .I1(n96), .CO(n28328));
    SB_LUT4 add_2345_5_lut (.I0(GND_net), .I1(n1763), .I2(n97), .I3(n28326), 
            .O(n6031)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2345_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2345_5 (.CI(n28326), .I0(n1763), .I1(n97), .CO(n28327));
    SB_LUT4 add_2345_4_lut (.I0(GND_net), .I1(n1764), .I2(n98), .I3(n28325), 
            .O(n6032)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2345_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2345_4 (.CI(n28325), .I0(n1764), .I1(n98), .CO(n28326));
    SB_LUT4 add_2345_3_lut (.I0(GND_net), .I1(n1765), .I2(n99), .I3(n28324), 
            .O(n6033)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2345_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2345_3 (.CI(n28324), .I0(n1765), .I1(n99), .CO(n28325));
    SB_LUT4 add_2345_2_lut (.I0(GND_net), .I1(n1055_adj_4734), .I2(n558), 
            .I3(VCC_net), .O(n6034)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2345_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2345_2 (.CI(VCC_net), .I0(n1055_adj_4734), .I1(n558), 
            .CO(n28324));
    SB_LUT4 add_2344_13_lut (.I0(GND_net), .I1(n1643), .I2(n89), .I3(n28323), 
            .O(n6008)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2344_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2344_12_lut (.I0(GND_net), .I1(n1644), .I2(n90), .I3(n28322), 
            .O(n6009)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2344_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2344_12 (.CI(n28322), .I0(n1644), .I1(n90), .CO(n28323));
    SB_LUT4 add_2344_11_lut (.I0(GND_net), .I1(n1645), .I2(n91), .I3(n28321), 
            .O(n6010)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2344_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2344_11 (.CI(n28321), .I0(n1645), .I1(n91), .CO(n28322));
    SB_LUT4 add_2344_10_lut (.I0(GND_net), .I1(n1646), .I2(n92), .I3(n28320), 
            .O(n6011)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2344_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2344_10 (.CI(n28320), .I0(n1646), .I1(n92), .CO(n28321));
    SB_LUT4 add_2344_9_lut (.I0(GND_net), .I1(n1647), .I2(n93), .I3(n28319), 
            .O(n6012)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2344_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2344_9 (.CI(n28319), .I0(n1647), .I1(n93), .CO(n28320));
    SB_LUT4 add_2344_8_lut (.I0(GND_net), .I1(n1648), .I2(n94), .I3(n28318), 
            .O(n6013)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2344_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2344_8 (.CI(n28318), .I0(n1648), .I1(n94), .CO(n28319));
    SB_LUT4 add_2344_7_lut (.I0(GND_net), .I1(n1649), .I2(n95), .I3(n28317), 
            .O(n6014)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2344_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2344_7 (.CI(n28317), .I0(n1649), .I1(n95), .CO(n28318));
    SB_LUT4 add_2344_6_lut (.I0(GND_net), .I1(n1650), .I2(n96), .I3(n28316), 
            .O(n6015)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2344_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2344_6 (.CI(n28316), .I0(n1650), .I1(n96), .CO(n28317));
    SB_LUT4 add_2344_5_lut (.I0(GND_net), .I1(n1651), .I2(n97), .I3(n28315), 
            .O(n6016)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2344_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2344_5 (.CI(n28315), .I0(n1651), .I1(n97), .CO(n28316));
    SB_LUT4 add_2344_4_lut (.I0(GND_net), .I1(n1652), .I2(n98), .I3(n28314), 
            .O(n6017)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2344_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2344_4 (.CI(n28314), .I0(n1652), .I1(n98), .CO(n28315));
    SB_LUT4 add_2344_3_lut (.I0(GND_net), .I1(n1653), .I2(n99), .I3(n28313), 
            .O(n6018)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2344_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2344_3 (.CI(n28313), .I0(n1653), .I1(n99), .CO(n28314));
    SB_LUT4 add_2344_2_lut (.I0(GND_net), .I1(n1054_adj_4733), .I2(n558), 
            .I3(VCC_net), .O(n6019)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2344_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2344_2 (.CI(VCC_net), .I0(n1054_adj_4733), .I1(n558), 
            .CO(n28313));
    SB_LUT4 add_2343_12_lut (.I0(GND_net), .I1(n1529), .I2(n90), .I3(n28312), 
            .O(n5995)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2343_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2343_11_lut (.I0(GND_net), .I1(n1530), .I2(n91), .I3(n28311), 
            .O(n5996)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2343_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2343_11 (.CI(n28311), .I0(n1530), .I1(n91), .CO(n28312));
    SB_LUT4 add_2343_10_lut (.I0(GND_net), .I1(n1531), .I2(n92), .I3(n28310), 
            .O(n5997)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2343_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2343_10 (.CI(n28310), .I0(n1531), .I1(n92), .CO(n28311));
    SB_LUT4 add_2343_9_lut (.I0(GND_net), .I1(n1532), .I2(n93), .I3(n28309), 
            .O(n5998)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2343_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2343_9 (.CI(n28309), .I0(n1532), .I1(n93), .CO(n28310));
    SB_LUT4 add_2343_8_lut (.I0(GND_net), .I1(n1533), .I2(n94), .I3(n28308), 
            .O(n5999)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2343_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2343_8 (.CI(n28308), .I0(n1533), .I1(n94), .CO(n28309));
    SB_LUT4 add_2343_7_lut (.I0(GND_net), .I1(n1534), .I2(n95), .I3(n28307), 
            .O(n6000)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2343_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2343_7 (.CI(n28307), .I0(n1534), .I1(n95), .CO(n28308));
    SB_LUT4 add_2343_6_lut (.I0(GND_net), .I1(n1535), .I2(n96), .I3(n28306), 
            .O(n6001)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2343_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2343_6 (.CI(n28306), .I0(n1535), .I1(n96), .CO(n28307));
    SB_LUT4 add_2343_5_lut (.I0(GND_net), .I1(n1536), .I2(n97), .I3(n28305), 
            .O(n6002)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2343_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_8_lut (.I0(GND_net), .I1(n2453_adj_4881), .I2(VCC_net), 
            .I3(n28897), .O(n2520)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2343_5 (.CI(n28305), .I0(n1536), .I1(n97), .CO(n28306));
    SB_CARRY rem_4_add_1653_8 (.CI(n28897), .I0(n2453_adj_4881), .I1(VCC_net), 
            .CO(n28898));
    SB_LUT4 add_2343_4_lut (.I0(GND_net), .I1(n1537), .I2(n98), .I3(n28304), 
            .O(n6003)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2343_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2343_4 (.CI(n28304), .I0(n1537), .I1(n98), .CO(n28305));
    SB_LUT4 add_2343_3_lut (.I0(GND_net), .I1(n1538), .I2(n99), .I3(n28303), 
            .O(n6004)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2343_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2343_3 (.CI(n28303), .I0(n1538), .I1(n99), .CO(n28304));
    SB_LUT4 add_2343_2_lut (.I0(GND_net), .I1(n1053_adj_4732), .I2(n558), 
            .I3(VCC_net), .O(n6005)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2343_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2343_2 (.CI(VCC_net), .I0(n1053_adj_4732), .I1(n558), 
            .CO(n28303));
    SB_LUT4 add_2342_11_lut (.I0(GND_net), .I1(n1412), .I2(n91), .I3(n28302), 
            .O(n5983)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2342_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2342_10_lut (.I0(GND_net), .I1(n1413), .I2(n92), .I3(n28301), 
            .O(n5984)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2342_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2342_10 (.CI(n28301), .I0(n1413), .I1(n92), .CO(n28302));
    SB_LUT4 add_2342_9_lut (.I0(GND_net), .I1(n1414), .I2(n93), .I3(n28300), 
            .O(n5985)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2342_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2342_9 (.CI(n28300), .I0(n1414), .I1(n93), .CO(n28301));
    SB_LUT4 add_2342_8_lut (.I0(GND_net), .I1(n1415), .I2(n94), .I3(n28299), 
            .O(n5986)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2342_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2342_8 (.CI(n28299), .I0(n1415), .I1(n94), .CO(n28300));
    SB_LUT4 add_2342_7_lut (.I0(GND_net), .I1(n1416), .I2(n95), .I3(n28298), 
            .O(n5987)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2342_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2342_7 (.CI(n28298), .I0(n1416), .I1(n95), .CO(n28299));
    SB_LUT4 add_2342_6_lut (.I0(GND_net), .I1(n1417_adj_4739), .I2(n96), 
            .I3(n28297), .O(n5988)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2342_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2342_6 (.CI(n28297), .I0(n1417_adj_4739), .I1(n96), .CO(n28298));
    SB_LUT4 add_2342_5_lut (.I0(GND_net), .I1(n1418_adj_4740), .I2(n97), 
            .I3(n28296), .O(n5989)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2342_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2342_5 (.CI(n28296), .I0(n1418_adj_4740), .I1(n97), .CO(n28297));
    SB_LUT4 add_2342_4_lut (.I0(GND_net), .I1(n1419_adj_4741), .I2(n98), 
            .I3(n28295), .O(n5990)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2342_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2342_4 (.CI(n28295), .I0(n1419_adj_4741), .I1(n98), .CO(n28296));
    SB_LUT4 add_2342_3_lut (.I0(GND_net), .I1(n1420), .I2(n99), .I3(n28294), 
            .O(n5991)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2342_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2342_3 (.CI(n28294), .I0(n1420), .I1(n99), .CO(n28295));
    SB_LUT4 add_2342_2_lut (.I0(GND_net), .I1(n1052_adj_4731), .I2(n558), 
            .I3(VCC_net), .O(n5992)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2342_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2342_2 (.CI(VCC_net), .I0(n1052_adj_4731), .I1(n558), 
            .CO(n28294));
    SB_LUT4 add_2341_10_lut (.I0(GND_net), .I1(n1292), .I2(n92), .I3(n28293), 
            .O(n5972)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2341_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2341_9_lut (.I0(GND_net), .I1(n1293), .I2(n93), .I3(n28292), 
            .O(n5973)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2341_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2341_9 (.CI(n28292), .I0(n1293), .I1(n93), .CO(n28293));
    SB_LUT4 add_2341_8_lut (.I0(GND_net), .I1(n1294), .I2(n94), .I3(n28291), 
            .O(n5974)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2341_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2341_8 (.CI(n28291), .I0(n1294), .I1(n94), .CO(n28292));
    SB_LUT4 add_2341_7_lut (.I0(GND_net), .I1(n1295), .I2(n95), .I3(n28290), 
            .O(n5975)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2341_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2341_7 (.CI(n28290), .I0(n1295), .I1(n95), .CO(n28291));
    SB_LUT4 add_2341_6_lut (.I0(GND_net), .I1(n1296), .I2(n96), .I3(n28289), 
            .O(n5976)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2341_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2341_6 (.CI(n28289), .I0(n1296), .I1(n96), .CO(n28290));
    SB_LUT4 add_2341_5_lut (.I0(GND_net), .I1(n1297), .I2(n97), .I3(n28288), 
            .O(n5977)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2341_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2341_5 (.CI(n28288), .I0(n1297), .I1(n97), .CO(n28289));
    SB_LUT4 add_2341_4_lut (.I0(GND_net), .I1(n1298), .I2(n98), .I3(n28287), 
            .O(n5978)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2341_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2341_4 (.CI(n28287), .I0(n1298), .I1(n98), .CO(n28288));
    SB_LUT4 add_2341_3_lut (.I0(GND_net), .I1(n1299), .I2(n99), .I3(n28286), 
            .O(n5979)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2341_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2341_3 (.CI(n28286), .I0(n1299), .I1(n99), .CO(n28287));
    SB_LUT4 add_2341_2_lut (.I0(GND_net), .I1(n1051), .I2(n558), .I3(VCC_net), 
            .O(n5980)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2341_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2341_2 (.CI(VCC_net), .I0(n1051), .I1(n558), .CO(n28286));
    SB_LUT4 add_2340_9_lut (.I0(GND_net), .I1(n1169), .I2(n93), .I3(n28285), 
            .O(n5962)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2340_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2340_8_lut (.I0(GND_net), .I1(n1170_adj_4738), .I2(n94), 
            .I3(n28284), .O(n5963)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2340_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2340_8 (.CI(n28284), .I0(n1170_adj_4738), .I1(n94), .CO(n28285));
    SB_LUT4 add_2340_7_lut (.I0(GND_net), .I1(n1171), .I2(n95), .I3(n28283), 
            .O(n5964)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2340_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2340_7 (.CI(n28283), .I0(n1171), .I1(n95), .CO(n28284));
    SB_LUT4 add_2340_6_lut (.I0(GND_net), .I1(n1172), .I2(n96), .I3(n28282), 
            .O(n5965)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2340_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2340_6 (.CI(n28282), .I0(n1172), .I1(n96), .CO(n28283));
    SB_LUT4 add_2340_5_lut (.I0(GND_net), .I1(n1173), .I2(n97), .I3(n28281), 
            .O(n5966)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2340_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2340_5 (.CI(n28281), .I0(n1173), .I1(n97), .CO(n28282));
    SB_LUT4 add_2340_4_lut (.I0(GND_net), .I1(n1174), .I2(n98), .I3(n28280), 
            .O(n5967)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2340_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2340_4 (.CI(n28280), .I0(n1174), .I1(n98), .CO(n28281));
    SB_LUT4 add_2340_3_lut (.I0(GND_net), .I1(n1175), .I2(n99), .I3(n28279), 
            .O(n5968)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2340_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2340_3 (.CI(n28279), .I0(n1175), .I1(n99), .CO(n28280));
    SB_LUT4 add_2340_2_lut (.I0(GND_net), .I1(n1050), .I2(n558), .I3(VCC_net), 
            .O(n5969)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2340_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2340_2 (.CI(VCC_net), .I0(n1050), .I1(n558), .CO(n28279));
    SB_LUT4 add_2339_8_lut (.I0(GND_net), .I1(n1043), .I2(n94), .I3(n28278), 
            .O(n5953)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2339_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2339_7_lut (.I0(GND_net), .I1(n1044), .I2(n95), .I3(n28277), 
            .O(n5954)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2339_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2339_7 (.CI(n28277), .I0(n1044), .I1(n95), .CO(n28278));
    SB_LUT4 add_2339_6_lut (.I0(GND_net), .I1(n1045), .I2(n96), .I3(n28276), 
            .O(n5955)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2339_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2339_6 (.CI(n28276), .I0(n1045), .I1(n96), .CO(n28277));
    SB_LUT4 add_2339_5_lut (.I0(GND_net), .I1(n1046), .I2(n97), .I3(n28275), 
            .O(n5956)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2339_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2339_5 (.CI(n28275), .I0(n1046), .I1(n97), .CO(n28276));
    SB_LUT4 add_2339_4_lut (.I0(GND_net), .I1(n1047), .I2(n98), .I3(n28274), 
            .O(n5957)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2339_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2339_4 (.CI(n28274), .I0(n1047), .I1(n98), .CO(n28275));
    SB_LUT4 add_2339_3_lut (.I0(GND_net), .I1(n1048), .I2(n99), .I3(n28273), 
            .O(n5958)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2339_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2339_3 (.CI(n28273), .I0(n1048), .I1(n99), .CO(n28274));
    SB_LUT4 add_2339_2_lut (.I0(GND_net), .I1(n1049), .I2(n558), .I3(VCC_net), 
            .O(n5959)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2339_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2339_2 (.CI(VCC_net), .I0(n1049), .I1(n558), .CO(n28273));
    SB_LUT4 add_2338_7_lut (.I0(GND_net), .I1(n914), .I2(n95), .I3(n28272), 
            .O(n5945)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2338_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2338_6_lut (.I0(GND_net), .I1(n915), .I2(n96), .I3(n28271), 
            .O(n5946)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2338_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2338_6 (.CI(n28271), .I0(n915), .I1(n96), .CO(n28272));
    SB_LUT4 add_2338_5_lut (.I0(GND_net), .I1(n916), .I2(n97), .I3(n28270), 
            .O(n5947)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2338_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2338_5 (.CI(n28270), .I0(n916), .I1(n97), .CO(n28271));
    SB_LUT4 add_2338_4_lut (.I0(GND_net), .I1(n917), .I2(n98), .I3(n28269), 
            .O(n5948)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2338_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2338_4 (.CI(n28269), .I0(n917), .I1(n98), .CO(n28270));
    SB_LUT4 add_2338_3_lut (.I0(GND_net), .I1(n918), .I2(n99), .I3(n28268), 
            .O(n5949)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2338_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2338_3 (.CI(n28268), .I0(n918), .I1(n99), .CO(n28269));
    SB_LUT4 i13160_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n13302), 
            .I3(GND_net), .O(n17899));   // verilog/coms.v(127[12] 295[6])
    defparam i13160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_add_2122_10_lut (.I0(GND_net), .I1(n3151), .I2(VCC_net), 
            .I3(n28678), .O(n3218)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_10 (.CI(n28678), .I0(n3151), .I1(VCC_net), 
            .CO(n28679));
    SB_LUT4 div_46_LessThan_1281_i43_2_lut (.I0(n1969), .I1(n88), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_5027));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1281_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i41_2_lut (.I0(n1970), .I1(n89), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_5026));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1281_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i39_2_lut (.I0(n1971), .I1(n90), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5025));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1281_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_3_lut_adj_1793 (.I0(n2256), .I1(n2257), .I2(n2258), .I3(GND_net), 
            .O(n36071));
    defparam i1_3_lut_adj_1793.LUT_INIT = 16'hfefe;
    SB_LUT4 div_46_LessThan_1281_i37_2_lut (.I0(n1972), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5024));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1281_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1653_7_lut (.I0(GND_net), .I1(n2454_adj_4879), .I2(GND_net), 
            .I3(n28896), .O(n2521)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_9_lut (.I0(GND_net), .I1(n3152), .I2(VCC_net), 
            .I3(n28677), .O(n3219)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_mux_3_i10_3_lut (.I0(encoder0_position[9]), .I1(n16_adj_4703), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n1057_adj_4736));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1794 (.I0(n2248), .I1(n2250), .I2(n2253), .I3(n2252), 
            .O(n26_adj_5245));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i11_4_lut_adj_1794.LUT_INIT = 16'hfffe;
    SB_LUT4 add_2338_2_lut (.I0(GND_net), .I1(n919), .I2(n558), .I3(VCC_net), 
            .O(n5950)) /* synthesis syn_instantiated=1 */ ;
    defparam add_2338_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2338_2 (.CI(VCC_net), .I0(n919), .I1(n558), .CO(n28268));
    SB_LUT4 div_46_LessThan_1281_i25_2_lut (.I0(n1978), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_5014));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1281_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i27_2_lut (.I0(n1977), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5016));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1281_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut (.I0(control_mode[0]), .I1(n15942), .I2(control_mode[1]), 
            .I3(GND_net), .O(n15_adj_4673));   // verilog/TinyFPGA_B.v(210[5:22])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_46_LessThan_1281_i29_2_lut (.I0(n1976), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5018));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1281_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_adj_1795 (.I0(control_mode[0]), .I1(n15942), 
            .I2(control_mode[1]), .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(210[5:22])
    defparam i1_2_lut_3_lut_adj_1795.LUT_INIT = 16'hefef;
    SB_LUT4 div_46_LessThan_1281_i31_2_lut (.I0(n1975), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5020));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1281_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i33_2_lut (.I0(n1974), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5021));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1281_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1281_i35_2_lut (.I0(n1973), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5023));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1281_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1283_1_lut (.I0(n1991), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1992));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1283_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1281_i23_2_lut (.I0(n1979), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_5012));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1281_i23_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1796 (.I0(n2254), .I1(n2246), .I2(n36071), .I3(n2255), 
            .O(n19_adj_5247));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i4_4_lut_adj_1796.LUT_INIT = 16'heccc;
    SB_LUT4 i34543_4_lut (.I0(n29_adj_5018), .I1(n27_adj_5016), .I2(n25_adj_5014), 
            .I3(n23_adj_5012), .O(n41390));
    defparam i34543_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34528_4_lut (.I0(n35_adj_5023), .I1(n33_adj_5021), .I2(n31_adj_5020), 
            .I3(n41390), .O(n41375));
    defparam i34528_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1281_i22_4_lut (.I0(n1057_adj_4736), .I1(n99), 
            .I2(n1980), .I3(n558), .O(n22_adj_5011));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1281_i22_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_1281_i30_3_lut (.I0(n28_adj_5017), .I1(n93), 
            .I2(n33_adj_5021), .I3(GND_net), .O(n30_adj_5019));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1281_i30_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i1_3_lut_4_lut (.I0(n99), .I1(n16003), .I2(n558), .I3(n224), 
            .O(n5_adj_5242));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h02ff;
    SB_LUT4 div_46_LessThan_1281_i34_3_lut (.I0(n26_adj_5015), .I1(n91), 
            .I2(n37_adj_5024), .I3(GND_net), .O(n34_adj_5022));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1281_i34_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i2_3_lut_4_lut_adj_1797 (.I0(n99), .I1(n16003), .I2(n224), 
            .I3(n558), .O(n248));
    defparam i2_3_lut_4_lut_adj_1797.LUT_INIT = 16'hdddf;
    SB_LUT4 i35876_4_lut (.I0(n34_adj_5022), .I1(n24_adj_5013), .I2(n37_adj_5024), 
            .I3(n41368), .O(n42723));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35876_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34532_3_lut_3_lut (.I0(n392), .I1(n558), .I2(n369), .I3(GND_net), 
            .O(n510));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34532_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_CARRY rem_4_add_2122_9 (.CI(n28677), .I0(n3152), .I1(VCC_net), 
            .CO(n28678));
    SB_LUT4 i35877_3_lut (.I0(n42723), .I1(n90), .I2(n39_adj_5025), .I3(GND_net), 
            .O(n42724));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35877_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35722_3_lut (.I0(n42724), .I1(n89), .I2(n41_adj_5026), .I3(GND_net), 
            .O(n42569));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35722_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35659_4_lut (.I0(n41_adj_5026), .I1(n39_adj_5025), .I2(n37_adj_5024), 
            .I3(n41375), .O(n42506));
    defparam i35659_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35864_4_lut (.I0(n30_adj_5019), .I1(n22_adj_5011), .I2(n33_adj_5021), 
            .I3(n41385), .O(n42711));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35864_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34871_3_lut (.I0(n42569), .I1(n88), .I2(n43_adj_5027), .I3(GND_net), 
            .O(n41718));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34871_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i274_4_lut_4_lut (.I0(n392), .I1(n99), .I2(n2_adj_5323), 
            .I3(n5_adj_5242), .O(n35676));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i274_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i34537_3_lut_3_lut (.I0(n533), .I1(n558), .I2(n511), .I3(GND_net), 
            .O(n649));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34537_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 i1_2_lut_adj_1798 (.I0(n2241), .I1(n2240), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_5248));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i1_2_lut_adj_1798.LUT_INIT = 16'heeee;
    SB_LUT4 i35949_4_lut (.I0(n41718), .I1(n42711), .I2(n43_adj_5027), 
            .I3(n42506), .O(n42796));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35949_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35950_3_lut (.I0(n42796), .I1(n87), .I2(n1968), .I3(GND_net), 
            .O(n42797));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35950_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_46_i367_4_lut_4_lut (.I0(n533), .I1(n98), .I2(n4_adj_5252), 
            .I3(n35676), .O(n35825));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i367_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i1_4_lut_adj_1799 (.I0(n42797), .I1(n15980), .I2(n86), .I3(n1967), 
            .O(n1991));
    defparam i1_4_lut_adj_1799.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i368_4_lut_4_lut (.I0(n533), .I1(n99), .I2(n2_adj_5268), 
            .I3(n510), .O(n648));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i368_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_46_LessThan_1210_i35_2_lut (.I0(n1868), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_5007));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1210_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i11_3_lut (.I0(encoder0_position[10]), .I1(n15_adj_4709), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n1056_adj_4735));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_1210_i33_2_lut (.I0(n1869), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_5006));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1210_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i39_2_lut (.I0(n1866), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_5010));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1210_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i37_2_lut (.I0(n1867), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_5009));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1210_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i9_4_lut_adj_1800 (.I0(n2242), .I1(n2244), .I2(n2243), .I3(n2245), 
            .O(n24_adj_5246));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i9_4_lut_adj_1800.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_1210_i27_2_lut (.I0(n1872), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_5000));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1210_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i29_2_lut (.I0(n1871), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_5002));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1210_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1210_i31_2_lut (.I0(n1870), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_5004));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1210_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i34542_3_lut_3_lut (.I0(n671), .I1(n558), .I2(n650), .I3(GND_net), 
            .O(n785));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34542_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_LUT4 div_46_i459_4_lut_4_lut (.I0(n671), .I1(n98), .I2(n4_adj_5269), 
            .I3(n648), .O(n783));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i459_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_46_i1212_1_lut (.I0(n1886), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1887));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1212_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1210_i25_2_lut (.I0(n1873), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_4998));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1210_i25_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i34605_4_lut (.I0(n31_adj_5004), .I1(n29_adj_5002), .I2(n27_adj_5000), 
            .I3(n25_adj_4998), .O(n41452));
    defparam i34605_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY rem_4_add_1653_7 (.CI(n28896), .I0(n2454_adj_4879), .I1(GND_net), 
            .CO(n28897));
    SB_LUT4 rem_4_add_1653_6_lut (.I0(GND_net), .I1(n2455_adj_4878), .I2(GND_net), 
            .I3(n28895), .O(n2522)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_6 (.CI(n28895), .I0(n2455_adj_4878), .I1(GND_net), 
            .CO(n28896));
    SB_LUT4 rem_4_add_2122_8_lut (.I0(GND_net), .I1(n3153), .I2(VCC_net), 
            .I3(n28676), .O(n3220)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_8 (.CI(n28676), .I0(n3153), .I1(VCC_net), 
            .CO(n28677));
    SB_LUT4 div_46_LessThan_1210_i36_3_lut (.I0(n28_adj_5001), .I1(n91), 
            .I2(n39_adj_5010), .I3(GND_net), .O(n36_adj_5008));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1210_i36_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_i460_4_lut_4_lut (.I0(n671), .I1(n99), .I2(n2_adj_5273), 
            .I3(n649), .O(n784));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i460_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 rem_4_add_2122_7_lut (.I0(GND_net), .I1(n3154), .I2(GND_net), 
            .I3(n28675), .O(n3221)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1653_5_lut (.I0(GND_net), .I1(n2456_adj_4877), .I2(VCC_net), 
            .I3(n28894), .O(n2523)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1653_5 (.CI(n28894), .I0(n2456_adj_4877), .I1(VCC_net), 
            .CO(n28895));
    SB_CARRY rem_4_add_2122_7 (.CI(n28675), .I0(n3154), .I1(GND_net), 
            .CO(n28676));
    SB_LUT4 rem_4_add_1653_4_lut (.I0(GND_net), .I1(n2457_adj_4876), .I2(VCC_net), 
            .I3(n28893), .O(n2524)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1210_i24_4_lut (.I0(n1056_adj_4735), .I1(n99), 
            .I2(n1874), .I3(n558), .O(n24_adj_4997));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1210_i24_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_1210_i32_3_lut (.I0(n30_adj_5003), .I1(n93), 
            .I2(n35_adj_5007), .I3(GND_net), .O(n32_adj_5005));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1210_i32_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34589_4_lut (.I0(n37_adj_5009), .I1(n35_adj_5007), .I2(n33_adj_5006), 
            .I3(n41452), .O(n41436));
    defparam i34589_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35884_4_lut (.I0(n36_adj_5008), .I1(n26_adj_4999), .I2(n39_adj_5010), 
            .I3(n41430), .O(n42731));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35884_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35568_4_lut (.I0(n32_adj_5005), .I1(n24_adj_4997), .I2(n35_adj_5007), 
            .I3(n41446), .O(n42415));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35568_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i36004_4_lut (.I0(n42415), .I1(n42731), .I2(n39_adj_5010), 
            .I3(n41436), .O(n42851));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36004_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36005_3_lut (.I0(n42851), .I1(n90), .I2(n1865), .I3(GND_net), 
            .O(n42852));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36005_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35956_3_lut (.I0(n42852), .I1(n89), .I2(n1864), .I3(GND_net), 
            .O(n42803));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35956_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_46_i458_4_lut_4_lut (.I0(n671), .I1(n97), .I2(n6_adj_5253), 
            .I3(n35825), .O(n35865));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i458_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i35570_3_lut (.I0(n42803), .I1(n88), .I2(n1863), .I3(GND_net), 
            .O(n42417));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35570_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1801 (.I0(n42417), .I1(n15893), .I2(n87), .I3(n1862), 
            .O(n1886));
    defparam i1_4_lut_adj_1801.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i550_4_lut_4_lut (.I0(n806), .I1(n99), .I2(n2), .I3(n785), 
            .O(n917));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i550_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 i13_4_lut_adj_1802 (.I0(n19_adj_5247), .I1(n26_adj_5245), .I2(n2247), 
            .I3(n2251), .O(n28_adj_5244));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i13_4_lut_adj_1802.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i547_4_lut_4_lut (.I0(n806), .I1(n96), .I2(n8_adj_4669), 
            .I3(n35865), .O(n914));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i547_4_lut_4_lut.LUT_INIT = 16'h14eb;
    SB_LUT4 div_46_LessThan_1137_i37_2_lut (.I0(n1759), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4993));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1137_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i34561_3_lut_3_lut (.I0(n806), .I1(n558), .I2(n786), .I3(GND_net), 
            .O(n918));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34561_3_lut_3_lut.LUT_INIT = 16'he1e1;
    SB_CARRY rem_4_add_1653_4 (.CI(n28893), .I0(n2457_adj_4876), .I1(VCC_net), 
            .CO(n28894));
    SB_LUT4 rem_4_add_2122_6_lut (.I0(GND_net), .I1(n3155), .I2(GND_net), 
            .I3(n28674), .O(n3222)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_6 (.CI(n28674), .I0(n3155), .I1(GND_net), 
            .CO(n28675));
    SB_LUT4 rem_4_add_1653_3_lut (.I0(GND_net), .I1(n2458_adj_4875), .I2(GND_net), 
            .I3(n28892), .O(n2525)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1653_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2122_5_lut (.I0(GND_net), .I1(n3156), .I2(VCC_net), 
            .I3(n28673), .O(n3223)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1137_i35_2_lut (.I0(n1760), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4992));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1137_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i12_3_lut (.I0(encoder0_position[11]), .I1(n14_adj_4710), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n1055_adj_4734));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1653_3 (.CI(n28892), .I0(n2458_adj_4875), .I1(GND_net), 
            .CO(n28893));
    SB_CARRY rem_4_add_2122_5 (.CI(n28673), .I0(n3156), .I1(VCC_net), 
            .CO(n28674));
    SB_LUT4 div_46_i548_4_lut_4_lut (.I0(n806), .I1(n97), .I2(n6_adj_4670), 
            .I3(n783), .O(n915));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i548_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_CARRY rem_4_add_1653_2 (.CI(VCC_net), .I0(n2558_adj_4856), .I1(VCC_net), 
            .CO(n28892));
    SB_LUT4 rem_4_add_2122_4_lut (.I0(GND_net), .I1(n3157), .I2(VCC_net), 
            .I3(n28672), .O(n3224)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_24_lut (.I0(n2570), .I1(n2537_adj_4873), .I2(VCC_net), 
            .I3(n28891), .O(n2636_adj_4847)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1720_23_lut (.I0(GND_net), .I1(n2538_adj_4872), .I2(VCC_net), 
            .I3(n28890), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2122_4 (.CI(n28672), .I0(n3157), .I1(VCC_net), 
            .CO(n28673));
    SB_LUT4 rem_4_add_2122_3_lut (.I0(GND_net), .I1(n3158), .I2(GND_net), 
            .I3(n28671), .O(n3225)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2122_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_23 (.CI(n28890), .I0(n2538_adj_4872), .I1(VCC_net), 
            .CO(n28891));
    SB_LUT4 rem_4_add_1720_22_lut (.I0(GND_net), .I1(n2539_adj_4871), .I2(VCC_net), 
            .I3(n28889), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1137_i41_2_lut (.I0(n1757), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4996));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1137_i41_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_2122_3 (.CI(n28671), .I0(n3158), .I1(GND_net), 
            .CO(n28672));
    SB_DFF communication_counter_1222__i2 (.Q(communication_counter[2]), .C(LED_c), 
           .D(n163));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_CARRY rem_4_add_1720_22 (.CI(n28889), .I0(n2539_adj_4871), .I1(VCC_net), 
            .CO(n28890));
    SB_CARRY rem_4_add_2122_2 (.CI(VCC_net), .I0(n3258), .I1(VCC_net), 
            .CO(n28671));
    SB_LUT4 rem_4_add_1720_21_lut (.I0(GND_net), .I1(n2540_adj_4870), .I2(VCC_net), 
            .I3(n28888), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_31_lut (.I0(n3263), .I1(n3230), .I2(VCC_net), 
            .I3(n28670), .O(n38464)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_31_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_1720_21 (.CI(n28888), .I0(n2540_adj_4870), .I1(VCC_net), 
            .CO(n28889));
    SB_LUT4 div_46_LessThan_1137_i39_2_lut (.I0(n1758), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4995));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1137_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_1720_20_lut (.I0(GND_net), .I1(n2541_adj_4869), .I2(VCC_net), 
            .I3(n28887), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_30_lut (.I0(GND_net), .I1(n3231), .I2(VCC_net), 
            .I3(n28669), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_30 (.CI(n28669), .I0(n3231), .I1(VCC_net), 
            .CO(n28670));
    SB_CARRY rem_4_add_1720_20 (.CI(n28887), .I0(n2541_adj_4869), .I1(VCC_net), 
            .CO(n28888));
    SB_LUT4 rem_4_add_2189_29_lut (.I0(GND_net), .I1(n3232), .I2(VCC_net), 
            .I3(n28668), .O(n3299)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_29_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i549_4_lut_4_lut (.I0(n806), .I1(n98), .I2(n4_adj_4672), 
            .I3(n784), .O(n916));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i549_4_lut_4_lut.LUT_INIT = 16'heb14;
    SB_LUT4 div_46_i637_3_lut_3_lut (.I0(n938), .I1(n5948), .I2(n917), 
            .I3(GND_net), .O(n1046));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i637_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1720_19_lut (.I0(GND_net), .I1(n2542_adj_4868), .I2(VCC_net), 
            .I3(n28886), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_29 (.CI(n28668), .I0(n3232), .I1(VCC_net), 
            .CO(n28669));
    SB_LUT4 div_46_LessThan_1137_i29_2_lut (.I0(n1763), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4988));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1137_i29_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1720_19 (.CI(n28886), .I0(n2542_adj_4868), .I1(VCC_net), 
            .CO(n28887));
    SB_LUT4 rem_4_add_2189_28_lut (.I0(GND_net), .I1(n3233), .I2(VCC_net), 
            .I3(n28667), .O(n3300)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_18_lut (.I0(GND_net), .I1(n2543_adj_4867), .I2(VCC_net), 
            .I3(n28885), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_28 (.CI(n28667), .I0(n3233), .I1(VCC_net), 
            .CO(n28668));
    SB_LUT4 div_46_LessThan_1137_i31_2_lut (.I0(n1762), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4990));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1137_i31_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1720_18 (.CI(n28885), .I0(n2543_adj_4867), .I1(VCC_net), 
            .CO(n28886));
    SB_LUT4 rem_4_add_2189_27_lut (.I0(GND_net), .I1(n3234), .I2(VCC_net), 
            .I3(n28666), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_17_lut (.I0(GND_net), .I1(n2544_adj_4866), .I2(VCC_net), 
            .I3(n28884), .O(n2611)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_27 (.CI(n28666), .I0(n3234), .I1(VCC_net), 
            .CO(n28667));
    SB_LUT4 div_46_LessThan_1137_i33_2_lut (.I0(n1761), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4991));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1137_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1139_1_lut (.I0(n1778), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1779));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1139_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY rem_4_add_1720_17 (.CI(n28884), .I0(n2544_adj_4866), .I1(VCC_net), 
            .CO(n28885));
    SB_LUT4 rem_4_add_2189_26_lut (.I0(GND_net), .I1(n3235), .I2(VCC_net), 
            .I3(n28665), .O(n3302)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_26_lut.LUT_INIT = 16'hC33C;
    SB_DFF communication_counter_1222__i3 (.Q(communication_counter[3]), .C(LED_c), 
           .D(n162));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i4 (.Q(communication_counter[4]), .C(LED_c), 
           .D(n161));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i5 (.Q(communication_counter[5]), .C(LED_c), 
           .D(n160));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i6 (.Q(communication_counter[6]), .C(LED_c), 
           .D(n159));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i7 (.Q(communication_counter[7]), .C(LED_c), 
           .D(n158));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i8 (.Q(communication_counter[8]), .C(LED_c), 
           .D(n157));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i9 (.Q(communication_counter[9]), .C(LED_c), 
           .D(n156));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i10 (.Q(communication_counter[10]), 
           .C(LED_c), .D(n155));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i11 (.Q(communication_counter[11]), 
           .C(LED_c), .D(n154));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i12 (.Q(communication_counter[12]), 
           .C(LED_c), .D(n153));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i13 (.Q(communication_counter[13]), 
           .C(LED_c), .D(n152));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i14 (.Q(communication_counter[14]), 
           .C(LED_c), .D(n151));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i15 (.Q(communication_counter[15]), 
           .C(LED_c), .D(n150));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i16 (.Q(communication_counter[16]), 
           .C(LED_c), .D(n149));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i17 (.Q(communication_counter[17]), 
           .C(LED_c), .D(n148));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i18 (.Q(communication_counter[18]), 
           .C(LED_c), .D(n147));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i19 (.Q(communication_counter[19]), 
           .C(LED_c), .D(n146));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i20 (.Q(communication_counter[20]), 
           .C(LED_c), .D(n145));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i21 (.Q(communication_counter[21]), 
           .C(LED_c), .D(n144));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i22 (.Q(communication_counter[22]), 
           .C(LED_c), .D(n143));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i23 (.Q(communication_counter[23]), 
           .C(LED_c), .D(n142));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i24 (.Q(communication_counter[24]), 
           .C(LED_c), .D(n141));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i25 (.Q(communication_counter[25]), 
           .C(LED_c), .D(n140));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i26 (.Q(communication_counter[26]), 
           .C(LED_c), .D(n139));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i27 (.Q(communication_counter[27]), 
           .C(LED_c), .D(n138));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i28 (.Q(communication_counter[28]), 
           .C(LED_c), .D(n137));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i29 (.Q(communication_counter[29]), 
           .C(LED_c), .D(n136));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i30 (.Q(communication_counter[30]), 
           .C(LED_c), .D(n135));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_DFF communication_counter_1222__i31 (.Q(communication_counter[31]), 
           .C(LED_c), .D(n134));   // verilog/TinyFPGA_B.v(52[28:51])
    SB_LUT4 rem_4_add_715_8_lut (.I0(n1085), .I1(n1052), .I2(VCC_net), 
            .I3(n28227), .O(n1151)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 div_46_LessThan_1137_i27_2_lut (.I0(n1764), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_4986));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1137_i27_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 rem_4_add_715_7_lut (.I0(GND_net), .I1(n1053), .I2(VCC_net), 
            .I3(n28226), .O(n1120)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_26 (.CI(n28665), .I0(n3235), .I1(VCC_net), 
            .CO(n28666));
    SB_LUT4 rem_4_add_1720_16_lut (.I0(GND_net), .I1(n2545_adj_4865), .I2(VCC_net), 
            .I3(n28883), .O(n2612)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_25_lut (.I0(GND_net), .I1(n3236), .I2(VCC_net), 
            .I3(n28664), .O(n3303)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_16 (.CI(n28883), .I0(n2545_adj_4865), .I1(VCC_net), 
            .CO(n28884));
    SB_LUT4 i33934_4_lut (.I0(n33_adj_4991), .I1(n31_adj_4990), .I2(n29_adj_4988), 
            .I3(n27_adj_4986), .O(n40780));
    defparam i33934_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY rem_4_add_2189_25 (.CI(n28664), .I0(n3236), .I1(VCC_net), 
            .CO(n28665));
    SB_CARRY rem_4_add_715_7 (.CI(n28226), .I0(n1053), .I1(VCC_net), .CO(n28227));
    SB_LUT4 rem_4_add_715_6_lut (.I0(GND_net), .I1(n1054), .I2(GND_net), 
            .I3(n28225), .O(n1121)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_6 (.CI(n28225), .I0(n1054), .I1(GND_net), .CO(n28226));
    SB_LUT4 rem_4_add_715_5_lut (.I0(GND_net), .I1(n1055), .I2(GND_net), 
            .I3(n28224), .O(n1122)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_5 (.CI(n28224), .I0(n1055), .I1(GND_net), .CO(n28225));
    SB_LUT4 rem_4_add_715_4_lut (.I0(GND_net), .I1(n1056), .I2(VCC_net), 
            .I3(n28223), .O(n1123)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i639_3_lut_3_lut (.I0(n938), .I1(n5950), .I2(n919), 
            .I3(GND_net), .O(n1048));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i639_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_715_4 (.CI(n28223), .I0(n1056), .I1(VCC_net), .CO(n28224));
    SB_LUT4 rem_4_add_715_3_lut (.I0(GND_net), .I1(n1057), .I2(VCC_net), 
            .I3(n28222), .O(n1124)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1137_i38_3_lut (.I0(n30_adj_4989), .I1(n91), 
            .I2(n41_adj_4996), .I3(GND_net), .O(n38_adj_4994));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1137_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1137_i26_4_lut (.I0(n1055_adj_4734), .I1(n99), 
            .I2(n1765), .I3(n558), .O(n26_adj_4985));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1137_i26_4_lut.LUT_INIT = 16'h0317;
    SB_CARRY rem_4_add_715_3 (.CI(n28222), .I0(n1057), .I1(VCC_net), .CO(n28223));
    SB_LUT4 rem_4_add_715_2_lut (.I0(GND_net), .I1(n1058), .I2(GND_net), 
            .I3(VCC_net), .O(n1125)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_715_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_715_2 (.CI(VCC_net), .I0(n1058), .I1(GND_net), 
            .CO(n28222));
    SB_LUT4 div_46_i638_3_lut_3_lut (.I0(n938), .I1(n5949), .I2(n918), 
            .I3(GND_net), .O(n1047));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i638_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i636_3_lut_3_lut (.I0(n938), .I1(n5947), .I2(n916), 
            .I3(GND_net), .O(n1045));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i636_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i634_3_lut_3_lut (.I0(n938), .I1(n5945), .I2(n914), 
            .I3(GND_net), .O(n1043));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i634_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_2189_24_lut (.I0(GND_net), .I1(n3237), .I2(VCC_net), 
            .I3(n28663), .O(n3304)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35746_3_lut (.I0(n26_adj_4985), .I1(n95), .I2(n33_adj_4991), 
            .I3(GND_net), .O(n42593));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35746_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_add_916_11_lut (.I0(n1382), .I1(n1349), .I2(VCC_net), 
            .I3(n28213), .O(n1448)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_916_10_lut (.I0(GND_net), .I1(n1350), .I2(VCC_net), 
            .I3(n28212), .O(n1417)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_10 (.CI(n28212), .I0(n1350), .I1(VCC_net), 
            .CO(n28213));
    SB_LUT4 i35747_3_lut (.I0(n42593), .I1(n94), .I2(n35_adj_4992), .I3(GND_net), 
            .O(n42594));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35747_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33926_4_lut (.I0(n39_adj_4995), .I1(n37_adj_4993), .I2(n35_adj_4992), 
            .I3(n40780), .O(n40772));
    defparam i33926_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35941_4_lut (.I0(n38_adj_4994), .I1(n28_adj_4987), .I2(n41_adj_4996), 
            .I3(n40768), .O(n42788));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35941_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 rem_4_add_1720_15_lut (.I0(GND_net), .I1(n2546_adj_4864), .I2(VCC_net), 
            .I3(n28882), .O(n2613)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_24 (.CI(n28663), .I0(n3237), .I1(VCC_net), 
            .CO(n28664));
    SB_LUT4 div_46_i635_3_lut_3_lut (.I0(n938), .I1(n5946), .I2(n915), 
            .I3(GND_net), .O(n1044));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i635_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_2189_23_lut (.I0(GND_net), .I1(n3238), .I2(VCC_net), 
            .I3(n28662), .O(n3305)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35565_3_lut (.I0(n42594), .I1(n93), .I2(n37_adj_4993), .I3(GND_net), 
            .O(n42412));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35565_3_lut.LUT_INIT = 16'h3a3a;
    SB_CARRY rem_4_add_2189_23 (.CI(n28662), .I0(n3238), .I1(VCC_net), 
            .CO(n28663));
    SB_LUT4 rem_4_add_916_9_lut (.I0(GND_net), .I1(n1351), .I2(VCC_net), 
            .I3(n28211), .O(n1418)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_15 (.CI(n28882), .I0(n2546_adj_4864), .I1(VCC_net), 
            .CO(n28883));
    SB_LUT4 rem_4_add_1720_14_lut (.I0(GND_net), .I1(n2547_adj_4863), .I2(VCC_net), 
            .I3(n28881), .O(n2614)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_22_lut (.I0(GND_net), .I1(n3239), .I2(VCC_net), 
            .I3(n28661), .O(n3306)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_22 (.CI(n28661), .I0(n3239), .I1(VCC_net), 
            .CO(n28662));
    SB_CARRY rem_4_add_916_9 (.CI(n28211), .I0(n1351), .I1(VCC_net), .CO(n28212));
    SB_CARRY rem_4_add_1720_14 (.CI(n28881), .I0(n2547_adj_4863), .I1(VCC_net), 
            .CO(n28882));
    SB_LUT4 rem_4_add_1720_13_lut (.I0(GND_net), .I1(n2548_adj_4862), .I2(VCC_net), 
            .I3(n28880), .O(n2615)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_21_lut (.I0(GND_net), .I1(n3240), .I2(VCC_net), 
            .I3(n28660), .O(n3307)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_13 (.CI(n28880), .I0(n2548_adj_4862), .I1(VCC_net), 
            .CO(n28881));
    SB_LUT4 rem_4_add_1720_12_lut (.I0(GND_net), .I1(n2549_adj_4861), .I2(VCC_net), 
            .I3(n28879), .O(n2616)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_21 (.CI(n28660), .I0(n3240), .I1(VCC_net), 
            .CO(n28661));
    SB_LUT4 rem_4_add_2189_20_lut (.I0(GND_net), .I1(n3241), .I2(VCC_net), 
            .I3(n28659), .O(n3308)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_916_8_lut (.I0(GND_net), .I1(n1352), .I2(VCC_net), 
            .I3(n28210), .O(n1419)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36020_4_lut (.I0(n42412), .I1(n42788), .I2(n41_adj_4996), 
            .I3(n40772), .O(n42867));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36020_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY rem_4_add_1720_12 (.CI(n28879), .I0(n2549_adj_4861), .I1(VCC_net), 
            .CO(n28880));
    SB_CARRY rem_4_add_2189_20 (.CI(n28659), .I0(n3241), .I1(VCC_net), 
            .CO(n28660));
    SB_CARRY rem_4_add_916_8 (.CI(n28210), .I0(n1352), .I1(VCC_net), .CO(n28211));
    SB_LUT4 rem_4_add_1720_11_lut (.I0(GND_net), .I1(n2550_adj_4860), .I2(VCC_net), 
            .I3(n28878), .O(n2617)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_11 (.CI(n28878), .I0(n2550_adj_4860), .I1(VCC_net), 
            .CO(n28879));
    SB_LUT4 rem_4_add_2189_19_lut (.I0(GND_net), .I1(n3242), .I2(VCC_net), 
            .I3(n28658), .O(n3309)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_19 (.CI(n28658), .I0(n3242), .I1(VCC_net), 
            .CO(n28659));
    SB_LUT4 rem_4_add_1720_10_lut (.I0(GND_net), .I1(n2551_adj_4859), .I2(VCC_net), 
            .I3(n28877), .O(n2618_adj_4855)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_18_lut (.I0(GND_net), .I1(n3243), .I2(VCC_net), 
            .I3(n28657), .O(n3310)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_18 (.CI(n28657), .I0(n3243), .I1(VCC_net), 
            .CO(n28658));
    SB_CARRY rem_4_add_1720_10 (.CI(n28877), .I0(n2551_adj_4859), .I1(VCC_net), 
            .CO(n28878));
    SB_LUT4 rem_4_add_916_7_lut (.I0(GND_net), .I1(n1353), .I2(VCC_net), 
            .I3(n28209), .O(n1420_adj_4880)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_7 (.CI(n28209), .I0(n1353), .I1(VCC_net), .CO(n28210));
    SB_LUT4 i36021_3_lut (.I0(n42867), .I1(n90), .I2(n1756), .I3(GND_net), 
            .O(n42868));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36021_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35999_3_lut (.I0(n42868), .I1(n89), .I2(n1755), .I3(GND_net), 
            .O(n42846));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35999_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 rem_4_add_1720_9_lut (.I0(GND_net), .I1(n2552_adj_4858), .I2(VCC_net), 
            .I3(n28876), .O(n2619_adj_4854)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_17_lut (.I0(GND_net), .I1(n3244), .I2(VCC_net), 
            .I3(n28656), .O(n3311)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_9 (.CI(n28876), .I0(n2552_adj_4858), .I1(VCC_net), 
            .CO(n28877));
    SB_CARRY rem_4_add_2189_17 (.CI(n28656), .I0(n3244), .I1(VCC_net), 
            .CO(n28657));
    SB_LUT4 div_46_LessThan_570_i42_3_lut_3_lut (.I0(n916), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n42_adj_4822));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_570_i42_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 rem_4_add_1720_8_lut (.I0(GND_net), .I1(n2553_adj_4857), .I2(VCC_net), 
            .I3(n28875), .O(n2620_adj_4853)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_16_lut (.I0(GND_net), .I1(n3245), .I2(VCC_net), 
            .I3(n28655), .O(n3312)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_16 (.CI(n28655), .I0(n3245), .I1(VCC_net), 
            .CO(n28656));
    SB_LUT4 rem_4_add_916_6_lut (.I0(GND_net), .I1(n1354), .I2(GND_net), 
            .I3(n28208), .O(n1421)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_8 (.CI(n28875), .I0(n2553_adj_4857), .I1(VCC_net), 
            .CO(n28876));
    SB_LUT4 rem_4_add_2189_15_lut (.I0(GND_net), .I1(n3246), .I2(VCC_net), 
            .I3(n28654), .O(n3313)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_15 (.CI(n28654), .I0(n3246), .I1(VCC_net), 
            .CO(n28655));
    SB_LUT4 i34103_3_lut_4_lut (.I0(n916), .I1(n97), .I2(n98), .I3(n917), 
            .O(n40949));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34103_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 rem_4_add_1720_7_lut (.I0(GND_net), .I1(n2554), .I2(GND_net), 
            .I3(n28874), .O(n2621_adj_4852)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_7 (.CI(n28874), .I0(n2554), .I1(GND_net), 
            .CO(n28875));
    SB_LUT4 rem_4_add_1720_6_lut (.I0(GND_net), .I1(n2555), .I2(GND_net), 
            .I3(n28873), .O(n2622_adj_4851)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_2189_14_lut (.I0(GND_net), .I1(n3247), .I2(VCC_net), 
            .I3(n28653), .O(n3314)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_6 (.CI(n28208), .I0(n1354), .I1(GND_net), .CO(n28209));
    SB_CARRY rem_4_add_2189_14 (.CI(n28653), .I0(n3247), .I1(VCC_net), 
            .CO(n28654));
    SB_CARRY rem_4_add_1720_6 (.CI(n28873), .I0(n2555), .I1(GND_net), 
            .CO(n28874));
    SB_LUT4 rem_4_add_2189_13_lut (.I0(GND_net), .I1(n3248), .I2(VCC_net), 
            .I3(n28652), .O(n3315)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1803 (.I0(n42846), .I1(n15977), .I2(n88), .I3(n1754), 
            .O(n1778));
    defparam i1_4_lut_adj_1803.LUT_INIT = 16'hceef;
    SB_LUT4 rem_4_add_916_5_lut (.I0(GND_net), .I1(n1355), .I2(GND_net), 
            .I3(n28207), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_5_lut (.I0(GND_net), .I1(n2556), .I2(VCC_net), 
            .I3(n28872), .O(n2623_adj_4850)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_5 (.CI(n28872), .I0(n2556), .I1(VCC_net), 
            .CO(n28873));
    SB_CARRY rem_4_add_2189_13 (.CI(n28652), .I0(n3248), .I1(VCC_net), 
            .CO(n28653));
    SB_LUT4 rem_4_add_2189_12_lut (.I0(GND_net), .I1(n3249), .I2(VCC_net), 
            .I3(n28651), .O(n3316)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1720_4_lut (.I0(GND_net), .I1(n2557), .I2(VCC_net), 
            .I3(n28871), .O(n2624_adj_4849)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_12 (.CI(n28651), .I0(n3249), .I1(VCC_net), 
            .CO(n28652));
    SB_CARRY rem_4_add_916_5 (.CI(n28207), .I0(n1355), .I1(GND_net), .CO(n28208));
    SB_LUT4 rem_4_add_2189_11_lut (.I0(GND_net), .I1(n3250), .I2(VCC_net), 
            .I3(n28650), .O(n3317)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_916_4_lut (.I0(GND_net), .I1(n1356), .I2(VCC_net), 
            .I3(n28206), .O(n1423)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_4 (.CI(n28871), .I0(n2557), .I1(VCC_net), 
            .CO(n28872));
    SB_CARRY rem_4_add_2189_11 (.CI(n28650), .I0(n3250), .I1(VCC_net), 
            .CO(n28651));
    SB_CARRY rem_4_add_916_4 (.CI(n28206), .I0(n1356), .I1(VCC_net), .CO(n28207));
    SB_LUT4 rem_4_add_2189_10_lut (.I0(GND_net), .I1(n3251), .I2(VCC_net), 
            .I3(n28649), .O(n3318)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_916_3_lut (.I0(GND_net), .I1(n1357), .I2(VCC_net), 
            .I3(n28205), .O(n1424)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_3 (.CI(n28205), .I0(n1357), .I1(VCC_net), .CO(n28206));
    SB_LUT4 rem_4_add_1720_3_lut (.I0(GND_net), .I1(n2558_adj_4856), .I2(GND_net), 
            .I3(n28870), .O(n2625_adj_4848)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1720_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_10 (.CI(n28649), .I0(n3251), .I1(VCC_net), 
            .CO(n28650));
    SB_LUT4 rem_4_add_916_2_lut (.I0(GND_net), .I1(n1358), .I2(GND_net), 
            .I3(VCC_net), .O(n1425)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_916_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_916_2 (.CI(VCC_net), .I0(n1358), .I1(GND_net), 
            .CO(n28205));
    SB_CARRY rem_4_add_1720_3 (.CI(n28870), .I0(n2558_adj_4856), .I1(GND_net), 
            .CO(n28871));
    SB_LUT4 rem_4_add_2189_9_lut (.I0(GND_net), .I1(n3252), .I2(VCC_net), 
            .I3(n28648), .O(n3319)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1720_2 (.CI(VCC_net), .I0(n2658), .I1(VCC_net), 
            .CO(n28870));
    SB_CARRY rem_4_add_2189_9 (.CI(n28648), .I0(n3252), .I1(VCC_net), 
            .CO(n28649));
    SB_LUT4 rem_4_add_1787_25_lut (.I0(n2669), .I1(n2636_adj_4847), .I2(VCC_net), 
            .I3(n28869), .O(n2735)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_2189_8_lut (.I0(GND_net), .I1(n3253), .I2(VCC_net), 
            .I3(n28647), .O(n3320)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_8_lut.LUT_INIT = 16'hC33C;
    GND i1 (.Y(GND_net));
    SB_LUT4 rem_4_add_1787_24_lut (.I0(GND_net), .I1(n2637_adj_4846), .I2(VCC_net), 
            .I3(n28868), .O(n2704_adj_4841)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_8 (.CI(n28647), .I0(n3253), .I1(VCC_net), 
            .CO(n28648));
    SB_CARRY rem_4_add_1787_24 (.CI(n28868), .I0(n2637_adj_4846), .I1(VCC_net), 
            .CO(n28869));
    SB_LUT4 rem_4_add_2189_7_lut (.I0(GND_net), .I1(n3254), .I2(GND_net), 
            .I3(n28646), .O(n3321)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_23_lut (.I0(GND_net), .I1(n2638_adj_4845), .I2(VCC_net), 
            .I3(n28867), .O(n2705_adj_4840)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_7 (.CI(n28646), .I0(n3254), .I1(GND_net), 
            .CO(n28647));
    SB_CARRY rem_4_add_1787_23 (.CI(n28867), .I0(n2638_adj_4845), .I1(VCC_net), 
            .CO(n28868));
    SB_LUT4 rem_4_add_2189_6_lut (.I0(GND_net), .I1(n3255), .I2(GND_net), 
            .I3(n28645), .O(n3322)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_22_lut (.I0(GND_net), .I1(n2639), .I2(VCC_net), 
            .I3(n28866), .O(n2706_adj_4839)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_6 (.CI(n28645), .I0(n3255), .I1(GND_net), 
            .CO(n28646));
    SB_LUT4 rem_4_add_2189_5_lut (.I0(GND_net), .I1(n3256), .I2(VCC_net), 
            .I3(n28644), .O(n3323)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_22 (.CI(n28866), .I0(n2639), .I1(VCC_net), 
            .CO(n28867));
    SB_LUT4 rem_4_unary_minus_2_add_3_33_lut (.I0(communication_counter[31]), 
            .I1(GND_net), .I2(n2_adj_5275), .I3(n29892), .O(n746)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_unary_minus_2_add_3_32_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_5276), .I3(n29891), .O(n3_adj_4806)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_32 (.CI(n29891), .I0(GND_net), .I1(n3_adj_5276), 
            .CO(n29892));
    SB_LUT4 rem_4_add_1787_21_lut (.I0(GND_net), .I1(n2640), .I2(VCC_net), 
            .I3(n28865), .O(n2707_adj_4838)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_5 (.CI(n28644), .I0(n3256), .I1(VCC_net), 
            .CO(n28645));
    SB_LUT4 rem_4_unary_minus_2_add_3_31_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_5277), .I3(n29890), .O(n4_adj_4805)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_31 (.CI(n29890), .I0(GND_net), .I1(n4_adj_5277), 
            .CO(n29891));
    SB_LUT4 rem_4_unary_minus_2_add_3_30_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_5278), .I3(n29889), .O(n5_adj_4804)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_30 (.CI(n29889), .I0(GND_net), .I1(n5_adj_5278), 
            .CO(n29890));
    SB_LUT4 rem_4_unary_minus_2_add_3_29_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_5279), .I3(n29888), .O(n6_adj_4803)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_21 (.CI(n28865), .I0(n2640), .I1(VCC_net), 
            .CO(n28866));
    SB_CARRY rem_4_unary_minus_2_add_3_29 (.CI(n29888), .I0(GND_net), .I1(n6_adj_5279), 
            .CO(n29889));
    SB_LUT4 rem_4_add_2189_4_lut (.I0(GND_net), .I1(n3257), .I2(VCC_net), 
            .I3(n28643), .O(n3324)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_20_lut (.I0(GND_net), .I1(n2641), .I2(VCC_net), 
            .I3(n28864), .O(n2708_adj_4837)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_4 (.CI(n28643), .I0(n3257), .I1(VCC_net), 
            .CO(n28644));
    SB_LUT4 rem_4_unary_minus_2_add_3_28_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_5280), .I3(n29887), .O(n7_adj_4802)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_28 (.CI(n29887), .I0(GND_net), .I1(n7_adj_5280), 
            .CO(n29888));
    SB_LUT4 rem_4_unary_minus_2_add_3_27_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n8_adj_5281), .I3(n29886), .O(n8_adj_4801)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_20 (.CI(n28864), .I0(n2641), .I1(VCC_net), 
            .CO(n28865));
    SB_LUT4 rem_4_add_2189_3_lut (.I0(GND_net), .I1(n3258), .I2(GND_net), 
            .I3(n28642), .O(n3325)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2189_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_27 (.CI(n29886), .I0(GND_net), .I1(n8_adj_5281), 
            .CO(n29887));
    SB_CARRY rem_4_add_2189_3 (.CI(n28642), .I0(n3258), .I1(GND_net), 
            .CO(n28643));
    SB_LUT4 rem_4_unary_minus_2_add_3_26_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n9_adj_5282), .I3(n29885), .O(n9_adj_4800)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_26 (.CI(n29885), .I0(GND_net), .I1(n9_adj_5282), 
            .CO(n29886));
    SB_LUT4 rem_4_unary_minus_2_add_3_25_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n10_adj_5283), .I3(n29884), .O(n10_adj_4799)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_25 (.CI(n29884), .I0(GND_net), .I1(n10_adj_5283), 
            .CO(n29885));
    SB_LUT4 rem_4_unary_minus_2_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n11_adj_5284), .I3(n29883), .O(n11_adj_4798)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_24 (.CI(n29883), .I0(GND_net), .I1(n11_adj_5284), 
            .CO(n29884));
    SB_LUT4 rem_4_add_1787_19_lut (.I0(GND_net), .I1(n2642_adj_4844), .I2(VCC_net), 
            .I3(n28863), .O(n2709_adj_4836)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n12_adj_5285), .I3(n29882), .O(n12_adj_4797)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2189_2 (.CI(VCC_net), .I0(n3358), .I1(VCC_net), 
            .CO(n28642));
    SB_CARRY rem_4_unary_minus_2_add_3_23 (.CI(n29882), .I0(GND_net), .I1(n12_adj_5285), 
            .CO(n29883));
    SB_LUT4 rem_4_unary_minus_2_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n13_adj_5286), .I3(n29881), .O(n13_adj_4796)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_22 (.CI(n29881), .I0(GND_net), .I1(n13_adj_5286), 
            .CO(n29882));
    SB_LUT4 rem_4_unary_minus_2_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n14_adj_5287), .I3(n29880), .O(n14_adj_4795)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_19 (.CI(n28863), .I0(n2642_adj_4844), .I1(VCC_net), 
            .CO(n28864));
    SB_LUT4 rem_4_add_1787_18_lut (.I0(GND_net), .I1(n2643_adj_4843), .I2(VCC_net), 
            .I3(n28862), .O(n2710_adj_4835)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_21 (.CI(n29880), .I0(GND_net), .I1(n14_adj_5287), 
            .CO(n29881));
    SB_LUT4 rem_4_add_2298_9_lut (.I0(n43565), .I1(n2_adj_5275), .I2(n3452), 
            .I3(n28641), .O(color_23__N_164[7])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_2298_8_lut (.I0(n43569), .I1(n2_adj_5275), .I2(n3453), 
            .I3(n28640), .O(color_23__N_164[6])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_unary_minus_2_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n15_adj_5288), .I3(n29879), .O(n15_adj_4794)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_18 (.CI(n28862), .I0(n2643_adj_4843), .I1(VCC_net), 
            .CO(n28863));
    SB_CARRY rem_4_add_2298_8 (.CI(n28640), .I0(n2_adj_5275), .I1(n3453), 
            .CO(n28641));
    SB_CARRY rem_4_unary_minus_2_add_3_20 (.CI(n29879), .I0(GND_net), .I1(n15_adj_5288), 
            .CO(n29880));
    SB_LUT4 rem_4_unary_minus_2_add_3_19_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n16_adj_5289), .I3(n29878), .O(n16_adj_4793)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_19 (.CI(n29878), .I0(GND_net), .I1(n16_adj_5289), 
            .CO(n29879));
    SB_LUT4 rem_4_unary_minus_2_add_3_18_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n17_adj_5290), .I3(n29877), .O(n17_adj_4792)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_17_lut (.I0(GND_net), .I1(n2644), .I2(VCC_net), 
            .I3(n28861), .O(n2711_adj_4834)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_18 (.CI(n29877), .I0(GND_net), .I1(n17_adj_5290), 
            .CO(n29878));
    SB_CARRY rem_4_add_1787_17 (.CI(n28861), .I0(n2644), .I1(VCC_net), 
            .CO(n28862));
    SB_LUT4 rem_4_add_2298_7_lut (.I0(n43572), .I1(n2_adj_5275), .I2(n3454), 
            .I3(n28639), .O(color_23__N_164[5])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_7 (.CI(n28639), .I0(n2_adj_5275), .I1(n3454), 
            .CO(n28640));
    SB_LUT4 rem_4_unary_minus_2_add_3_17_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n18_adj_5291), .I3(n29876), .O(n18_adj_4791)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_17 (.CI(n29876), .I0(GND_net), .I1(n18_adj_5291), 
            .CO(n29877));
    SB_LUT4 rem_4_unary_minus_2_add_3_16_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n19_adj_5292), .I3(n29875), .O(n19_adj_4790)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_16 (.CI(n29875), .I0(GND_net), .I1(n19_adj_5292), 
            .CO(n29876));
    SB_LUT4 rem_4_unary_minus_2_add_3_15_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n20_adj_5293), .I3(n29874), .O(n20_adj_4789)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_16_lut (.I0(GND_net), .I1(n2645), .I2(VCC_net), 
            .I3(n28860), .O(n2712_adj_4833)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_15 (.CI(n29874), .I0(GND_net), .I1(n20_adj_5293), 
            .CO(n29875));
    SB_LUT4 rem_4_add_2298_6_lut (.I0(n43575), .I1(n2_adj_5275), .I2(n3455), 
            .I3(n28638), .O(color_23__N_164[4])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_unary_minus_2_add_3_14_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n21_adj_5294), .I3(n29873), .O(n21_adj_4788)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_14 (.CI(n29873), .I0(GND_net), .I1(n21_adj_5294), 
            .CO(n29874));
    SB_LUT4 rem_4_unary_minus_2_add_3_13_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n22_adj_5295), .I3(n29872), .O(n22_adj_4787)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_13 (.CI(n29872), .I0(GND_net), .I1(n22_adj_5295), 
            .CO(n29873));
    SB_LUT4 rem_4_add_782_9_lut (.I0(n1184), .I1(n1151), .I2(VCC_net), 
            .I3(n28195), .O(n1250)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_9_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_1787_16 (.CI(n28860), .I0(n2645), .I1(VCC_net), 
            .CO(n28861));
    SB_LUT4 rem_4_unary_minus_2_add_3_12_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n23_adj_5296), .I3(n29871), .O(n23_adj_4786)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2298_6 (.CI(n28638), .I0(n2_adj_5275), .I1(n3455), 
            .CO(n28639));
    SB_CARRY rem_4_unary_minus_2_add_3_12 (.CI(n29871), .I0(GND_net), .I1(n23_adj_5296), 
            .CO(n29872));
    SB_LUT4 rem_4_add_782_8_lut (.I0(GND_net), .I1(n1152), .I2(VCC_net), 
            .I3(n28194), .O(n1219)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_11_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n24_adj_5297), .I3(n29870), .O(n24_adj_4785)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_8 (.CI(n28194), .I0(n1152), .I1(VCC_net), .CO(n28195));
    SB_CARRY rem_4_unary_minus_2_add_3_11 (.CI(n29870), .I0(GND_net), .I1(n24_adj_5297), 
            .CO(n29871));
    SB_LUT4 rem_4_add_782_7_lut (.I0(GND_net), .I1(n1153), .I2(VCC_net), 
            .I3(n28193), .O(n1220)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n25_adj_5298), .I3(n29869), .O(n25_adj_4784)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_15_lut (.I0(GND_net), .I1(n2646), .I2(VCC_net), 
            .I3(n28859), .O(n2713_adj_4832)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_7 (.CI(n28193), .I0(n1153), .I1(VCC_net), .CO(n28194));
    SB_LUT4 rem_4_add_2298_5_lut (.I0(n43578), .I1(n2_adj_5275), .I2(n3456), 
            .I3(n28637), .O(color_23__N_164[3])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_5_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_782_6_lut (.I0(GND_net), .I1(n1154), .I2(GND_net), 
            .I3(n28192), .O(n1221)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_6 (.CI(n28192), .I0(n1154), .I1(GND_net), .CO(n28193));
    SB_LUT4 rem_4_add_782_5_lut (.I0(GND_net), .I1(n1155), .I2(GND_net), 
            .I3(n28191), .O(n1222)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_5 (.CI(n28191), .I0(n1155), .I1(GND_net), .CO(n28192));
    SB_LUT4 rem_4_add_782_4_lut (.I0(GND_net), .I1(n1156), .I2(VCC_net), 
            .I3(n28190), .O(n1223)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_15 (.CI(n28859), .I0(n2646), .I1(VCC_net), 
            .CO(n28860));
    SB_CARRY rem_4_unary_minus_2_add_3_10 (.CI(n29869), .I0(GND_net), .I1(n25_adj_5298), 
            .CO(n29870));
    SB_CARRY rem_4_add_2298_5 (.CI(n28637), .I0(n2_adj_5275), .I1(n3456), 
            .CO(n28638));
    SB_LUT4 rem_4_unary_minus_2_add_3_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n26_adj_5299), .I3(n29868), .O(n26_adj_4783)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_9 (.CI(n29868), .I0(GND_net), .I1(n26_adj_5299), 
            .CO(n29869));
    SB_LUT4 rem_4_unary_minus_2_add_3_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n27_adj_5300), .I3(n29867), .O(n27_adj_4782)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_8 (.CI(n29867), .I0(GND_net), .I1(n27_adj_5300), 
            .CO(n29868));
    SB_LUT4 rem_4_unary_minus_2_add_3_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n28_adj_5301), .I3(n29866), .O(n28_adj_4781)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_7 (.CI(n29866), .I0(GND_net), .I1(n28_adj_5301), 
            .CO(n29867));
    SB_LUT4 rem_4_unary_minus_2_add_3_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n29_adj_5302), .I3(n29865), .O(n29_adj_4780)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_14_lut (.I0(GND_net), .I1(n2647), .I2(VCC_net), 
            .I3(n28858), .O(n2714_adj_4831)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_6 (.CI(n29865), .I0(GND_net), .I1(n29_adj_5302), 
            .CO(n29866));
    SB_LUT4 rem_4_add_2298_4_lut (.I0(n43581), .I1(n2_adj_5275), .I2(n38575), 
            .I3(n28636), .O(color_23__N_164[2])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_782_4 (.CI(n28190), .I0(n1156), .I1(VCC_net), .CO(n28191));
    SB_LUT4 rem_4_add_782_3_lut (.I0(GND_net), .I1(n1157), .I2(VCC_net), 
            .I3(n28189), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_782_3 (.CI(n28189), .I0(n1157), .I1(VCC_net), .CO(n28190));
    SB_LUT4 rem_4_add_782_2_lut (.I0(GND_net), .I1(n1158), .I2(GND_net), 
            .I3(VCC_net), .O(n1225)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_782_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n30_adj_5303), .I3(n29864), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_5 (.CI(n29864), .I0(GND_net), .I1(n30_adj_5303), 
            .CO(n29865));
    SB_CARRY rem_4_add_782_2 (.CI(VCC_net), .I0(n1158), .I1(GND_net), 
            .CO(n28189));
    SB_LUT4 rem_4_unary_minus_2_add_3_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n31_adj_5304), .I3(n29863), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_25_lut (.I0(GND_net), .I1(displacement_23__N_229[23]), 
            .I2(n3_adj_4689), .I3(n28188), .O(displacement_23__N_80[23])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_14 (.CI(n28858), .I0(n2647), .I1(VCC_net), 
            .CO(n28859));
    SB_CARRY rem_4_unary_minus_2_add_3_4 (.CI(n29863), .I0(GND_net), .I1(n31_adj_5304), 
            .CO(n29864));
    SB_LUT4 displacement_23__I_0_add_2_24_lut (.I0(GND_net), .I1(displacement_23__N_229[22]), 
            .I2(n3_adj_4689), .I3(n28187), .O(displacement_23__N_80[22])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_2298_4 (.CI(n28636), .I0(n2_adj_5275), .I1(n38575), 
            .CO(n28637));
    SB_CARRY displacement_23__I_0_add_2_24 (.CI(n28187), .I0(displacement_23__N_229[22]), 
            .I1(n3_adj_4689), .CO(n28188));
    SB_LUT4 rem_4_unary_minus_2_add_3_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n32_adj_5305), .I3(n29862), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_3 (.CI(n29862), .I0(GND_net), .I1(n32_adj_5305), 
            .CO(n29863));
    SB_LUT4 displacement_23__I_0_add_2_23_lut (.I0(GND_net), .I1(displacement_23__N_229[21]), 
            .I2(n3_adj_4689), .I3(n28186), .O(displacement_23__N_80[21])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_unary_minus_2_add_3_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n33_adj_5306), .I3(VCC_net), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_unary_minus_2_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n33_adj_5306), 
            .CO(n29862));
    SB_LUT4 rem_4_add_2298_3_lut (.I0(communication_counter[1]), .I1(n2_adj_5275), 
            .I2(n3458), .I3(n28635), .O(color_23__N_164[1])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_3 (.CI(n28635), .I0(n2_adj_5275), .I1(n3458), 
            .CO(n28636));
    SB_LUT4 rem_4_add_1787_13_lut (.I0(GND_net), .I1(n2648), .I2(VCC_net), 
            .I3(n28857), .O(n2715_adj_4830)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_13 (.CI(n28857), .I0(n2648), .I1(VCC_net), 
            .CO(n28858));
    SB_LUT4 rem_4_add_2298_2_lut (.I0(communication_counter[0]), .I1(n2_adj_5275), 
            .I2(n3360), .I3(VCC_net), .O(color_23__N_164[0])) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_2298_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_2298_2 (.CI(VCC_net), .I0(n2_adj_5275), .I1(n3360), 
            .CO(n28635));
    SB_LUT4 rem_4_add_1787_12_lut (.I0(GND_net), .I1(n2649), .I2(VCC_net), 
            .I3(n28856), .O(n2716_adj_4829)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_23 (.CI(n28186), .I0(displacement_23__N_229[21]), 
            .I1(n3_adj_4689), .CO(n28187));
    SB_LUT4 displacement_23__I_0_add_2_22_lut (.I0(GND_net), .I1(displacement_23__N_229[20]), 
            .I2(n3_adj_4689), .I3(n28185), .O(displacement_23__N_80[20])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_22 (.CI(n28185), .I0(displacement_23__N_229[20]), 
            .I1(n3_adj_4689), .CO(n28186));
    SB_CARRY rem_4_add_1787_12 (.CI(n28856), .I0(n2649), .I1(VCC_net), 
            .CO(n28857));
    SB_LUT4 displacement_23__I_0_add_2_21_lut (.I0(GND_net), .I1(displacement_23__N_229[19]), 
            .I2(n6_adj_4683), .I3(n28184), .O(displacement_23__N_80[19])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_11_lut (.I0(GND_net), .I1(n2650), .I2(VCC_net), 
            .I3(n28855), .O(n2717_adj_4828)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_21 (.CI(n28184), .I0(displacement_23__N_229[19]), 
            .I1(n6_adj_4683), .CO(n28185));
    SB_LUT4 displacement_23__I_0_add_2_20_lut (.I0(GND_net), .I1(displacement_23__N_229[18]), 
            .I2(n7_adj_4682), .I3(n28183), .O(displacement_23__N_80[18])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_11 (.CI(n28855), .I0(n2650), .I1(VCC_net), 
            .CO(n28856));
    SB_LUT4 rem_4_add_1050_13_lut (.I0(n1580), .I1(n1547), .I2(VCC_net), 
            .I3(n29063), .O(n1646_adj_4813)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1787_10_lut (.I0(GND_net), .I1(n2651), .I2(VCC_net), 
            .I3(n28854), .O(n2718_adj_4827)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_20 (.CI(n28183), .I0(displacement_23__N_229[18]), 
            .I1(n7_adj_4682), .CO(n28184));
    SB_CARRY rem_4_add_1787_10 (.CI(n28854), .I0(n2651), .I1(VCC_net), 
            .CO(n28855));
    SB_LUT4 displacement_23__I_0_add_2_19_lut (.I0(GND_net), .I1(displacement_23__N_229[17]), 
            .I2(n8_adj_4681), .I3(n28182), .O(displacement_23__N_80[17])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_19 (.CI(n28182), .I0(displacement_23__N_229[17]), 
            .I1(n8_adj_4681), .CO(n28183));
    SB_LUT4 rem_4_add_1787_9_lut (.I0(GND_net), .I1(n2652), .I2(VCC_net), 
            .I3(n28853), .O(n2719_adj_4826)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_12_lut (.I0(GND_net), .I1(n1548), .I2(VCC_net), 
            .I3(n29062), .O(n1615)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_9 (.CI(n28853), .I0(n2652), .I1(VCC_net), 
            .CO(n28854));
    SB_LUT4 displacement_23__I_0_add_2_18_lut (.I0(GND_net), .I1(displacement_23__N_229[16]), 
            .I2(n9_adj_4677), .I3(n28181), .O(displacement_23__N_80[16])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_8_lut (.I0(GND_net), .I1(n2653), .I2(VCC_net), 
            .I3(n28852), .O(n2720_adj_4825)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_18 (.CI(n28181), .I0(displacement_23__N_229[16]), 
            .I1(n9_adj_4677), .CO(n28182));
    SB_CARRY rem_4_add_1050_12 (.CI(n29062), .I0(n1548), .I1(VCC_net), 
            .CO(n29063));
    SB_LUT4 displacement_23__I_0_add_2_17_lut (.I0(GND_net), .I1(displacement_23__N_229[15]), 
            .I2(n10_adj_4676), .I3(n28180), .O(displacement_23__N_80[15])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_11_lut (.I0(GND_net), .I1(n1549), .I2(VCC_net), 
            .I3(n29061), .O(n1616)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_8 (.CI(n28852), .I0(n2653), .I1(VCC_net), 
            .CO(n28853));
    SB_CARRY displacement_23__I_0_add_2_17 (.CI(n28180), .I0(displacement_23__N_229[15]), 
            .I1(n10_adj_4676), .CO(n28181));
    SB_LUT4 displacement_23__I_0_add_2_16_lut (.I0(GND_net), .I1(displacement_23__N_229[14]), 
            .I2(n11_adj_4664), .I3(n28179), .O(displacement_23__N_80[14])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_16 (.CI(n28179), .I0(displacement_23__N_229[14]), 
            .I1(n11_adj_4664), .CO(n28180));
    SB_LUT4 displacement_23__I_0_add_2_15_lut (.I0(GND_net), .I1(displacement_23__N_229[13]), 
            .I2(n12_adj_4716), .I3(n28178), .O(displacement_23__N_80[13])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_11 (.CI(n29061), .I0(n1549), .I1(VCC_net), 
            .CO(n29062));
    SB_LUT4 rem_4_add_1787_7_lut (.I0(GND_net), .I1(n2654), .I2(GND_net), 
            .I3(n28851), .O(n2721)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_15 (.CI(n28178), .I0(displacement_23__N_229[13]), 
            .I1(n12_adj_4716), .CO(n28179));
    SB_LUT4 displacement_23__I_0_add_2_14_lut (.I0(GND_net), .I1(displacement_23__N_229[12]), 
            .I2(n13_adj_4717), .I3(n28177), .O(displacement_23__N_80[12])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_14 (.CI(n28177), .I0(displacement_23__N_229[12]), 
            .I1(n13_adj_4717), .CO(n28178));
    SB_CARRY rem_4_add_1787_7 (.CI(n28851), .I0(n2654), .I1(GND_net), 
            .CO(n28852));
    SB_LUT4 displacement_23__I_0_add_2_13_lut (.I0(GND_net), .I1(displacement_23__N_229[11]), 
            .I2(n14_adj_4718), .I3(n28176), .O(displacement_23__N_80[11])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_13 (.CI(n28176), .I0(displacement_23__N_229[11]), 
            .I1(n14_adj_4718), .CO(n28177));
    SB_LUT4 rem_4_add_1050_10_lut (.I0(GND_net), .I1(n1550), .I2(VCC_net), 
            .I3(n29060), .O(n1617)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_12_lut (.I0(GND_net), .I1(displacement_23__N_229[10]), 
            .I2(n15_adj_4719), .I3(n28175), .O(displacement_23__N_80[10])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_10 (.CI(n29060), .I0(n1550), .I1(VCC_net), 
            .CO(n29061));
    SB_LUT4 rem_4_add_1787_6_lut (.I0(GND_net), .I1(n2655), .I2(GND_net), 
            .I3(n28850), .O(n2722)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_9_lut (.I0(GND_net), .I1(n1551), .I2(VCC_net), 
            .I3(n29059), .O(n1618)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_6 (.CI(n28850), .I0(n2655), .I1(GND_net), 
            .CO(n28851));
    SB_CARRY displacement_23__I_0_add_2_12 (.CI(n28175), .I0(displacement_23__N_229[10]), 
            .I1(n15_adj_4719), .CO(n28176));
    SB_LUT4 displacement_23__I_0_add_2_11_lut (.I0(GND_net), .I1(displacement_23__N_229[9]), 
            .I2(n16_adj_4720), .I3(n28174), .O(displacement_23__N_80[9])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_11 (.CI(n28174), .I0(displacement_23__N_229[9]), 
            .I1(n16_adj_4720), .CO(n28175));
    SB_LUT4 displacement_23__I_0_add_2_10_lut (.I0(GND_net), .I1(displacement_23__N_229[8]), 
            .I2(n17_adj_4721), .I3(n28173), .O(displacement_23__N_80[8])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_10 (.CI(n28173), .I0(displacement_23__N_229[8]), 
            .I1(n17_adj_4721), .CO(n28174));
    SB_LUT4 displacement_23__I_0_add_2_9_lut (.I0(GND_net), .I1(displacement_23__N_229[7]), 
            .I2(n18_adj_4722), .I3(n28172), .O(displacement_23__N_80[7])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_9 (.CI(n28172), .I0(displacement_23__N_229[7]), 
            .I1(n18_adj_4722), .CO(n28173));
    SB_CARRY rem_4_add_1050_9 (.CI(n29059), .I0(n1551), .I1(VCC_net), 
            .CO(n29060));
    SB_LUT4 rem_4_add_1050_8_lut (.I0(GND_net), .I1(n1552), .I2(VCC_net), 
            .I3(n29058), .O(n1619)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_5_lut (.I0(GND_net), .I1(n2656), .I2(VCC_net), 
            .I3(n28849), .O(n2723_adj_4824)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 displacement_23__I_0_add_2_8_lut (.I0(GND_net), .I1(displacement_23__N_229[6]), 
            .I2(n19_adj_4723), .I3(n28171), .O(displacement_23__N_80[6])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_8 (.CI(n28171), .I0(displacement_23__N_229[6]), 
            .I1(n19_adj_4723), .CO(n28172));
    SB_LUT4 displacement_23__I_0_add_2_7_lut (.I0(GND_net), .I1(displacement_23__N_229[5]), 
            .I2(n20_adj_4724), .I3(n28170), .O(displacement_23__N_80[5])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_7 (.CI(n28170), .I0(displacement_23__N_229[5]), 
            .I1(n20_adj_4724), .CO(n28171));
    SB_LUT4 displacement_23__I_0_add_2_6_lut (.I0(GND_net), .I1(displacement_23__N_229[4]), 
            .I2(n21_adj_4725), .I3(n28169), .O(displacement_23__N_80[4])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_8 (.CI(n29058), .I0(n1552), .I1(VCC_net), 
            .CO(n29059));
    SB_CARRY rem_4_add_1787_5 (.CI(n28849), .I0(n2656), .I1(VCC_net), 
            .CO(n28850));
    SB_LUT4 rem_4_add_1787_4_lut (.I0(GND_net), .I1(n2657), .I2(VCC_net), 
            .I3(n28848), .O(n2724_adj_4823)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_6 (.CI(n28169), .I0(displacement_23__N_229[4]), 
            .I1(n21_adj_4725), .CO(n28170));
    SB_LUT4 displacement_23__I_0_add_2_5_lut (.I0(GND_net), .I1(displacement_23__N_229[3]), 
            .I2(n22_adj_4726), .I3(n28168), .O(displacement_23__N_80[3])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY displacement_23__I_0_add_2_5 (.CI(n28168), .I0(displacement_23__N_229[3]), 
            .I1(n22_adj_4726), .CO(n28169));
    SB_LUT4 displacement_23__I_0_add_2_4_lut (.I0(GND_net), .I1(displacement_23__N_229[2]), 
            .I2(n23_adj_4727), .I3(n28167), .O(displacement_23__N_80[2])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_4 (.CI(n28848), .I0(n2657), .I1(VCC_net), 
            .CO(n28849));
    SB_CARRY displacement_23__I_0_add_2_4 (.CI(n28167), .I0(displacement_23__N_229[2]), 
            .I1(n23_adj_4727), .CO(n28168));
    SB_LUT4 displacement_23__I_0_add_2_3_lut (.I0(GND_net), .I1(displacement_23__N_229[1]), 
            .I2(n24_adj_4728), .I3(n28166), .O(displacement_23__N_80[1])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1787_3_lut (.I0(GND_net), .I1(n2658), .I2(GND_net), 
            .I3(n28847), .O(n2725)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1787_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_3 (.CI(n28847), .I0(n2658), .I1(GND_net), 
            .CO(n28848));
    SB_CARRY displacement_23__I_0_add_2_3 (.CI(n28166), .I0(displacement_23__N_229[1]), 
            .I1(n24_adj_4728), .CO(n28167));
    SB_LUT4 displacement_23__I_0_add_2_2_lut (.I0(GND_net), .I1(displacement_23__N_229[0]), 
            .I2(n25_adj_4729), .I3(VCC_net), .O(displacement_23__N_80[0])) /* synthesis syn_instantiated=1 */ ;
    defparam displacement_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1787_2 (.CI(VCC_net), .I0(n2758), .I1(VCC_net), 
            .CO(n28847));
    SB_CARRY displacement_23__I_0_add_2_2 (.CI(VCC_net), .I0(displacement_23__N_229[0]), 
            .I1(n25_adj_4729), .CO(n28166));
    SB_LUT4 rem_4_add_1050_7_lut (.I0(GND_net), .I1(n1553), .I2(VCC_net), 
            .I3(n29057), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_7 (.CI(n29057), .I0(n1553), .I1(VCC_net), 
            .CO(n29058));
    SB_LUT4 rem_4_add_1854_26_lut (.I0(n2768), .I1(n2735), .I2(VCC_net), 
            .I3(n28846), .O(n2834)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1854_25_lut (.I0(GND_net), .I1(n2736), .I2(VCC_net), 
            .I3(n28845), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_6_lut (.I0(GND_net), .I1(n1554), .I2(GND_net), 
            .I3(n29056), .O(n1621)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_25 (.CI(n28845), .I0(n2736), .I1(VCC_net), 
            .CO(n28846));
    SB_LUT4 rem_4_add_1854_24_lut (.I0(GND_net), .I1(n2737), .I2(VCC_net), 
            .I3(n28844), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_24 (.CI(n28844), .I0(n2737), .I1(VCC_net), 
            .CO(n28845));
    SB_LUT4 rem_4_add_1854_23_lut (.I0(GND_net), .I1(n2738), .I2(VCC_net), 
            .I3(n28843), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_6 (.CI(n29056), .I0(n1554), .I1(GND_net), 
            .CO(n29057));
    SB_CARRY rem_4_add_1854_23 (.CI(n28843), .I0(n2738), .I1(VCC_net), 
            .CO(n28844));
    SB_LUT4 rem_4_add_1050_5_lut (.I0(GND_net), .I1(n1555), .I2(GND_net), 
            .I3(n29055), .O(n1622)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i723_3_lut_3_lut (.I0(n1067), .I1(n5957), .I2(n1047), 
            .I3(GND_net), .O(n1173));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i723_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_1050_5 (.CI(n29055), .I0(n1555), .I1(GND_net), 
            .CO(n29056));
    SB_LUT4 rem_4_add_1854_22_lut (.I0(GND_net), .I1(n2739), .I2(VCC_net), 
            .I3(n28842), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_4_lut (.I0(GND_net), .I1(n1556), .I2(VCC_net), 
            .I3(n29054), .O(n1623)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_22 (.CI(n28842), .I0(n2739), .I1(VCC_net), 
            .CO(n28843));
    SB_LUT4 rem_4_add_1854_21_lut (.I0(GND_net), .I1(n2740), .I2(VCC_net), 
            .I3(n28841), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i724_3_lut_3_lut (.I0(n1067), .I1(n5958), .I2(n1048), 
            .I3(GND_net), .O(n1174));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i724_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i725_3_lut_3_lut (.I0(n1067), .I1(n5959), .I2(n1049), 
            .I3(GND_net), .O(n1175));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i725_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i722_3_lut_3_lut (.I0(n1067), .I1(n5956), .I2(n1046), 
            .I3(GND_net), .O(n1172));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i722_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i721_3_lut_3_lut (.I0(n1067), .I1(n5955), .I2(n1045), 
            .I3(GND_net), .O(n1171));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i721_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i719_3_lut_3_lut (.I0(n1067), .I1(n5953), .I2(n1043), 
            .I3(GND_net), .O(n1169));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i720_3_lut_3_lut (.I0(n1067), .I1(n5954), .I2(n1044), 
            .I3(GND_net), .O(n1170_adj_4738));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i720_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_983_12_lut (.I0(n1481), .I1(n1448), .I2(VCC_net), 
            .I3(n28142), .O(n1547)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_983_11_lut (.I0(GND_net), .I1(n1449), .I2(VCC_net), 
            .I3(n28141), .O(n1516)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14_4_lut_adj_1804 (.I0(n2249), .I1(n28_adj_5244), .I2(n24_adj_5246), 
            .I3(n16_adj_5248), .O(n2273_adj_4953));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i14_4_lut_adj_1804.LUT_INIT = 16'hfffe;
    SB_CARRY rem_4_add_983_11 (.CI(n28141), .I0(n1449), .I1(VCC_net), 
            .CO(n28142));
    SB_LUT4 div_46_LessThan_657_i40_3_lut_3_lut (.I0(n1046), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n40_adj_4936));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_657_i40_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_CARRY rem_4_add_1050_4 (.CI(n29054), .I0(n1556), .I1(VCC_net), 
            .CO(n29055));
    SB_CARRY rem_4_add_1854_21 (.CI(n28841), .I0(n2740), .I1(VCC_net), 
            .CO(n28842));
    SB_LUT4 rem_4_add_983_10_lut (.I0(GND_net), .I1(n1450), .I2(VCC_net), 
            .I3(n28140), .O(n1517)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_20_lut (.I0(GND_net), .I1(n2741), .I2(VCC_net), 
            .I3(n28840), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_3_lut (.I0(GND_net), .I1(n1557), .I2(VCC_net), 
            .I3(n29053), .O(n1624)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1050_3 (.CI(n29053), .I0(n1557), .I1(VCC_net), 
            .CO(n29054));
    SB_CARRY rem_4_add_1854_20 (.CI(n28840), .I0(n2741), .I1(VCC_net), 
            .CO(n28841));
    SB_CARRY rem_4_add_983_10 (.CI(n28140), .I0(n1450), .I1(VCC_net), 
            .CO(n28141));
    SB_LUT4 rem_4_add_983_9_lut (.I0(GND_net), .I1(n1451), .I2(VCC_net), 
            .I3(n28139), .O(n1518)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_9 (.CI(n28139), .I0(n1451), .I1(VCC_net), .CO(n28140));
    SB_LUT4 rem_4_add_983_8_lut (.I0(GND_net), .I1(n1452), .I2(VCC_net), 
            .I3(n28138), .O(n1519)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_8 (.CI(n28138), .I0(n1452), .I1(VCC_net), .CO(n28139));
    SB_LUT4 rem_4_add_983_7_lut (.I0(GND_net), .I1(n1453), .I2(VCC_net), 
            .I3(n28137), .O(n1520)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_7 (.CI(n28137), .I0(n1453), .I1(VCC_net), .CO(n28138));
    SB_LUT4 rem_4_add_983_6_lut (.I0(GND_net), .I1(n1454), .I2(GND_net), 
            .I3(n28136), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_6 (.CI(n28136), .I0(n1454), .I1(GND_net), .CO(n28137));
    SB_LUT4 rem_4_add_983_5_lut (.I0(GND_net), .I1(n1455), .I2(GND_net), 
            .I3(n28135), .O(n1522)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_5 (.CI(n28135), .I0(n1455), .I1(GND_net), .CO(n28136));
    SB_LUT4 rem_4_add_983_4_lut (.I0(GND_net), .I1(n1456), .I2(VCC_net), 
            .I3(n28134), .O(n1523)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1050_2_lut (.I0(GND_net), .I1(n1558), .I2(GND_net), 
            .I3(VCC_net), .O(n1625)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1050_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_19_lut (.I0(GND_net), .I1(n2742), .I2(VCC_net), 
            .I3(n28839), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_4 (.CI(n28134), .I0(n1456), .I1(VCC_net), .CO(n28135));
    SB_CARRY rem_4_add_1854_19 (.CI(n28839), .I0(n2742), .I1(VCC_net), 
            .CO(n28840));
    SB_CARRY rem_4_add_1050_2 (.CI(VCC_net), .I0(n1558), .I1(GND_net), 
            .CO(n29053));
    SB_LUT4 rem_4_add_1854_18_lut (.I0(GND_net), .I1(n2743), .I2(VCC_net), 
            .I3(n28838), .O(n2810)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_983_3_lut (.I0(GND_net), .I1(n1457), .I2(VCC_net), 
            .I3(n28133), .O(n1524)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_983_3 (.CI(n28133), .I0(n1457), .I1(VCC_net), .CO(n28134));
    SB_LUT4 rem_4_add_983_2_lut (.I0(GND_net), .I1(n1458), .I2(GND_net), 
            .I3(VCC_net), .O(n1525)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_983_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1117_15_lut (.I0(n1679), .I1(n1646_adj_4813), .I2(VCC_net), 
            .I3(n29052), .O(n1745)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY rem_4_add_1854_18 (.CI(n28838), .I0(n2743), .I1(VCC_net), 
            .CO(n28839));
    SB_CARRY rem_4_add_983_2 (.CI(VCC_net), .I0(n1458), .I1(GND_net), 
            .CO(n28133));
    SB_LUT4 rem_4_add_1117_14_lut (.I0(GND_net), .I1(n1647_adj_4814), .I2(VCC_net), 
            .I3(n29051), .O(n1714)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_17_lut (.I0(GND_net), .I1(n2744), .I2(VCC_net), 
            .I3(n28837), .O(n2811)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_14 (.CI(n29051), .I0(n1647_adj_4814), .I1(VCC_net), 
            .CO(n29052));
    SB_CARRY rem_4_add_1854_17 (.CI(n28837), .I0(n2744), .I1(VCC_net), 
            .CO(n28838));
    SB_LUT4 rem_4_add_1117_13_lut (.I0(GND_net), .I1(n1648_adj_4815), .I2(VCC_net), 
            .I3(n29050), .O(n1715)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_16_lut (.I0(GND_net), .I1(n2745), .I2(VCC_net), 
            .I3(n28836), .O(n2812)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_13 (.CI(n29050), .I0(n1648_adj_4815), .I1(VCC_net), 
            .CO(n29051));
    SB_CARRY rem_4_add_1854_16 (.CI(n28836), .I0(n2745), .I1(VCC_net), 
            .CO(n28837));
    SB_LUT4 rem_4_add_1117_12_lut (.I0(GND_net), .I1(n1649_adj_4816), .I2(VCC_net), 
            .I3(n29049), .O(n1716)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_15_lut (.I0(GND_net), .I1(n2746), .I2(VCC_net), 
            .I3(n28835), .O(n2813)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_15 (.CI(n28835), .I0(n2746), .I1(VCC_net), 
            .CO(n28836));
    SB_CARRY rem_4_add_1117_12 (.CI(n29049), .I0(n1649_adj_4816), .I1(VCC_net), 
            .CO(n29050));
    SB_LUT4 rem_4_add_1854_14_lut (.I0(GND_net), .I1(n2747), .I2(VCC_net), 
            .I3(n28834), .O(n2814)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_562_24_lut (.I0(duty[22]), .I1(n43653), .I2(n3), .I3(n28122), 
            .O(pwm_setpoint_22__N_57[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_562_23_lut (.I0(duty[21]), .I1(n43653), .I2(n4_adj_4658), 
            .I3(n28121), .O(pwm_setpoint_22__N_57[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_562_23 (.CI(n28121), .I0(n43653), .I1(n4_adj_4658), .CO(n28122));
    SB_LUT4 add_562_22_lut (.I0(duty[20]), .I1(n43653), .I2(n5), .I3(n28120), 
            .O(pwm_setpoint_22__N_57[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1854_14 (.CI(n28834), .I0(n2747), .I1(VCC_net), 
            .CO(n28835));
    SB_LUT4 rem_4_add_1117_11_lut (.I0(GND_net), .I1(n1650_adj_4817), .I2(VCC_net), 
            .I3(n29048), .O(n1717)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_13_lut (.I0(GND_net), .I1(n2748), .I2(VCC_net), 
            .I3(n28833), .O(n2815)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_562_22 (.CI(n28120), .I0(n43653), .I1(n5), .CO(n28121));
    SB_CARRY rem_4_add_1854_13 (.CI(n28833), .I0(n2748), .I1(VCC_net), 
            .CO(n28834));
    SB_LUT4 add_562_21_lut (.I0(duty[19]), .I1(n43653), .I2(n6), .I3(n28119), 
            .O(pwm_setpoint_22__N_57[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_562_21 (.CI(n28119), .I0(n43653), .I1(n6), .CO(n28120));
    SB_LUT4 add_562_20_lut (.I0(duty[18]), .I1(n43653), .I2(n7), .I3(n28118), 
            .O(pwm_setpoint_22__N_57[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_562_20 (.CI(n28118), .I0(n43653), .I1(n7), .CO(n28119));
    SB_LUT4 add_562_19_lut (.I0(duty[17]), .I1(n43653), .I2(n8), .I3(n28117), 
            .O(pwm_setpoint_22__N_57[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_562_19 (.CI(n28117), .I0(n43653), .I1(n8), .CO(n28118));
    SB_LUT4 add_562_18_lut (.I0(duty[16]), .I1(n43653), .I2(n9), .I3(n28116), 
            .O(pwm_setpoint_22__N_57[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_562_18 (.CI(n28116), .I0(n43653), .I1(n9), .CO(n28117));
    SB_CARRY rem_4_add_1117_11 (.CI(n29048), .I0(n1650_adj_4817), .I1(VCC_net), 
            .CO(n29049));
    SB_LUT4 rem_4_add_1854_12_lut (.I0(GND_net), .I1(n2749), .I2(VCC_net), 
            .I3(n28832), .O(n2816)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_562_17_lut (.I0(duty[15]), .I1(n43653), .I2(n10_adj_4659), 
            .I3(n28115), .O(pwm_setpoint_22__N_57[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_562_17 (.CI(n28115), .I0(n43653), .I1(n10_adj_4659), 
            .CO(n28116));
    SB_LUT4 add_562_16_lut (.I0(duty[14]), .I1(n43653), .I2(n11), .I3(n28114), 
            .O(pwm_setpoint_22__N_57[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_16_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_562_16 (.CI(n28114), .I0(n43653), .I1(n11), .CO(n28115));
    SB_LUT4 add_562_15_lut (.I0(duty[13]), .I1(n43653), .I2(n12), .I3(n28113), 
            .O(pwm_setpoint_22__N_57[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_15_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_562_15 (.CI(n28113), .I0(n43653), .I1(n12), .CO(n28114));
    SB_LUT4 rem_4_add_1117_10_lut (.I0(GND_net), .I1(n1651_adj_4818), .I2(VCC_net), 
            .I3(n29047), .O(n1718)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34053_3_lut_4_lut (.I0(n1046), .I1(n97), .I2(n98), .I3(n1047), 
            .O(n40899));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34053_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 add_562_14_lut (.I0(duty[12]), .I1(n43653), .I2(n13), .I3(n28112), 
            .O(pwm_setpoint_22__N_57[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1854_12 (.CI(n28832), .I0(n2749), .I1(VCC_net), 
            .CO(n28833));
    SB_CARRY add_562_14 (.CI(n28112), .I0(n43653), .I1(n13), .CO(n28113));
    SB_LUT4 add_562_13_lut (.I0(duty[11]), .I1(n43653), .I2(n14), .I3(n28111), 
            .O(pwm_setpoint_22__N_57[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_562_13 (.CI(n28111), .I0(n43653), .I1(n14), .CO(n28112));
    SB_LUT4 add_562_12_lut (.I0(duty[10]), .I1(n43653), .I2(n15_adj_4660), 
            .I3(n28110), .O(pwm_setpoint_22__N_57[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_562_12 (.CI(n28110), .I0(n43653), .I1(n15_adj_4660), 
            .CO(n28111));
    SB_LUT4 add_562_11_lut (.I0(duty[9]), .I1(n43653), .I2(n16_adj_4661), 
            .I3(n28109), .O(pwm_setpoint_22__N_57[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_562_11 (.CI(n28109), .I0(n43653), .I1(n16_adj_4661), 
            .CO(n28110));
    SB_LUT4 add_562_10_lut (.I0(duty[8]), .I1(n43653), .I2(n17), .I3(n28108), 
            .O(pwm_setpoint_22__N_57[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY rem_4_add_1117_10 (.CI(n29047), .I0(n1651_adj_4818), .I1(VCC_net), 
            .CO(n29048));
    SB_CARRY add_562_10 (.CI(n28108), .I0(n43653), .I1(n17), .CO(n28109));
    SB_LUT4 add_562_9_lut (.I0(duty[7]), .I1(n43653), .I2(n18_adj_4662), 
            .I3(n28107), .O(pwm_setpoint_22__N_57[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 div_46_LessThan_1062_i39_2_lut (.I0(n1647), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4980));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1062_i39_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY add_562_9 (.CI(n28107), .I0(n43653), .I1(n18_adj_4662), .CO(n28108));
    SB_LUT4 add_562_8_lut (.I0(duty[6]), .I1(n43653), .I2(n19), .I3(n28106), 
            .O(pwm_setpoint_22__N_57[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1854_11_lut (.I0(GND_net), .I1(n2750), .I2(VCC_net), 
            .I3(n28831), .O(n2817)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_562_8 (.CI(n28106), .I0(n43653), .I1(n19), .CO(n28107));
    SB_LUT4 add_562_7_lut (.I0(duty[5]), .I1(n43653), .I2(n20_adj_4663), 
            .I3(n28105), .O(pwm_setpoint_22__N_57[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_562_7 (.CI(n28105), .I0(n43653), .I1(n20_adj_4663), .CO(n28106));
    SB_LUT4 add_562_6_lut (.I0(duty[4]), .I1(n43653), .I2(n21), .I3(n28104), 
            .O(pwm_setpoint_22__N_57[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 rem_4_add_1117_9_lut (.I0(GND_net), .I1(n1652_adj_4819), .I2(VCC_net), 
            .I3(n29046), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_562_6 (.CI(n28104), .I0(n43653), .I1(n21), .CO(n28105));
    SB_CARRY rem_4_add_1854_11 (.CI(n28831), .I0(n2750), .I1(VCC_net), 
            .CO(n28832));
    SB_LUT4 add_562_5_lut (.I0(duty[3]), .I1(n43653), .I2(n22), .I3(n28103), 
            .O(pwm_setpoint_22__N_57[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_562_5 (.CI(n28103), .I0(n43653), .I1(n22), .CO(n28104));
    SB_LUT4 add_562_4_lut (.I0(duty[2]), .I1(n43653), .I2(n23), .I3(n28102), 
            .O(pwm_setpoint_22__N_57[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_562_4 (.CI(n28102), .I0(n43653), .I1(n23), .CO(n28103));
    SB_LUT4 add_562_3_lut (.I0(duty[1]), .I1(n43653), .I2(n24), .I3(n28101), 
            .O(pwm_setpoint_22__N_57[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_562_3 (.CI(n28101), .I0(n43653), .I1(n24), .CO(n28102));
    SB_LUT4 add_562_2_lut (.I0(duty[0]), .I1(n43653), .I2(n25), .I3(VCC_net), 
            .O(pwm_setpoint_22__N_57[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_562_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_562_2 (.CI(VCC_net), .I0(n43653), .I1(n25), .CO(n28101));
    SB_CARRY rem_4_add_1117_9 (.CI(n29046), .I0(n1652_adj_4819), .I1(VCC_net), 
            .CO(n29047));
    SB_LUT4 rem_4_add_1854_10_lut (.I0(GND_net), .I1(n2751), .I2(VCC_net), 
            .I3(n28830), .O(n2818)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1117_8_lut (.I0(GND_net), .I1(n1653_adj_4820), .I2(VCC_net), 
            .I3(n29045), .O(n1720)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_8 (.CI(n29045), .I0(n1653_adj_4820), .I1(VCC_net), 
            .CO(n29046));
    SB_CARRY rem_4_add_1854_10 (.CI(n28830), .I0(n2751), .I1(VCC_net), 
            .CO(n28831));
    SB_LUT4 div_46_i808_3_lut_3_lut (.I0(n1193), .I1(n5968), .I2(n1175), 
            .I3(GND_net), .O(n1298));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i808_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1117_7_lut (.I0(GND_net), .I1(n1654), .I2(GND_net), 
            .I3(n29044), .O(n1721)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_9_lut (.I0(GND_net), .I1(n2752), .I2(VCC_net), 
            .I3(n28829), .O(n2819)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_7 (.CI(n29044), .I0(n1654), .I1(GND_net), 
            .CO(n29045));
    SB_CARRY rem_4_add_1854_9 (.CI(n28829), .I0(n2752), .I1(VCC_net), 
            .CO(n28830));
    SB_LUT4 div_46_i809_3_lut_3_lut (.I0(n1193), .I1(n5969), .I2(n1050), 
            .I3(GND_net), .O(n1299));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i809_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1117_6_lut (.I0(GND_net), .I1(n1655), .I2(GND_net), 
            .I3(n29043), .O(n1722)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_6 (.CI(n29043), .I0(n1655), .I1(GND_net), 
            .CO(n29044));
    SB_LUT4 rem_4_add_1854_8_lut (.I0(GND_net), .I1(n2753), .I2(VCC_net), 
            .I3(n28828), .O(n2820)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_8 (.CI(n28828), .I0(n2753), .I1(VCC_net), 
            .CO(n28829));
    SB_LUT4 div_46_i805_3_lut_3_lut (.I0(n1193), .I1(n5965), .I2(n1172), 
            .I3(GND_net), .O(n1295));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i805_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i804_3_lut_3_lut (.I0(n1193), .I1(n5964), .I2(n1171), 
            .I3(GND_net), .O(n1294));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i804_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_1117_5_lut (.I0(GND_net), .I1(n1656), .I2(VCC_net), 
            .I3(n29042), .O(n1723)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_7_lut (.I0(GND_net), .I1(n2754), .I2(GND_net), 
            .I3(n28827), .O(n2821)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_i1467_3_lut (.I0(n2154), .I1(n2221), .I2(n2174_adj_4984), 
            .I3(GND_net), .O(n2253));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1467_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY rem_4_add_1117_5 (.CI(n29042), .I0(n1656), .I1(VCC_net), 
            .CO(n29043));
    SB_CARRY rem_4_add_1854_7 (.CI(n28827), .I0(n2754), .I1(GND_net), 
            .CO(n28828));
    SB_LUT4 rem_4_add_1854_6_lut (.I0(GND_net), .I1(n2755), .I2(GND_net), 
            .I3(n28826), .O(n2822)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1117_4_lut (.I0(GND_net), .I1(n1657), .I2(VCC_net), 
            .I3(n29041), .O(n1724)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_LessThan_1062_i37_2_lut (.I0(n1648), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4979));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1062_i37_2_lut.LUT_INIT = 16'h9999;
    SB_CARRY rem_4_add_1117_4 (.CI(n29041), .I0(n1657), .I1(VCC_net), 
            .CO(n29042));
    SB_CARRY rem_4_add_1854_6 (.CI(n28826), .I0(n2755), .I1(GND_net), 
            .CO(n28827));
    SB_LUT4 rem_4_add_1117_3_lut (.I0(GND_net), .I1(n1658), .I2(GND_net), 
            .I3(n29040), .O(n1725)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1117_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_1854_5_lut (.I0(GND_net), .I1(n2756), .I2(VCC_net), 
            .I3(n28825), .O(n2823)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1117_3 (.CI(n29040), .I0(n1658), .I1(GND_net), 
            .CO(n29041));
    SB_CARRY rem_4_add_1854_5 (.CI(n28825), .I0(n2756), .I1(VCC_net), 
            .CO(n28826));
    SB_LUT4 rem_4_add_1854_4_lut (.I0(GND_net), .I1(n2757), .I2(VCC_net), 
            .I3(n28824), .O(n2824)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF blink_53 (.Q(blink), .C(LED_c), .D(blink_N_255));   // verilog/TinyFPGA_B.v(51[8] 74[4])
    SB_CARRY rem_4_add_1117_2 (.CI(VCC_net), .I0(n1758_adj_4811), .I1(VCC_net), 
            .CO(n29040));
    SB_CARRY rem_4_add_1854_4 (.CI(n28824), .I0(n2757), .I1(VCC_net), 
            .CO(n28825));
    SB_LUT4 div_46_i806_3_lut_3_lut (.I0(n1193), .I1(n5966), .I2(n1173), 
            .I3(GND_net), .O(n1296));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i806_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_849_10_lut (.I0(n1283), .I1(n1250), .I2(VCC_net), 
            .I3(n29039), .O(n1349)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_1854_3_lut (.I0(GND_net), .I1(n2758), .I2(GND_net), 
            .I3(n28823), .O(n2825)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_1854_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_849_9_lut (.I0(GND_net), .I1(n1251), .I2(VCC_net), 
            .I3(n29038), .O(n1318)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_1854_3 (.CI(n28823), .I0(n2758), .I1(GND_net), 
            .CO(n28824));
    SB_CARRY rem_4_add_849_9 (.CI(n29038), .I0(n1251), .I1(VCC_net), .CO(n29039));
    SB_CARRY rem_4_add_1854_2 (.CI(VCC_net), .I0(n2858), .I1(VCC_net), 
            .CO(n28823));
    SB_LUT4 div_46_unary_minus_2_add_3_25_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(n2_adj_4912), .I3(n28822), .O(n224)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 rem_4_add_849_8_lut (.I0(GND_net), .I1(n1252), .I2(VCC_net), 
            .I3(n29037), .O(n1319)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_8 (.CI(n29037), .I0(n1252), .I1(VCC_net), .CO(n29038));
    SB_LUT4 div_46_unary_minus_2_add_3_24_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n3_adj_4913), .I3(n28821), .O(n3_adj_4694)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i803_3_lut_3_lut (.I0(n1193), .I1(n5963), .I2(n1170_adj_4738), 
            .I3(GND_net), .O(n1293));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i803_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_add_849_7_lut (.I0(GND_net), .I1(n1253), .I2(VCC_net), 
            .I3(n29036), .O(n1320)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_24 (.CI(n28821), .I0(GND_net), .I1(n3_adj_4913), 
            .CO(n28822));
    SB_CARRY rem_4_add_849_7 (.CI(n29036), .I0(n1253), .I1(VCC_net), .CO(n29037));
    SB_LUT4 div_46_unary_minus_2_add_3_23_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n4_adj_4914), .I3(n28820), .O(n4_adj_4693)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 rem_4_add_849_6_lut (.I0(GND_net), .I1(n1254), .I2(GND_net), 
            .I3(n29035), .O(n1321)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_23 (.CI(n28820), .I0(GND_net), .I1(n4_adj_4914), 
            .CO(n28821));
    SB_CARRY rem_4_add_849_6 (.CI(n29035), .I0(n1254), .I1(GND_net), .CO(n29036));
    SB_LUT4 rem_4_add_849_5_lut (.I0(GND_net), .I1(n1255), .I2(GND_net), 
            .I3(n29034), .O(n1322)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_unary_minus_2_add_3_22_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n5_adj_4915), .I3(n28819), .O(n5_adj_4692)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY rem_4_add_849_5 (.CI(n29034), .I0(n1255), .I1(GND_net), .CO(n29035));
    SB_CARRY div_46_unary_minus_2_add_3_22 (.CI(n28819), .I0(GND_net), .I1(n5_adj_4915), 
            .CO(n28820));
    SB_LUT4 rem_4_add_849_4_lut (.I0(GND_net), .I1(n1256), .I2(VCC_net), 
            .I3(n29033), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i802_3_lut_3_lut (.I0(n1193), .I1(n5962), .I2(n1169), 
            .I3(GND_net), .O(n1292));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i802_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_CARRY rem_4_add_849_4 (.CI(n29033), .I0(n1256), .I1(VCC_net), .CO(n29034));
    SB_LUT4 div_46_unary_minus_2_add_3_21_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n6_adj_4916), .I3(n28818), .O(n6_adj_4706)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_21 (.CI(n28818), .I0(GND_net), .I1(n6_adj_4916), 
            .CO(n28819));
    SB_LUT4 rem_4_add_849_3_lut (.I0(GND_net), .I1(n1257), .I2(VCC_net), 
            .I3(n29032), .O(n1324)) /* synthesis syn_instantiated=1 */ ;
    defparam rem_4_add_849_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 div_46_i807_3_lut_3_lut (.I0(n1193), .I1(n5967), .I2(n1174), 
            .I3(GND_net), .O(n1297));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i807_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_mux_3_i13_3_lut (.I0(encoder0_position[12]), .I1(n13_adj_4697), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n1054_adj_4733));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_unary_minus_2_add_3_20_lut (.I0(GND_net), .I1(GND_net), 
            .I2(n7_adj_4917), .I3(n28817), .O(n7_adj_4705)) /* synthesis syn_instantiated=1 */ ;
    defparam div_46_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY div_46_unary_minus_2_add_3_20 (.CI(n28817), .I0(GND_net), .I1(n7_adj_4917), 
            .CO(n28818));
    SB_LUT4 div_46_LessThan_1062_i43_2_lut (.I0(n1645), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4983));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1062_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i35318_3_lut (.I0(n2152), .I1(n2219), .I2(n2174_adj_4984), 
            .I3(GND_net), .O(n2251));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i35318_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_742_i38_3_lut_3_lut (.I0(n1173), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n38_adj_4943));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_742_i38_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_4_lut_adj_1805 (.I0(n5_adj_4766), .I1(n122), .I2(n2774), 
            .I3(n63_adj_4745), .O(n6_adj_5357));   // verilog/coms.v(127[12] 295[6])
    defparam i1_4_lut_adj_1805.LUT_INIT = 16'heaaa;
    SB_LUT4 i34043_3_lut_4_lut (.I0(n1173), .I1(n97), .I2(n98), .I3(n1174), 
            .O(n40889));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34043_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1062_i31_2_lut (.I0(n1651), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4975));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1062_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1062_i33_2_lut (.I0(n1650), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4977));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1062_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1062_i35_2_lut (.I0(n1649), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4978));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1062_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_1062_i41_2_lut (.I0(n1646), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4982));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1062_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i1064_1_lut (.I0(n1667), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1668));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1064_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_1062_i29_2_lut (.I0(n1652), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_4973));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1062_i29_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33959_4_lut (.I0(n35_adj_4978), .I1(n33_adj_4977), .I2(n31_adj_4975), 
            .I3(n29_adj_4973), .O(n40805));
    defparam i33959_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 div_46_LessThan_1062_i40_3_lut (.I0(n32_adj_4976), .I1(n91), 
            .I2(n43_adj_4983), .I3(GND_net), .O(n40_adj_4981));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1062_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_1062_i28_4_lut (.I0(n1054_adj_4733), .I1(n99), 
            .I2(n1653), .I3(n558), .O(n28_adj_4972));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1062_i28_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35750_3_lut (.I0(n28_adj_4972), .I1(n95), .I2(n35_adj_4978), 
            .I3(GND_net), .O(n42597));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35750_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35751_3_lut (.I0(n42597), .I1(n94), .I2(n37_adj_4979), .I3(GND_net), 
            .O(n42598));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35751_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33952_4_lut (.I0(n41_adj_4982), .I1(n39_adj_4980), .I2(n37_adj_4979), 
            .I3(n40805), .O(n40798));
    defparam i33952_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35748_4_lut (.I0(n40_adj_4981), .I1(n30_adj_4974), .I2(n43_adj_4983), 
            .I3(n40794), .O(n42595));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35748_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35561_3_lut (.I0(n42598), .I1(n93), .I2(n39_adj_4980), .I3(GND_net), 
            .O(n42408));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35561_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35932_4_lut (.I0(n42408), .I1(n42595), .I2(n43_adj_4983), 
            .I3(n40798), .O(n42779));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35932_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35933_3_lut (.I0(n42779), .I1(n90), .I2(n1644), .I3(GND_net), 
            .O(n42780));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35933_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1806 (.I0(n42780), .I1(n15889), .I2(n89), .I3(n1643), 
            .O(n1667));
    defparam i1_4_lut_adj_1806.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_985_i39_2_lut (.I0(n1533), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4967));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_985_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_985_i41_2_lut (.I0(n1532), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4968));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_985_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i14_3_lut (.I0(encoder0_position[13]), .I1(n12_adj_4698), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n1053_adj_4732));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1807 (.I0(n44342), .I1(n6_adj_5357), .I2(n15994), 
            .I3(n3894), .O(n8_adj_5243));   // verilog/coms.v(127[12] 295[6])
    defparam i3_4_lut_adj_1807.LUT_INIT = 16'hcfce;
    SB_LUT4 div_46_LessThan_985_i45_2_lut (.I0(n1530), .I1(n91), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4971));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_985_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_985_i33_2_lut (.I0(n1536), .I1(n97), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_4963));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_985_i33_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_985_i35_2_lut (.I0(n1535), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4965));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_985_i35_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_985_i37_2_lut (.I0(n1534), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_4966));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_985_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_985_i43_2_lut (.I0(n1531), .I1(n92), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4970));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_985_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i987_1_lut (.I0(n1553_adj_4742), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1554_adj_4743));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i987_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_985_i31_2_lut (.I0(n1537), .I1(n98), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_4961));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_985_i31_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i33982_4_lut (.I0(n37_adj_4966), .I1(n35_adj_4965), .I2(n33_adj_4963), 
            .I3(n31_adj_4961), .O(n40828));
    defparam i33982_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 rem_4_i1535_rep_57_3_lut (.I0(n2254), .I1(n2321), .I2(n2273_adj_4953), 
            .I3(GND_net), .O(n2353));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1535_rep_57_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_985_i42_3_lut (.I0(n34_adj_4964), .I1(n91), 
            .I2(n45_adj_4971), .I3(GND_net), .O(n42_adj_4969));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_985_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_LessThan_985_i30_4_lut (.I0(n1053_adj_4732), .I1(n99), 
            .I2(n1538), .I3(n558), .O(n30_adj_4960));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_985_i30_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35754_3_lut (.I0(n30_adj_4960), .I1(n95), .I2(n37_adj_4966), 
            .I3(GND_net), .O(n42601));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35754_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i4_4_lut_adj_1808 (.I0(n122), .I1(n8_adj_5243), .I2(n63_adj_4657), 
            .I3(n5_adj_5338), .O(n43830));   // verilog/coms.v(127[12] 295[6])
    defparam i4_4_lut_adj_1808.LUT_INIT = 16'hefcf;
    SB_LUT4 i35755_3_lut (.I0(n42601), .I1(n94), .I2(n39_adj_4967), .I3(GND_net), 
            .O(n42602));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35755_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i33974_4_lut (.I0(n43_adj_4970), .I1(n41_adj_4968), .I2(n39_adj_4967), 
            .I3(n40828), .O(n40820));
    defparam i33974_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35310_4_lut (.I0(n42_adj_4969), .I1(n32_adj_4962), .I2(n45_adj_4971), 
            .I3(n40818), .O(n42157));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35310_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 rem_4_mux_3_i13_3_lut (.I0(communication_counter[12]), .I1(n21_adj_4788), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2358_adj_4940));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35557_3_lut (.I0(n42602), .I1(n93), .I2(n41_adj_4968), .I3(GND_net), 
            .O(n42404));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35557_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 rem_4_i1538_3_lut (.I0(n2257), .I1(n2324), .I2(n2273_adj_4953), 
            .I3(GND_net), .O(n2356));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35776_4_lut (.I0(n42404), .I1(n42157), .I2(n45_adj_4971), 
            .I3(n40820), .O(n42623));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35776_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_4_lut_adj_1809 (.I0(n42623), .I1(n15974), .I2(n90), .I3(n1529), 
            .O(n1553_adj_4742));
    defparam i1_4_lut_adj_1809.LUT_INIT = 16'hceef;
    SB_LUT4 i13161_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n13302), 
            .I3(GND_net), .O(n17900));   // verilog/coms.v(127[12] 295[6])
    defparam i13161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13162_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n13302), 
            .I3(GND_net), .O(n17901));   // verilog/coms.v(127[12] 295[6])
    defparam i13162_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_LessThan_906_i43_2_lut (.I0(n1414), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4959));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_906_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_906_i41_2_lut (.I0(n1415), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4958));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_906_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_906_i37_2_lut (.I0(n1417_adj_4739), .I1(n96), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4956));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_906_i37_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_906_i39_2_lut (.I0(n1416), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4957));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_906_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i15_3_lut (.I0(encoder0_position[14]), .I1(n11_adj_4707), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n1052_adj_4731));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i908_1_lut (.I0(n1436), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1437));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i908_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4917));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_906_i32_4_lut (.I0(n1052_adj_4731), .I1(n99), 
            .I2(n1420), .I3(n558), .O(n32_adj_4954));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_906_i32_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35758_3_lut (.I0(n32_adj_4954), .I1(n95), .I2(n39_adj_4957), 
            .I3(GND_net), .O(n42605));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35758_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35759_3_lut (.I0(n42605), .I1(n94), .I2(n41_adj_4958), .I3(GND_net), 
            .O(n42606));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35759_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34704_4_lut (.I0(n41_adj_4958), .I1(n39_adj_4957), .I2(n37_adj_4956), 
            .I3(n40846), .O(n41551));
    defparam i34704_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_46_i890_3_lut_3_lut (.I0(n1316), .I1(n5979), .I2(n1299), 
            .I3(GND_net), .O(n1419_adj_4741));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i890_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i35308_3_lut (.I0(n34_adj_4955), .I1(n96), .I2(n37_adj_4956), 
            .I3(GND_net), .O(n42155));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35308_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35551_3_lut (.I0(n42606), .I1(n93), .I2(n43_adj_4959), .I3(GND_net), 
            .O(n42398));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35551_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35756_4_lut (.I0(n42398), .I1(n42155), .I2(n43_adj_4959), 
            .I3(n41551), .O(n42603));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35756_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 div_46_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4916));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35757_3_lut (.I0(n42603), .I1(n92), .I2(n1413), .I3(GND_net), 
            .O(n42604));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35757_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_46_i889_3_lut_3_lut (.I0(n1316), .I1(n5978), .I2(n1298), 
            .I3(GND_net), .O(n1418_adj_4740));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i889_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1810 (.I0(n42604), .I1(n15883), .I2(n91), .I3(n1412), 
            .O(n1436));
    defparam i1_4_lut_adj_1810.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_825_i45_2_lut (.I0(n1293), .I1(n93), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_4952));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_825_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4915));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_825_i39_2_lut (.I0(n1296), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_4948));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_825_i39_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_825_i43_2_lut (.I0(n1294), .I1(n94), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_4950));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_825_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_LessThan_825_i41_2_lut (.I0(n1295), .I1(n95), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4949));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_825_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i16_3_lut (.I0(encoder0_position[15]), .I1(n10_adj_4708), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n1051));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i827_1_lut (.I0(n1316), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1317));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i827_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_825_i34_4_lut (.I0(n1051), .I1(n99), .I2(n1299), 
            .I3(n558), .O(n34));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_825_i34_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35762_3_lut (.I0(n34), .I1(n95), .I2(n41_adj_4949), .I3(GND_net), 
            .O(n42609));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35762_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35763_3_lut (.I0(n42609), .I1(n94), .I2(n43_adj_4950), .I3(GND_net), 
            .O(n42610));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35763_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34714_4_lut (.I0(n43_adj_4950), .I1(n41_adj_4949), .I2(n39_adj_4948), 
            .I3(n40867), .O(n41561));
    defparam i34714_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 div_46_LessThan_825_i38_3_lut (.I0(n36_adj_4946), .I1(n96), 
            .I2(n39_adj_4948), .I3(GND_net), .O(n38_adj_4947));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_825_i38_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35547_3_lut (.I0(n42610), .I1(n93), .I2(n45_adj_4952), .I3(GND_net), 
            .O(n44_adj_4951));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35547_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35306_4_lut (.I0(n44_adj_4951), .I1(n38_adj_4947), .I2(n45_adj_4952), 
            .I3(n41561), .O(n42153));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35306_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1811 (.I0(n42153), .I1(n15880), .I2(n92), .I3(n1292), 
            .O(n1316));
    defparam i1_4_lut_adj_1811.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_LessThan_742_i41_2_lut (.I0(n1172), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4945));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_742_i41_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i17_3_lut (.I0(encoder0_position[16]), .I1(n9_adj_4695), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n1050));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i744_1_lut (.I0(n1193), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1194));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i744_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i891_3_lut_3_lut (.I0(n1316), .I1(n5980), .I2(n1051), 
            .I3(GND_net), .O(n1420));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i891_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_742_i36_4_lut (.I0(n1050), .I1(n99), .I2(n1175), 
            .I3(n558), .O(n36_adj_4942));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_742_i36_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_742_i40_3_lut (.I0(n38_adj_4943), .I1(n96), 
            .I2(n41_adj_4945), .I3(GND_net), .O(n40_adj_4944));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_742_i40_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35939_4_lut (.I0(n40_adj_4944), .I1(n36_adj_4942), .I2(n41_adj_4945), 
            .I3(n40889), .O(n42786));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35939_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35940_3_lut (.I0(n42786), .I1(n95), .I2(n1171), .I3(GND_net), 
            .O(n42787));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35940_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35869_3_lut (.I0(n42787), .I1(n94), .I2(n1170_adj_4738), 
            .I3(GND_net), .O(n42716));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35869_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 div_46_i887_3_lut_3_lut (.I0(n1316), .I1(n5976), .I2(n1296), 
            .I3(GND_net), .O(n1416));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i887_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1812 (.I0(n42716), .I1(n15877), .I2(n93), .I3(n1169), 
            .O(n1193));
    defparam i1_4_lut_adj_1812.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_i888_3_lut_3_lut (.I0(n1316), .I1(n5977), .I2(n1297), 
            .I3(GND_net), .O(n1417_adj_4739));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i888_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13163_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n13302), 
            .I3(GND_net), .O(n17902));   // verilog/coms.v(127[12] 295[6])
    defparam i13163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i886_3_lut_3_lut (.I0(n1316), .I1(n5975), .I2(n1295), 
            .I3(GND_net), .O(n1415));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i886_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_657_i43_2_lut (.I0(n1045), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n43));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_657_i43_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_i885_3_lut_3_lut (.I0(n1316), .I1(n5974), .I2(n1294), 
            .I3(GND_net), .O(n1414));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i885_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_mux_3_i18_3_lut (.I0(encoder0_position[17]), .I1(n8_adj_4696), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n1049));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i884_3_lut_3_lut (.I0(n1316), .I1(n5973), .I2(n1293), 
            .I3(GND_net), .O(n1413));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i884_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i659_1_lut (.I0(n1067), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n1068));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i659_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i883_3_lut_3_lut (.I0(n1316), .I1(n5972), .I2(n1292), 
            .I3(GND_net), .O(n1412));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i883_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4914));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34021_3_lut_4_lut (.I0(n1297), .I1(n97), .I2(n98), .I3(n1298), 
            .O(n40867));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34021_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_657_i38_4_lut (.I0(n1049), .I1(n99), .I2(n1048), 
            .I3(n558), .O(n38));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_657_i38_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_825_i36_3_lut_3_lut (.I0(n1297), .I1(n97), .I2(n98), 
            .I3(GND_net), .O(n36_adj_4946));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_825_i36_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_657_i42_3_lut (.I0(n40_adj_4936), .I1(n96), 
            .I2(n43), .I3(GND_net), .O(n42_adj_4937));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_657_i42_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 div_46_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4913));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35770_4_lut (.I0(n42_adj_4937), .I1(n38), .I2(n43), .I3(n40899), 
            .O(n42617));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35770_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35771_3_lut (.I0(n42617), .I1(n95), .I2(n1044), .I3(GND_net), 
            .O(n42618));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35771_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1813 (.I0(n42618), .I1(n15874), .I2(n94), .I3(n1043), 
            .O(n1067));
    defparam i1_4_lut_adj_1813.LUT_INIT = 16'hceef;
    SB_LUT4 div_46_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4912));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i22715_3_lut (.I0(n783), .I1(n97), .I2(n6_adj_4670), .I3(GND_net), 
            .O(n8_adj_4669));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i22715_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i22707_3_lut (.I0(n784), .I1(n98), .I2(n4_adj_4672), .I3(GND_net), 
            .O(n6_adj_4670));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i22707_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 div_46_LessThan_570_i45_2_lut (.I0(n915), .I1(n96), .I2(GND_net), 
            .I3(GND_net), .O(n45));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_570_i45_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 div_46_mux_3_i19_3_lut (.I0(encoder0_position[18]), .I1(n7_adj_4705), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n919));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22691_2_lut (.I0(n786), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i22691_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_i572_1_lut (.I0(n938), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n939));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i572_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_570_i40_4_lut (.I0(n919), .I1(n99), .I2(n918), 
            .I3(n558), .O(n40_adj_4821));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_570_i40_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 div_46_LessThan_570_i44_3_lut (.I0(n42_adj_4822), .I1(n96), 
            .I2(n45), .I3(GND_net), .O(n44));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_570_i44_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i35286_4_lut (.I0(n44), .I1(n40_adj_4821), .I2(n45), .I3(n40949), 
            .O(n42133));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35286_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i1_4_lut_adj_1814 (.I0(n42133), .I1(n15864), .I2(n95), .I3(n914), 
            .O(n938));
    defparam i1_4_lut_adj_1814.LUT_INIT = 16'hceef;
    SB_LUT4 i22747_3_lut (.I0(n648), .I1(n98), .I2(n4_adj_5269), .I3(GND_net), 
            .O(n6_adj_5253));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i22747_3_lut.LUT_INIT = 16'he8e8;
    SB_LUT4 i22731_2_lut (.I0(n650), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_5273));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i22731_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_mux_3_i20_3_lut (.I0(encoder0_position[19]), .I1(n6_adj_4706), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n786));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i483_1_lut (.I0(n806), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n807));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i483_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_481_i42_4_lut (.I0(n786), .I1(n99), .I2(n785), 
            .I3(n558), .O(n42_adj_4778));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_481_i42_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35742_3_lut (.I0(n42_adj_4778), .I1(n98), .I2(n784), .I3(GND_net), 
            .O(n42589));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35742_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i35743_3_lut (.I0(n42589), .I1(n97), .I2(n783), .I3(GND_net), 
            .O(n42590));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35743_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1815 (.I0(n42590), .I1(n15971), .I2(n96), .I3(n35865), 
            .O(n806));
    defparam i1_4_lut_adj_1815.LUT_INIT = 16'hefce;
    SB_LUT4 i36042_2_lut (.I0(blink), .I1(n25734), .I2(GND_net), .I3(GND_net), 
            .O(blink_N_255));
    defparam i36042_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 i13164_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n13302), 
            .I3(GND_net), .O(n17903));   // verilog/coms.v(127[12] 295[6])
    defparam i13164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13165_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n13302), .I3(GND_net), .O(n17904));   // verilog/coms.v(127[12] 295[6])
    defparam i13165_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22763_2_lut (.I0(n511), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_5268));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i22763_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_mux_3_i21_3_lut (.I0(encoder0_position[20]), .I1(n5_adj_4692), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n650));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i392_1_lut (.I0(n671), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n672));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i392_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_390_i44_4_lut (.I0(n650), .I1(n99), .I2(n649), 
            .I3(n558), .O(n44_adj_4842));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_390_i44_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i35294_3_lut (.I0(n44_adj_4842), .I1(n98), .I2(n648), .I3(GND_net), 
            .O(n42141));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i35294_3_lut.LUT_INIT = 16'h2b2b;
    SB_LUT4 i1_4_lut_adj_1816 (.I0(n42141), .I1(n15966), .I2(n97), .I3(n35825), 
            .O(n671));
    defparam i1_4_lut_adj_1816.LUT_INIT = 16'hefce;
    SB_LUT4 i1_2_lut_adj_1817 (.I0(n2356), .I1(n2358_adj_4940), .I2(GND_net), 
            .I3(GND_net), .O(n38171));
    defparam i1_2_lut_adj_1817.LUT_INIT = 16'heeee;
    SB_LUT4 i13166_3_lut (.I0(\data_out_frame[18] [1]), .I1(displacement[17]), 
            .I2(n13302), .I3(GND_net), .O(n17905));   // verilog/coms.v(127[12] 295[6])
    defparam i13166_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13440_3_lut (.I0(encoder0_position[23]), .I1(n2993), .I2(count_enable), 
            .I3(GND_net), .O(n18179));   // quad.v(35[10] 41[6])
    defparam i13440_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i22787_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n2_adj_5323));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i22787_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 div_46_mux_3_i22_3_lut (.I0(encoder0_position[21]), .I1(n4_adj_4693), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n511));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i299_1_lut (.I0(n533), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n534));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i299_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_LessThan_297_i46_4_lut (.I0(n511), .I1(n99), .I2(n510), 
            .I3(n558), .O(n46));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_297_i46_4_lut.LUT_INIT = 16'h0317;
    SB_LUT4 i1_4_lut_adj_1818 (.I0(n46), .I1(n15996), .I2(n98), .I3(n35676), 
            .O(n533));
    defparam i1_4_lut_adj_1818.LUT_INIT = 16'hefce;
    SB_LUT4 div_46_mux_3_i23_3_lut (.I0(encoder0_position[22]), .I1(n3_adj_4694), 
            .I2(encoder0_position[23]), .I3(GND_net), .O(n369));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i204_1_lut (.I0(n392), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i204_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34174_2_lut (.I0(n369), .I1(n558), .I2(GND_net), .I3(GND_net), 
            .O(n40651));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34174_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_4_lut_adj_1819 (.I0(n40651), .I1(n16003), .I2(n99), .I3(n5_adj_5242), 
            .O(n392));
    defparam i1_4_lut_adj_1819.LUT_INIT = 16'hefce;
    SB_LUT4 div_46_mux_5_i23_3_lut (.I0(gearBoxRatio[22]), .I1(n53), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n78));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i23_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1820 (.I0(n78), .I1(n77), .I2(GND_net), .I3(GND_net), 
            .O(n15910));
    defparam i1_2_lut_adj_1820.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i22_3_lut (.I0(gearBoxRatio[21]), .I1(n54), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n79));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i22_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i21_3_lut (.I0(gearBoxRatio[20]), .I1(n55), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n80));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i21_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i20_3_lut (.I0(gearBoxRatio[19]), .I1(n56), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n81));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i20_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1821 (.I0(n81), .I1(n15987), .I2(GND_net), .I3(GND_net), 
            .O(n15983));
    defparam i1_2_lut_adj_1821.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i19_3_lut (.I0(gearBoxRatio[18]), .I1(n57), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n82));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i19_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i18_3_lut (.I0(gearBoxRatio[17]), .I1(n58), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n83));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i18_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i17_3_lut (.I0(gearBoxRatio[16]), .I1(n59), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n84));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i17_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1822 (.I0(n84), .I1(n15901), .I2(GND_net), .I3(GND_net), 
            .O(n15897));
    defparam i1_2_lut_adj_1822.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i16_3_lut (.I0(gearBoxRatio[15]), .I1(n60), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n85));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i16_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i15_3_lut (.I0(gearBoxRatio[14]), .I1(n61), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n86));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i15_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i14_3_lut (.I0(gearBoxRatio[13]), .I1(n62), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n87));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i14_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1823 (.I0(n87), .I1(n15893), .I2(GND_net), .I3(GND_net), 
            .O(n15977));
    defparam i1_2_lut_adj_1823.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_mux_5_i13_3_lut (.I0(gearBoxRatio[12]), .I1(n63), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n88));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i13_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i12_3_lut (.I0(gearBoxRatio[11]), .I1(n64), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n89));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i12_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_i970_3_lut_3_lut (.I0(n1436), .I1(n5991), .I2(n1420), 
            .I3(GND_net), .O(n1537));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i970_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_mux_5_i11_3_lut (.I0(gearBoxRatio[10]), .I1(n65), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n90));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i11_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1824 (.I0(n90), .I1(n15974), .I2(GND_net), .I3(GND_net), 
            .O(n15883));
    defparam i1_2_lut_adj_1824.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_i964_3_lut_3_lut (.I0(n1436), .I1(n5985), .I2(n1414), 
            .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i964_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_mux_5_i10_3_lut (.I0(gearBoxRatio[9]), .I1(n66), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n91));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i10_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i9_3_lut (.I0(gearBoxRatio[8]), .I1(n67), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n92));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i9_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i8_3_lut (.I0(gearBoxRatio[7]), .I1(n68), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n93));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i8_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1825 (.I0(n93), .I1(n15877), .I2(GND_net), .I3(GND_net), 
            .O(n15874));
    defparam i1_2_lut_adj_1825.LUT_INIT = 16'hdddd;
    SB_LUT4 unary_minus_28_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_mux_5_i7_3_lut (.I0(gearBoxRatio[6]), .I1(n69), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n94));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i7_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 unary_minus_28_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_mux_5_i6_3_lut (.I0(gearBoxRatio[5]), .I1(n70), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n95));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i6_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_mux_5_i5_3_lut (.I0(gearBoxRatio[4]), .I1(n71), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n96));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 unary_minus_28_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1826 (.I0(n96), .I1(n15971), .I2(GND_net), .I3(GND_net), 
            .O(n15966));
    defparam i1_2_lut_adj_1826.LUT_INIT = 16'hdddd;
    SB_LUT4 div_46_i968_3_lut_3_lut (.I0(n1436), .I1(n5989), .I2(n1418_adj_4740), 
            .I3(GND_net), .O(n1535));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i968_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_mux_5_i4_3_lut (.I0(gearBoxRatio[3]), .I1(n72), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n97));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i4_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 unary_minus_28_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4663));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i12802_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n23989), 
            .I3(n15851), .O(n17541));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12802_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 div_46_mux_5_i3_3_lut (.I0(gearBoxRatio[2]), .I1(n73), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n98));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i3_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 unary_minus_28_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_mux_5_i2_3_lut (.I0(gearBoxRatio[1]), .I1(n74), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n99));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 unary_minus_28_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18_adj_4662));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i969_3_lut_3_lut (.I0(n1436), .I1(n5990), .I2(n1419_adj_4741), 
            .I3(GND_net), .O(n1536));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i969_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_mux_5_i1_3_lut (.I0(gearBoxRatio[0]), .I1(n75), .I2(gearBoxRatio[23]), 
            .I3(GND_net), .O(n558));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_mux_5_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 div_46_i967_3_lut_3_lut (.I0(n1436), .I1(n5988), .I2(n1417_adj_4739), 
            .I3(GND_net), .O(n1534));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i967_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 unary_minus_28_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4661));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4660));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36790_2_lut (.I0(encoder0_position[23]), .I1(gearBoxRatio[23]), 
            .I2(GND_net), .I3(GND_net), .O(n43635));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i36790_2_lut.LUT_INIT = 16'h9999;
    SB_LUT4 unary_minus_28_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_mux_3_i3_3_lut (.I0(communication_counter[2]), .I1(n31), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3358));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4659));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2219_3_lut (.I0(n3258), .I1(n3325), .I2(n3263), .I3(GND_net), 
            .O(n3357));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2218_3_lut (.I0(n3257), .I1(n3324), .I2(n3263), .I3(GND_net), 
            .O(n3356));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2218_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i963_3_lut_3_lut (.I0(n1436), .I1(n5984), .I2(n1413), 
            .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i963_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 unary_minus_28_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2217_3_lut (.I0(n3256), .I1(n3323), .I2(n3263), .I3(GND_net), 
            .O(n3355));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2216_3_lut (.I0(n3255), .I1(n3322), .I2(n3263), .I3(GND_net), 
            .O(n3354));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34844_3_lut (.I0(n3051), .I1(n3118), .I2(n3065), .I3(GND_net), 
            .O(n3150));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i34844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34845_3_lut (.I0(n3150), .I1(n3217), .I2(n3164), .I3(GND_net), 
            .O(n3249));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i34845_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2140_3_lut (.I0(n3147), .I1(n3214), .I2(n3164), .I3(GND_net), 
            .O(n3246));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2140_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2130_3_lut (.I0(n3137), .I1(n3204), .I2(n3164), .I3(GND_net), 
            .O(n3236));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2130_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i971_3_lut_3_lut (.I0(n1436), .I1(n5992), .I2(n1052_adj_4731), 
            .I3(GND_net), .O(n1538));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i971_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i2127_3_lut (.I0(n3134), .I1(n3201), .I2(n3164), .I3(GND_net), 
            .O(n3233));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2127_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2129_3_lut (.I0(n3136), .I1(n3203), .I2(n3164), .I3(GND_net), 
            .O(n3235));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2129_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2126_3_lut (.I0(n3133), .I1(n3200), .I2(n3164), .I3(GND_net), 
            .O(n3232));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2135_3_lut (.I0(n3142), .I1(n3209), .I2(n3164), .I3(GND_net), 
            .O(n3241));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2135_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2134_3_lut (.I0(n3141), .I1(n3208), .I2(n3164), .I3(GND_net), 
            .O(n3240));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2134_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2133_3_lut (.I0(n3140), .I1(n3207), .I2(n3164), .I3(GND_net), 
            .O(n3239));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2133_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2132_3_lut (.I0(n3139), .I1(n3206), .I2(n3164), .I3(GND_net), 
            .O(n3238));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2132_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2131_3_lut (.I0(n3138), .I1(n3205), .I2(n3164), .I3(GND_net), 
            .O(n3237));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2131_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2128_3_lut (.I0(n3135), .I1(n3202), .I2(n3164), .I3(GND_net), 
            .O(n3234));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2128_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35483_3_lut (.I0(n3046), .I1(n3113), .I2(n3065), .I3(GND_net), 
            .O(n3145));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i35483_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35293_3_lut (.I0(n3145), .I1(n3212), .I2(n3164), .I3(GND_net), 
            .O(n3244));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i35293_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2139_3_lut (.I0(n3146), .I1(n3213), .I2(n3164), .I3(GND_net), 
            .O(n3245));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2139_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2147_3_lut (.I0(n3154), .I1(n3221), .I2(n3164), .I3(GND_net), 
            .O(n3253));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2141_3_lut (.I0(n3148), .I1(n3215), .I2(n3164), .I3(GND_net), 
            .O(n3247));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2125_3_lut (.I0(n3132), .I1(n3199), .I2(n3164), .I3(GND_net), 
            .O(n3231));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2125_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2146_3_lut (.I0(n3153), .I1(n3220), .I2(n3164), .I3(GND_net), 
            .O(n3252));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2137_3_lut (.I0(n3144), .I1(n3211), .I2(n3164), .I3(GND_net), 
            .O(n3243));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2137_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35290_3_lut (.I0(n38584), .I1(n2852), .I2(n41601), .I3(GND_net), 
            .O(n3149));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i35290_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35291_3_lut (.I0(n3149), .I1(n3216), .I2(n3164), .I3(GND_net), 
            .O(n3248));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i35291_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2145_3_lut (.I0(n3152), .I1(n3219), .I2(n3164), .I3(GND_net), 
            .O(n3251));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2136_3_lut (.I0(n3143), .I1(n3210), .I2(n3164), .I3(GND_net), 
            .O(n3242));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2136_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2149_3_lut (.I0(n3156), .I1(n3223), .I2(n3164), .I3(GND_net), 
            .O(n3255));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34842_3_lut (.I0(n3052), .I1(n3119), .I2(n3065), .I3(GND_net), 
            .O(n3151));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i34842_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34843_3_lut (.I0(n3151), .I1(n3218), .I2(n3164), .I3(GND_net), 
            .O(n3250));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i34843_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2072_3_lut (.I0(n3047), .I1(n3114), .I2(n3065), .I3(GND_net), 
            .O(n3146));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2072_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i966_3_lut_3_lut (.I0(n1436), .I1(n5987), .I2(n1416), 
            .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i966_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i2073_3_lut (.I0(n3048), .I1(n3115), .I2(n3065), .I3(GND_net), 
            .O(n3147));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2073_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2070_3_lut (.I0(n3045), .I1(n3112), .I2(n3065), .I3(GND_net), 
            .O(n3144));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2058_3_lut (.I0(n3033), .I1(n3100), .I2(n3065), .I3(GND_net), 
            .O(n3132));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2058_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_28_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4658));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_28_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(149[23:28])
    defparam unary_minus_28_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2079_3_lut (.I0(n3054), .I1(n3121), .I2(n3065), .I3(GND_net), 
            .O(n3153));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i965_3_lut_3_lut (.I0(n1436), .I1(n5986), .I2(n1415), 
            .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i965_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i2074_3_lut (.I0(n3049), .I1(n3116), .I2(n3065), .I3(GND_net), 
            .O(n3148));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2074_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35298_3_lut (.I0(n2947_adj_4655), .I1(n3014_adj_4749), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3046));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i35298_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1827 (.I0(n2354), .I1(n38171), .I2(n2355), .I3(n2357_adj_4941), 
            .O(n36008));
    defparam i1_4_lut_adj_1827.LUT_INIT = 16'ha080;
    SB_LUT4 rem_4_i2069_3_lut (.I0(n3044), .I1(n3111), .I2(n3065), .I3(GND_net), 
            .O(n3143));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13439_3_lut (.I0(encoder0_position[22]), .I1(n2994), .I2(count_enable), 
            .I3(GND_net), .O(n18178));   // quad.v(35[10] 41[6])
    defparam i13439_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13438_3_lut (.I0(encoder0_position[21]), .I1(n2995), .I2(count_enable), 
            .I3(GND_net), .O(n18177));   // quad.v(35[10] 41[6])
    defparam i13438_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2066_3_lut (.I0(n3041), .I1(n3108), .I2(n3065), .I3(GND_net), 
            .O(n3140));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2065_3_lut (.I0(n3040), .I1(n3107), .I2(n3065), .I3(GND_net), 
            .O(n3139));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2065_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2064_3_lut (.I0(n3039), .I1(n3106), .I2(n3065), .I3(GND_net), 
            .O(n3138));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2062_3_lut (.I0(n3037), .I1(n3104), .I2(n3065), .I3(GND_net), 
            .O(n3136));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2062_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2063_3_lut (.I0(n3038), .I1(n3105), .I2(n3065), .I3(GND_net), 
            .O(n3137));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2061_3_lut (.I0(n3036), .I1(n3103), .I2(n3065), .I3(GND_net), 
            .O(n3135));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2061_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2060_3_lut (.I0(n3035), .I1(n3102), .I2(n3065), .I3(GND_net), 
            .O(n3134));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2060_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2059_3_lut (.I0(n3034), .I1(n3101), .I2(n3065), .I3(GND_net), 
            .O(n3133));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2059_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2081_3_lut (.I0(n3056), .I1(n3123), .I2(n3065), .I3(GND_net), 
            .O(n3155));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2080_3_lut (.I0(n3055), .I1(n3122), .I2(n3065), .I3(GND_net), 
            .O(n3154));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2067_3_lut (.I0(n3042), .I1(n3109), .I2(n3065), .I3(GND_net), 
            .O(n3141));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34754_3_lut (.I0(n3065), .I1(n2966_adj_4763), .I2(n2867), 
            .I3(GND_net), .O(n41601));
    defparam i34754_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 rem_4_i1941_rep_26_3_lut (.I0(n2919), .I1(n3018), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n38596));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1941_rep_26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2008_rep_14_3_lut (.I0(n38596), .I1(n3117), .I2(n3065), 
            .I3(GND_net), .O(n38584));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2008_rep_14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2068_3_lut (.I0(n3043), .I1(n3110), .I2(n3065), .I3(GND_net), 
            .O(n3142));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2068_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2078_3_lut (.I0(n3053), .I1(n3120), .I2(n3065), .I3(GND_net), 
            .O(n3152));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1991_3_lut (.I0(n2934), .I1(n3001_adj_4762), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13437_3_lut (.I0(encoder0_position[20]), .I1(n2996), .I2(count_enable), 
            .I3(GND_net), .O(n18176));   // quad.v(35[10] 41[6])
    defparam i13437_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34852_3_lut (.I0(n2847), .I1(n2914), .I2(n2867), .I3(GND_net), 
            .O(n2946_adj_4776));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i34852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34853_3_lut (.I0(n2946_adj_4776), .I1(n3013_adj_4750), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3045));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i34853_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13451_3_lut (.I0(encoder1_position[10]), .I1(n2956), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18190));   // quad.v(35[10] 41[6])
    defparam i13451_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2002_3_lut (.I0(n2945_adj_4654), .I1(n3012_adj_4751), 
            .I2(n2966_adj_4763), .I3(GND_net), .O(n3044));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2002_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34850_3_lut (.I0(n2852), .I1(n2919), .I2(n2867), .I3(GND_net), 
            .O(n2951_adj_4772));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i34850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34851_3_lut (.I0(n2951_adj_4772), .I1(n3018), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3050));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i34851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2007_3_lut (.I0(n2950_adj_4773), .I1(n3017), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3049));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2009_rep_17_3_lut (.I0(n2952_adj_4771), .I1(n3019), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3051));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2009_rep_17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2006_3_lut (.I0(n2949_adj_4774), .I1(n3016_adj_4747), 
            .I2(n2966_adj_4763), .I3(GND_net), .O(n3048));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2006_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2005_3_lut (.I0(n2948_adj_4775), .I1(n3015_adj_4748), 
            .I2(n2966_adj_4763), .I3(GND_net), .O(n3047));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2005_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2011_3_lut (.I0(n2954_adj_4769), .I1(n3021), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3053));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1995_3_lut (.I0(n2938), .I1(n3005_adj_4758), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3037));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1993_3_lut (.I0(n2936), .I1(n3003_adj_4760), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3035));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1994_3_lut (.I0(n2937), .I1(n3004_adj_4759), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3036));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1992_3_lut (.I0(n2935), .I1(n3002_adj_4761), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3034));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2001_3_lut (.I0(n2944_adj_4777), .I1(n3011_adj_4752), 
            .I2(n2966_adj_4763), .I3(GND_net), .O(n3043));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2010_rep_15_3_lut (.I0(n2953_adj_4770), .I1(n3020), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3052));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2010_rep_15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1999_3_lut (.I0(n2942), .I1(n3009_adj_4754), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3041));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1997_3_lut (.I0(n2940), .I1(n3007_adj_4756), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3039));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1998_3_lut (.I0(n2941), .I1(n3008_adj_4755), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3040));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1996_3_lut (.I0(n2939), .I1(n3006_adj_4757), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3038));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2013_3_lut (.I0(n2956_adj_4767), .I1(n3023), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3055));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2000_3_lut (.I0(n2943_adj_4656), .I1(n3010_adj_4753), 
            .I2(n2966_adj_4763), .I3(GND_net), .O(n3042));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2000_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2012_3_lut (.I0(n2955_adj_4768), .I1(n3022), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3054));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35539_3_lut (.I0(n2846), .I1(n2913), .I2(n2867), .I3(GND_net), 
            .O(n2945_adj_4654));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i35539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1934_3_lut (.I0(n2845), .I1(n2912), .I2(n2867), .I3(GND_net), 
            .O(n2944_adj_4777));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13450_3_lut (.I0(encoder1_position[9]), .I1(n2957), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18189));   // quad.v(35[10] 41[6])
    defparam i13450_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13449_3_lut (.I0(encoder1_position[8]), .I1(n2958), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18188));   // quad.v(35[10] 41[6])
    defparam i13449_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13448_3_lut (.I0(encoder1_position[7]), .I1(n2959), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18187));   // quad.v(35[10] 41[6])
    defparam i13448_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1933_3_lut (.I0(n2844), .I1(n2911), .I2(n2867), .I3(GND_net), 
            .O(n2943_adj_4656));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1933_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13447_3_lut (.I0(encoder1_position[6]), .I1(n2960), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18186));   // quad.v(35[10] 41[6])
    defparam i13447_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1940_3_lut (.I0(n2851), .I1(n2918), .I2(n2867), .I3(GND_net), 
            .O(n2950_adj_4773));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1940_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i962_3_lut_3_lut (.I0(n1436), .I1(n5983), .I2(n1412), 
            .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i962_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1943_3_lut (.I0(n2854), .I1(n2921), .I2(n2867), .I3(GND_net), 
            .O(n2953_adj_4770));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1943_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34000_3_lut_4_lut (.I0(n1418_adj_4740), .I1(n97), .I2(n98), 
            .I3(n1419_adj_4741), .O(n40846));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i34000_3_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 rem_4_i1942_3_lut (.I0(n2853), .I1(n2920), .I2(n2867), .I3(GND_net), 
            .O(n2952_adj_4771));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1942_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1939_3_lut (.I0(n2850), .I1(n2917), .I2(n2867), .I3(GND_net), 
            .O(n2949_adj_4774));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1939_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1937_rep_22_3_lut (.I0(n2848), .I1(n2915), .I2(n2867), 
            .I3(GND_net), .O(n2947_adj_4655));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1937_rep_22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1932_3_lut (.I0(n2843), .I1(n2910), .I2(n2867), .I3(GND_net), 
            .O(n2942));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1932_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1931_3_lut (.I0(n2842), .I1(n2909), .I2(n2867), .I3(GND_net), 
            .O(n2941));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1926_3_lut (.I0(n2837), .I1(n2904), .I2(n2867), .I3(GND_net), 
            .O(n2936));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1925_3_lut (.I0(n2836), .I1(n2903), .I2(n2867), .I3(GND_net), 
            .O(n2935));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1924_3_lut (.I0(n2835), .I1(n2902), .I2(n2867), .I3(GND_net), 
            .O(n2934));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1930_3_lut (.I0(n2841), .I1(n2908), .I2(n2867), .I3(GND_net), 
            .O(n2940));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1930_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1928_3_lut (.I0(n2839), .I1(n2906), .I2(n2867), .I3(GND_net), 
            .O(n2938));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1929_3_lut (.I0(n2840), .I1(n2907), .I2(n2867), .I3(GND_net), 
            .O(n2939));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1929_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1927_3_lut (.I0(n2838), .I1(n2905), .I2(n2867), .I3(GND_net), 
            .O(n2937));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1945_3_lut (.I0(n2856), .I1(n2923), .I2(n2867), .I3(GND_net), 
            .O(n2955_adj_4768));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1938_3_lut (.I0(n2849), .I1(n2916), .I2(n2867), .I3(GND_net), 
            .O(n2948_adj_4775));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1938_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1944_3_lut (.I0(n2855), .I1(n2922), .I2(n2867), .I3(GND_net), 
            .O(n2954_adj_4769));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1947_3_lut (.I0(n2858), .I1(n2925), .I2(n2867), .I3(GND_net), 
            .O(n2957_adj_4765));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1947_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1828 (.I0(n2353), .I1(n2349), .I2(n2350), .I3(n2352), 
            .O(n28));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i12_4_lut_adj_1828.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_LessThan_906_i34_3_lut_3_lut (.I0(n1418_adj_4740), .I1(n97), 
            .I2(n98), .I3(GND_net), .O(n34_adj_4955));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_906_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 rem_4_i1946_3_lut (.I0(n2857), .I1(n2924), .I2(n2867), .I3(GND_net), 
            .O(n2956_adj_4767));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1829 (.I0(n2956_adj_4767), .I1(n2957_adj_4765), 
            .I2(n2958_adj_4764), .I3(GND_net), .O(n36043));
    defparam i1_3_lut_adj_1829.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1830 (.I0(n2954_adj_4769), .I1(n2948_adj_4775), 
            .I2(n36043), .I3(n2955_adj_4768), .O(n28_adj_5356));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i6_4_lut_adj_1830.LUT_INIT = 16'heccc;
    SB_LUT4 i13_4_lut_adj_1831 (.I0(n2937), .I1(n2939), .I2(n2938), .I3(n2940), 
            .O(n35_adj_5354));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i13_4_lut_adj_1831.LUT_INIT = 16'hfffe;
    SB_LUT4 i13446_3_lut (.I0(encoder1_position[5]), .I1(n2961), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18185));   // quad.v(35[10] 41[6])
    defparam i13446_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1832 (.I0(n2934), .I1(n2935), .I2(n2933), .I3(n2936), 
            .O(n34_adj_5355));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i12_4_lut_adj_1832.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1833 (.I0(n35_adj_5354), .I1(n2941), .I2(n28_adj_5356), 
            .I3(n2942), .O(n40_adj_5342));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i18_4_lut_adj_1833.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n2947_adj_4655), .I1(n2949_adj_4774), .I2(n2952_adj_4771), 
            .I3(n2953_adj_4770), .O(n38_adj_5344));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_3_lut (.I0(n2951_adj_4772), .I1(n34_adj_5355), .I2(n2950_adj_4773), 
            .I3(GND_net), .O(n39_adj_5343));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1834 (.I0(n2943_adj_4656), .I1(n2944_adj_4777), 
            .I2(n2945_adj_4654), .I3(n2946_adj_4776), .O(n37_adj_5347));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i15_4_lut_adj_1834.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1835 (.I0(n37_adj_5347), .I1(n39_adj_5343), .I2(n38_adj_5344), 
            .I3(n40_adj_5342), .O(n2966_adj_4763));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i21_4_lut_adj_1835.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i7_3_lut (.I0(communication_counter[6]), .I1(n27_adj_4782), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2958_adj_4764));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2015_3_lut (.I0(n2958_adj_4764), .I1(n3025), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3057));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2014_3_lut (.I0(n2957_adj_4765), .I1(n3024), .I2(n2966_adj_4763), 
            .I3(GND_net), .O(n3056));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13445_3_lut (.I0(encoder1_position[4]), .I1(n2962), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n18184));   // quad.v(35[10] 41[6])
    defparam i13445_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1836 (.I0(n3056), .I1(n3057), .I2(n3058), .I3(GND_net), 
            .O(n36105));
    defparam i1_3_lut_adj_1836.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1837 (.I0(n3054), .I1(n3042), .I2(n36105), .I3(n3055), 
            .O(n29_adj_4730));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i6_4_lut_adj_1837.LUT_INIT = 16'heccc;
    SB_LUT4 div_46_i1048_3_lut_3_lut (.I0(n1553_adj_4742), .I1(n6004), .I2(n1538), 
            .I3(GND_net), .O(n1652));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1048_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14_4_lut_adj_1838 (.I0(n3038), .I1(n3040), .I2(n3039), .I3(n3041), 
            .O(n37));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i14_4_lut_adj_1838.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1839 (.I0(n3034), .I1(n3036), .I2(n3035), .I3(n3037), 
            .O(n36));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i13_4_lut_adj_1839.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1042_3_lut_3_lut (.I0(n1553_adj_4742), .I1(n5998), .I2(n1532), 
            .I3(GND_net), .O(n1646));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1042_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i19_4_lut (.I0(n37), .I1(n29_adj_4730), .I2(n3052), .I3(n3043), 
            .O(n42));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n3053), .I1(n3047), .I2(n3048), .I3(n3051), 
            .O(n40));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1840 (.I0(n3045), .I1(n36), .I2(n3033), .I3(n3032), 
            .O(n41));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i18_4_lut_adj_1840.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1841 (.I0(n3049), .I1(n3050), .I2(n3044), .I3(n3046), 
            .O(n39));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i16_4_lut_adj_1841.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1842 (.I0(n39), .I1(n41), .I2(n40), .I3(n42), 
            .O(n3065));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i22_4_lut_adj_1842.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i6_3_lut (.I0(communication_counter[5]), .I1(n28_adj_4781), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3058));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2083_3_lut (.I0(n3058), .I1(n3125), .I2(n3065), .I3(GND_net), 
            .O(n3157));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2082_3_lut (.I0(n3057), .I1(n3124), .I2(n3065), .I3(GND_net), 
            .O(n3156));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2082_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1843 (.I0(n3156), .I1(n3157), .I2(n3158), .I3(GND_net), 
            .O(n36053));
    defparam i1_3_lut_adj_1843.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1844 (.I0(n3141), .I1(n3154), .I2(n36053), .I3(n3155), 
            .O(n30_adj_5352));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i6_4_lut_adj_1844.LUT_INIT = 16'heaaa;
    SB_LUT4 i16_4_lut_adj_1845 (.I0(n3150), .I1(n3152), .I2(n3142), .I3(n3149), 
            .O(n40_adj_5350));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i16_4_lut_adj_1845.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_2_lut (.I0(n3133), .I1(n3134), .I2(GND_net), .I3(GND_net), 
            .O(n26_adj_5353));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i14_4_lut_adj_1846 (.I0(n3135), .I1(n3137), .I2(n3136), .I3(n3138), 
            .O(n38_adj_5351));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i14_4_lut_adj_1846.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut (.I0(n3139), .I1(n40_adj_5350), .I2(n30_adj_5352), 
            .I3(n3140), .O(n44_adj_5345));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1847 (.I0(n3143), .I1(n3145), .I2(n3148), .I3(n3153), 
            .O(n42_adj_5348));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i18_4_lut_adj_1847.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1848 (.I0(n3132), .I1(n38_adj_5351), .I2(n26_adj_5353), 
            .I3(n3131), .O(n43_adj_5346));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i19_4_lut_adj_1848.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1849 (.I0(n3144), .I1(n3147), .I2(n3151), .I3(n3146), 
            .O(n41_adj_5349));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i17_4_lut_adj_1849.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(n41_adj_5349), .I1(n43_adj_5346), .I2(n42_adj_5348), 
            .I3(n44_adj_5345), .O(n3164));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i5_3_lut (.I0(communication_counter[4]), .I1(n29_adj_4780), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3158));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_mux_3_i4_3_lut (.I0(communication_counter[3]), .I1(n30), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3258));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2151_3_lut (.I0(n3158), .I1(n3225), .I2(n3164), .I3(GND_net), 
            .O(n3257));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2150_3_lut (.I0(n3157), .I1(n3224), .I2(n3164), .I3(GND_net), 
            .O(n3256));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1850 (.I0(n3256), .I1(n3257), .I2(n3258), .I3(GND_net), 
            .O(n36110));
    defparam i1_3_lut_adj_1850.LUT_INIT = 16'hfefe;
    SB_LUT4 i7_4_lut_adj_1851 (.I0(n3254), .I1(n3250), .I2(n36110), .I3(n3255), 
            .O(n32_adj_5313));
    defparam i7_4_lut_adj_1851.LUT_INIT = 16'heccc;
    SB_LUT4 i17_4_lut_adj_1852 (.I0(n3242), .I1(n3251), .I2(n3248), .I3(n3243), 
            .O(n42_adj_5309));
    defparam i17_4_lut_adj_1852.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1853 (.I0(n2343), .I1(n2345), .I2(n2344), .I3(n36008), 
            .O(n26));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i10_4_lut_adj_1853.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1854 (.I0(n2346), .I1(n2351), .I2(n2347), .I3(n2348), 
            .O(n27));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i11_4_lut_adj_1854.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1855 (.I0(n2340), .I1(n2341), .I2(n2339), .I3(n2342), 
            .O(n25_adj_4667));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i9_4_lut_adj_1855.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1856 (.I0(n25_adj_4667), .I1(n27), .I2(n26), 
            .I3(n28), .O(n2372_adj_4939));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i15_4_lut_adj_1856.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1047_3_lut_3_lut (.I0(n1553_adj_4742), .I1(n6003), .I2(n1537), 
            .I3(GND_net), .O(n1651));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1047_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_71_i1_4_lut (.I0(encoder1_position[0]), .I1(displacement[0]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[0]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12_3_lut_adj_1857 (.I0(bit_ctr[8]), .I1(n40707), .I2(n4483), 
            .I3(GND_net), .O(n33633));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1857.LUT_INIT = 16'hacac;
    SB_LUT4 mux_70_i1_3_lut (.I0(encoder0_position[0]), .I1(motor_state_23__N_106[0]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1539_3_lut (.I0(n2258), .I1(n2325), .I2(n2273_adj_4953), 
            .I3(GND_net), .O(n2357_adj_4941));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1539_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i2_4_lut (.I0(encoder1_position[1]), .I1(displacement[1]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[1]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i2_3_lut (.I0(encoder0_position[1]), .I1(motor_state_23__N_106[1]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1046_3_lut_3_lut (.I0(n1553_adj_4742), .I1(n6002), .I2(n1536), 
            .I3(GND_net), .O(n1650));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1046_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1045_3_lut_3_lut (.I0(n1553_adj_4742), .I1(n6001), .I2(n1535), 
            .I3(GND_net), .O(n1649));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1045_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1041_3_lut_3_lut (.I0(n1553_adj_4742), .I1(n5997), .I2(n1531), 
            .I3(GND_net), .O(n1645));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1041_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_71_i3_4_lut (.I0(encoder1_position[2]), .I1(displacement[2]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[2]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12_3_lut_adj_1858 (.I0(bit_ctr[7]), .I1(n40706), .I2(n4483), 
            .I3(GND_net), .O(n33631));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1858.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1049_3_lut_3_lut (.I0(n1553_adj_4742), .I1(n6005), .I2(n1053_adj_4732), 
            .I3(GND_net), .O(n1653));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1049_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1044_3_lut_3_lut (.I0(n1553_adj_4742), .I1(n6000), .I2(n1534), 
            .I3(GND_net), .O(n1648));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1044_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1043_3_lut_3_lut (.I0(n1553_adj_4742), .I1(n5999), .I2(n1533), 
            .I3(GND_net), .O(n1647));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1043_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_70_i3_3_lut (.I0(encoder0_position[2]), .I1(motor_state_23__N_106[2]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1040_3_lut_3_lut (.I0(n1553_adj_4742), .I1(n5996), .I2(n1530), 
            .I3(GND_net), .O(n1644));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1040_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13520_3_lut (.I0(\half_duty[0] [7]), .I1(half_duty_new[7]), 
            .I2(n1170), .I3(GND_net), .O(n18259));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1039_3_lut_3_lut (.I0(n1553_adj_4742), .I1(n5995), .I2(n1529), 
            .I3(GND_net), .O(n1643));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1039_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13519_3_lut (.I0(\half_duty[0] [6]), .I1(half_duty_new[6]), 
            .I2(n1170), .I3(GND_net), .O(n18258));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13519_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i4_4_lut (.I0(encoder1_position[3]), .I1(displacement[3]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[3]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 rem_4_mux_3_i12_3_lut (.I0(communication_counter[11]), .I1(n22_adj_4787), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2458_adj_4875));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_70_i4_3_lut (.I0(encoder0_position[3]), .I1(motor_state_23__N_106[3]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1123_3_lut_3_lut (.I0(n1667), .I1(n6017), .I2(n1652), 
            .I3(GND_net), .O(n1763));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1123_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_71_i5_4_lut (.I0(encoder1_position[4]), .I1(displacement[4]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[4]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i5_3_lut (.I0(encoder0_position[4]), .I1(motor_state_23__N_106[4]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1122_3_lut_3_lut (.I0(n1667), .I1(n6016), .I2(n1651), 
            .I3(GND_net), .O(n1762));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1122_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_71_i6_4_lut (.I0(encoder1_position[5]), .I1(displacement[5]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[5]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13517_3_lut (.I0(\half_duty[0] [4]), .I1(half_duty_new[4]), 
            .I2(n1170), .I3(GND_net), .O(n18256));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_70_i6_3_lut (.I0(encoder0_position[5]), .I1(motor_state_23__N_106[5]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1124_3_lut_3_lut (.I0(n1667), .I1(n6018), .I2(n1653), 
            .I3(GND_net), .O(n1764));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1124_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13516_3_lut (.I0(\half_duty[0] [3]), .I1(half_duty_new[3]), 
            .I2(n1170), .I3(GND_net), .O(n18255));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i7_4_lut (.I0(encoder1_position[6]), .I1(displacement[6]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[6]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i7_3_lut (.I0(encoder0_position[6]), .I1(motor_state_23__N_106[6]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1118_3_lut_3_lut (.I0(n1667), .I1(n6012), .I2(n1647), 
            .I3(GND_net), .O(n1758));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1118_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1117_3_lut_3_lut (.I0(n1667), .I1(n6011), .I2(n1646), 
            .I3(GND_net), .O(n1757));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1117_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1125_3_lut_3_lut (.I0(n1667), .I1(n6019), .I2(n1054_adj_4733), 
            .I3(GND_net), .O(n1765));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1125_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4918));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1120_3_lut_3_lut (.I0(n1667), .I1(n6014), .I2(n1649), 
            .I3(GND_net), .O(n1760));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1120_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_71_i8_4_lut (.I0(encoder1_position[7]), .I1(displacement[7]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[7]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i8_3_lut (.I0(encoder0_position[7]), .I1(motor_state_23__N_106[7]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1119_3_lut_3_lut (.I0(n1667), .I1(n6013), .I2(n1648), 
            .I3(GND_net), .O(n1759));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1119_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_71_i9_4_lut (.I0(encoder1_position[8]), .I1(displacement[8]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[8]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i9_3_lut (.I0(encoder0_position[8]), .I1(motor_state_23__N_106[8]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1116_3_lut_3_lut (.I0(n1667), .I1(n6010), .I2(n1645), 
            .I3(GND_net), .O(n1756));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1116_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1115_3_lut_3_lut (.I0(n1667), .I1(n6009), .I2(n1644), 
            .I3(GND_net), .O(n1755));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1115_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1606_3_lut (.I0(n2357_adj_4941), .I1(n2424), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2456_adj_4877));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i10_4_lut (.I0(encoder1_position[9]), .I1(displacement[9]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[9]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 div_46_i1114_3_lut_3_lut (.I0(n1667), .I1(n6008), .I2(n1643), 
            .I3(GND_net), .O(n1754));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1114_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13515_3_lut (.I0(\half_duty[0] [2]), .I1(half_duty_new[2]), 
            .I2(n1170), .I3(GND_net), .O(n18254));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13515_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_70_i10_3_lut (.I0(encoder0_position[9]), .I1(motor_state_23__N_106[9]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1121_3_lut_3_lut (.I0(n1667), .I1(n6015), .I2(n1650), 
            .I3(GND_net), .O(n1761));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1121_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_71_i11_4_lut (.I0(encoder1_position[10]), .I1(displacement[10]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[10]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i11_3_lut (.I0(encoder0_position[10]), .I1(motor_state_23__N_106[10]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1198_3_lut_3_lut (.I0(n1778), .I1(n6033), .I2(n1765), 
            .I3(GND_net), .O(n1873));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1198_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1589_3_lut (.I0(n2340), .I1(n2407), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2439));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13514_3_lut (.I0(\half_duty[0] [1]), .I1(half_duty_new[1]), 
            .I2(n1170), .I3(GND_net), .O(n18253));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i13514_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_71_i12_4_lut (.I0(encoder1_position[11]), .I1(displacement[11]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[11]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i12_3_lut (.I0(encoder0_position[11]), .I1(motor_state_23__N_106[11]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1187_3_lut_3_lut (.I0(n1778), .I1(n6022), .I2(n1754), 
            .I3(GND_net), .O(n1862));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1187_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12_3_lut_adj_1859 (.I0(bit_ctr[20]), .I1(n40715), .I2(n4483), 
            .I3(GND_net), .O(n33651));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1859.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1860 (.I0(bit_ctr[19]), .I1(n40714), .I2(n4483), 
            .I3(GND_net), .O(n33649));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1860.LUT_INIT = 16'hacac;
    SB_LUT4 mux_71_i13_4_lut (.I0(encoder1_position[12]), .I1(displacement[12]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[12]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i13_3_lut (.I0(encoder0_position[12]), .I1(motor_state_23__N_106[12]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1197_3_lut_3_lut (.I0(n1778), .I1(n6032), .I2(n1764), 
            .I3(GND_net), .O(n1872));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1197_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_71_i14_4_lut (.I0(encoder1_position[13]), .I1(displacement[13]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[13]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12_3_lut_adj_1861 (.I0(bit_ctr[30]), .I1(n40725), .I2(n4483), 
            .I3(GND_net), .O(n33671));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1861.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1862 (.I0(n2439), .I1(n2438), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_5328));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i1_2_lut_adj_1862.LUT_INIT = 16'heeee;
    SB_LUT4 mux_70_i14_3_lut (.I0(encoder0_position[13]), .I1(motor_state_23__N_106[13]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1195_3_lut_3_lut (.I0(n1778), .I1(n6030), .I2(n1762), 
            .I3(GND_net), .O(n1870));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1195_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1196_3_lut_3_lut (.I0(n1778), .I1(n6031), .I2(n1763), 
            .I3(GND_net), .O(n1871));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1196_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1192_3_lut_3_lut (.I0(n1778), .I1(n6027), .I2(n1759), 
            .I3(GND_net), .O(n1867));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1192_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12_3_lut_adj_1863 (.I0(bit_ctr[29]), .I1(n40724), .I2(n4483), 
            .I3(GND_net), .O(n33669));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1863.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1864 (.I0(bit_ctr[28]), .I1(n40723), .I2(n4483), 
            .I3(GND_net), .O(n33667));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1864.LUT_INIT = 16'hacac;
    SB_LUT4 mux_71_i15_4_lut (.I0(encoder1_position[14]), .I1(displacement[14]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[14]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_adj_1865 (.I0(n2456_adj_4877), .I1(n2458_adj_4875), 
            .I2(GND_net), .I3(GND_net), .O(n38425));
    defparam i1_2_lut_adj_1865.LUT_INIT = 16'heeee;
    SB_LUT4 mux_70_i15_3_lut (.I0(encoder0_position[14]), .I1(motor_state_23__N_106[14]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1191_3_lut_3_lut (.I0(n1778), .I1(n6026), .I2(n1758), 
            .I3(GND_net), .O(n1866));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1191_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12898_3_lut (.I0(n17385), .I1(r_Bit_Index_adj_5402[0]), .I2(n17256), 
            .I3(GND_net), .O(n17637));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12898_3_lut.LUT_INIT = 16'h1414;
    SB_LUT4 mux_71_i16_4_lut (.I0(encoder1_position[15]), .I1(displacement[15]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[15]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12_3_lut_adj_1866 (.I0(bit_ctr[14]), .I1(n40704), .I2(n4483), 
            .I3(GND_net), .O(n33623));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1866.LUT_INIT = 16'hacac;
    SB_LUT4 mux_70_i16_3_lut (.I0(encoder0_position[15]), .I1(motor_state_23__N_106[15]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1194_3_lut_3_lut (.I0(n1778), .I1(n6029), .I2(n1761), 
            .I3(GND_net), .O(n1869));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1194_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12801_4_lut (.I0(n17376), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(n17250), .O(n17540));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12801_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 mux_71_i17_4_lut (.I0(encoder1_position[16]), .I1(displacement[16]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[16]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i17_3_lut (.I0(encoder0_position[16]), .I1(motor_state_23__N_106[16]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_3_lut_adj_1867 (.I0(bit_ctr[31]), .I1(n40726), .I2(n4483), 
            .I3(GND_net), .O(n33673));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1867.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1199_3_lut_3_lut (.I0(n1778), .I1(n6034), .I2(n1055_adj_4734), 
            .I3(GND_net), .O(n1874));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1199_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1193_3_lut_3_lut (.I0(n1778), .I1(n6028), .I2(n1760), 
            .I3(GND_net), .O(n1868));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1193_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_71_i18_4_lut (.I0(encoder1_position[17]), .I1(displacement[17]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[17]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_adj_1868 (.I0(n2454_adj_4879), .I1(n38425), .I2(n2455_adj_4878), 
            .I3(n2457_adj_4876), .O(n36076));
    defparam i1_4_lut_adj_1868.LUT_INIT = 16'ha080;
    SB_LUT4 mux_70_i18_3_lut (.I0(encoder0_position[17]), .I1(motor_state_23__N_106[17]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1190_3_lut_3_lut (.I0(n1778), .I1(n6025), .I2(n1757), 
            .I3(GND_net), .O(n1865));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1190_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1189_3_lut_3_lut (.I0(n1778), .I1(n6024), .I2(n1756), 
            .I3(GND_net), .O(n1864));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1189_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1188_3_lut_3_lut (.I0(n1778), .I1(n6023), .I2(n1755), 
            .I3(GND_net), .O(n1863));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1188_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_71_i19_4_lut (.I0(encoder1_position[18]), .I1(displacement[18]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[18]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i19_3_lut (.I0(encoder0_position[18]), .I1(motor_state_23__N_106[18]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_4_lut_adj_1869 (.I0(n2449_adj_4885), .I1(n2450_adj_4884), 
            .I2(n2451_adj_4883), .I3(n18_adj_5328), .O(n30_adj_5324));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i13_4_lut_adj_1869.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_71_i20_4_lut (.I0(encoder1_position[19]), .I1(displacement[19]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[19]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i20_3_lut (.I0(encoder0_position[19]), .I1(motor_state_23__N_106[19]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1266_3_lut_3_lut (.I0(n1886), .I1(n6045), .I2(n1870), 
            .I3(GND_net), .O(n1975));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1266_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1260_3_lut_3_lut (.I0(n1886), .I1(n6039), .I2(n1864), 
            .I3(GND_net), .O(n1969));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1260_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_71_i21_4_lut (.I0(encoder1_position[20]), .I1(displacement[20]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[20]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i12_3_lut_adj_1870 (.I0(byte_transmit_counter[1]), .I1(n40746), 
            .I2(n24918), .I3(GND_net), .O(n34419));   // verilog/coms.v(127[12] 295[6])
    defparam i12_3_lut_adj_1870.LUT_INIT = 16'hacac;
    SB_LUT4 mux_70_i21_3_lut (.I0(encoder0_position[20]), .I1(motor_state_23__N_106[20]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1259_3_lut_3_lut (.I0(n1886), .I1(n6038), .I2(n1863), 
            .I3(GND_net), .O(n1968));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1259_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i11_4_lut_adj_1871 (.I0(n2444), .I1(n2445), .I2(n36076), .I3(n2446), 
            .O(n28_adj_5326));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i11_4_lut_adj_1871.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1258_3_lut_3_lut (.I0(n1886), .I1(n6037), .I2(n1862), 
            .I3(GND_net), .O(n1967));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1258_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 mux_71_i22_4_lut (.I0(encoder1_position[21]), .I1(displacement[21]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[21]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i22_3_lut (.I0(encoder0_position[21]), .I1(motor_state_23__N_106[21]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1264_3_lut_3_lut (.I0(n1886), .I1(n6043), .I2(n1868), 
            .I3(GND_net), .O(n1973));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1264_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12_4_lut_adj_1872 (.I0(n2448_adj_4886), .I1(n2447_adj_4887), 
            .I2(n2453_adj_4881), .I3(n2452_adj_4882), .O(n29_adj_5325));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i12_4_lut_adj_1872.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_71_i23_4_lut (.I0(encoder1_position[22]), .I1(displacement[22]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[22]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i23_3_lut (.I0(encoder0_position[22]), .I1(motor_state_23__N_106[22]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1265_3_lut_3_lut (.I0(n1886), .I1(n6044), .I2(n1869), 
            .I3(GND_net), .O(n1974));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1265_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i4_4_lut_adj_1873 (.I0(control_mode[3]), .I1(control_mode[5]), 
            .I2(control_mode[4]), .I3(control_mode[7]), .O(n10_adj_5230));   // verilog/TinyFPGA_B.v(211[5:22])
    defparam i4_4_lut_adj_1873.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(control_mode[6]), .I1(n10_adj_5230), .I2(control_mode[2]), 
            .I3(GND_net), .O(n15942));   // verilog/TinyFPGA_B.v(211[5:22])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut (.I0(control_mode[0]), .I1(control_mode[1]), .I2(n15942), 
            .I3(GND_net), .O(n15_adj_4665));   // verilog/TinyFPGA_B.v(211[5:22])
    defparam i2_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 mux_71_i24_4_lut (.I0(encoder1_position[23]), .I1(displacement[23]), 
            .I2(n15_adj_4665), .I3(n15), .O(motor_state_23__N_106[23]));   // verilog/TinyFPGA_B.v(211[5] 214[10])
    defparam mux_71_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 mux_70_i24_3_lut (.I0(encoder0_position[23]), .I1(motor_state_23__N_106[23]), 
            .I2(n15_adj_4673), .I3(GND_net), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(210[5] 214[10])
    defparam mux_70_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1270_3_lut_3_lut (.I0(n1886), .I1(n6049), .I2(n1874), 
            .I3(GND_net), .O(n1979));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1270_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i10_4_lut_adj_1874 (.I0(n2440), .I1(n2442), .I2(n2441), .I3(n2443), 
            .O(n27_adj_5327));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i10_4_lut_adj_1874.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1269_3_lut_3_lut (.I0(n1886), .I1(n6048), .I2(n1873), 
            .I3(GND_net), .O(n1978));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1269_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i16_4_lut_adj_1875 (.I0(n27_adj_5327), .I1(n29_adj_5325), .I2(n28_adj_5326), 
            .I3(n30_adj_5324), .O(n2471_adj_4874));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i16_4_lut_adj_1875.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1267_3_lut_3_lut (.I0(n1886), .I1(n6046), .I2(n1871), 
            .I3(GND_net), .O(n1976));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1267_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1591_3_lut (.I0(n2342), .I1(n2409), .I2(n2372_adj_4939), 
            .I3(GND_net), .O(n2441));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1268_3_lut_3_lut (.I0(n1886), .I1(n6047), .I2(n1872), 
            .I3(GND_net), .O(n1977));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1268_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1658_3_lut (.I0(n2441), .I1(n2508), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2540_adj_4870));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12798_4_lut (.I0(n17376), .I1(r_Bit_Index[2]), .I2(n4698), 
            .I3(n17250), .O(n17537));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12798_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 rem_4_i1657_3_lut (.I0(n2440), .I1(n2507), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2539_adj_4871));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1656_3_lut (.I0(n2439), .I1(n2506), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2538_adj_4872));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4729));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4728));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4727));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4726));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4725));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1271_3_lut_3_lut (.I0(n1886), .I1(n6050), .I2(n1056_adj_4735), 
            .I3(GND_net), .O(n1980));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1271_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1263_3_lut_3_lut (.I0(n1886), .I1(n6042), .I2(n1867), 
            .I3(GND_net), .O(n1972));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1263_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1262_3_lut_3_lut (.I0(n1886), .I1(n6041), .I2(n1866), 
            .I3(GND_net), .O(n1971));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1262_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1261_3_lut_3_lut (.I0(n1886), .I1(n6040), .I2(n1865), 
            .I3(GND_net), .O(n1970));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1261_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1340_3_lut_3_lut (.I0(n1991), .I1(n6066), .I2(n1980), 
            .I3(GND_net), .O(n2082));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1340_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12_3_lut_adj_1876 (.I0(n40744), .I1(byte_transmit_counter[3]), 
            .I2(n24918), .I3(GND_net), .O(n34315));   // verilog/coms.v(127[12] 295[6])
    defparam i12_3_lut_adj_1876.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4724));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1332_3_lut_3_lut (.I0(n1991), .I1(n6058), .I2(n1972), 
            .I3(GND_net), .O(n2074));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1332_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12_3_lut_adj_1877 (.I0(byte_transmit_counter[2]), .I1(n40747), 
            .I2(n24918), .I3(GND_net), .O(n34421));   // verilog/coms.v(127[12] 295[6])
    defparam i12_3_lut_adj_1877.LUT_INIT = 16'hacac;
    SB_LUT4 i10_4_lut_adj_1878 (.I0(n2538_adj_4872), .I1(n2539_adj_4871), 
            .I2(n2537_adj_4873), .I3(n2540_adj_4870), .O(n28_adj_5322));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i10_4_lut_adj_1878.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1879 (.I0(n2556), .I1(n2558_adj_4856), .I2(GND_net), 
            .I3(GND_net), .O(n38205));
    defparam i1_2_lut_adj_1879.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1880 (.I0(n2554), .I1(n38205), .I2(n2555), .I3(n2557), 
            .O(n36012));
    defparam i1_4_lut_adj_1880.LUT_INIT = 16'ha080;
    SB_LUT4 div_46_i1330_3_lut_3_lut (.I0(n1991), .I1(n6056), .I2(n1970), 
            .I3(GND_net), .O(n2072));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1330_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1329_3_lut_3_lut (.I0(n1991), .I1(n6055), .I2(n1969), 
            .I3(GND_net), .O(n2071));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1329_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i14_3_lut (.I0(n2548_adj_4862), .I1(n28_adj_5322), .I2(n2547_adj_4863), 
            .I3(GND_net), .O(n32_adj_5318));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i14_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 displacement_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4723));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1328_3_lut_3_lut (.I0(n1991), .I1(n6054), .I2(n1968), 
            .I3(GND_net), .O(n2070));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1328_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12_3_lut_adj_1881 (.I0(n40742), .I1(byte_transmit_counter[5]), 
            .I2(n24918), .I3(GND_net), .O(n34225));   // verilog/coms.v(127[12] 295[6])
    defparam i12_3_lut_adj_1881.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1327_3_lut_3_lut (.I0(n1991), .I1(n6053), .I2(n1967), 
            .I3(GND_net), .O(n2069));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1327_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12_4_lut_adj_1882 (.I0(n36012), .I1(n2546_adj_4864), .I2(n2545_adj_4865), 
            .I3(n2549_adj_4861), .O(n30_adj_5320));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i12_4_lut_adj_1882.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_3_lut_adj_1883 (.I0(n40743), .I1(byte_transmit_counter[4]), 
            .I2(n24918), .I3(GND_net), .O(n34267));   // verilog/coms.v(127[12] 295[6])
    defparam i12_3_lut_adj_1883.LUT_INIT = 16'hcaca;
    SB_LUT4 i13_4_lut_adj_1884 (.I0(n2552_adj_4858), .I1(n2551_adj_4859), 
            .I2(n2550_adj_4860), .I3(n2553_adj_4857), .O(n31_adj_5319));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i13_4_lut_adj_1884.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_3_lut_adj_1885 (.I0(n40740), .I1(byte_transmit_counter[7]), 
            .I2(n24918), .I3(GND_net), .O(n34167));   // verilog/coms.v(127[12] 295[6])
    defparam i12_3_lut_adj_1885.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1886 (.I0(n2541_adj_4869), .I1(n2543_adj_4867), 
            .I2(n2542_adj_4868), .I3(n2544_adj_4866), .O(n29_adj_5321));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i11_4_lut_adj_1886.LUT_INIT = 16'hfffe;
    SB_LUT4 displacement_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4722));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4721));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i17_4_lut_adj_1887 (.I0(n29_adj_5321), .I1(n31_adj_5319), .I2(n30_adj_5320), 
            .I3(n32_adj_5318), .O(n2570));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i17_4_lut_adj_1887.LUT_INIT = 16'hfffe;
    SB_LUT4 displacement_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4720));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1660_3_lut (.I0(n2443), .I1(n2510), .I2(n2471_adj_4874), 
            .I3(GND_net), .O(n2542_adj_4868));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1336_3_lut_3_lut (.I0(n1991), .I1(n6062), .I2(n1976), 
            .I3(GND_net), .O(n2078));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1336_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i1727_3_lut (.I0(n2542_adj_4868), .I1(n2609), .I2(n2570), 
            .I3(GND_net), .O(n2641));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1727_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1725_3_lut (.I0(n2540_adj_4870), .I1(n2607), .I2(n2570), 
            .I3(GND_net), .O(n2639));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1725_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1726_3_lut (.I0(n2541_adj_4869), .I1(n2608), .I2(n2570), 
            .I3(GND_net), .O(n2640));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1726_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i1724_3_lut (.I0(n2539_adj_4871), .I1(n2606), .I2(n2570), 
            .I3(GND_net), .O(n2638_adj_4845));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1724_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1334_3_lut_3_lut (.I0(n1991), .I1(n6060), .I2(n1974), 
            .I3(GND_net), .O(n2076));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1334_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i11_4_lut_adj_1888 (.I0(n2638_adj_4845), .I1(n2640), .I2(n2639), 
            .I3(n2641), .O(n30_adj_5266));
    defparam i11_4_lut_adj_1888.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1889 (.I0(n2656), .I1(n2658), .I2(GND_net), .I3(GND_net), 
            .O(n38429));
    defparam i1_2_lut_adj_1889.LUT_INIT = 16'heeee;
    SB_LUT4 displacement_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4719));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4718));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4717));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1890 (.I0(n2654), .I1(n38429), .I2(n2655), .I3(n2657), 
            .O(n36089));
    defparam i1_4_lut_adj_1890.LUT_INIT = 16'ha080;
    SB_LUT4 i15_4_lut_adj_1891 (.I0(n2653), .I1(n30_adj_5266), .I2(n2637_adj_4846), 
            .I3(n2636_adj_4847), .O(n34_adj_5262));
    defparam i15_4_lut_adj_1891.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1892 (.I0(n2645), .I1(n2651), .I2(n2646), .I3(n2649), 
            .O(n32_adj_5264));
    defparam i13_4_lut_adj_1892.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1893 (.I0(n2650), .I1(n2652), .I2(n2648), .I3(n2647), 
            .O(n33_adj_5263));
    defparam i14_4_lut_adj_1893.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1894 (.I0(n2642_adj_4844), .I1(n36089), .I2(n2643_adj_4843), 
            .I3(n2644), .O(n31_adj_5265));
    defparam i12_4_lut_adj_1894.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1335_3_lut_3_lut (.I0(n1991), .I1(n6061), .I2(n1975), 
            .I3(GND_net), .O(n2077));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1335_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1338_3_lut_3_lut (.I0(n1991), .I1(n6064), .I2(n1978), 
            .I3(GND_net), .O(n2080));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1338_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i18_4_lut_adj_1895 (.I0(n31_adj_5265), .I1(n33_adj_5263), .I2(n32_adj_5264), 
            .I3(n34_adj_5262), .O(n2669));
    defparam i18_4_lut_adj_1895.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i10_3_lut (.I0(communication_counter[9]), .I1(n24_adj_4785), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2658));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4716));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1811_3_lut (.I0(n2658), .I1(n2725), .I2(n2669), .I3(GND_net), 
            .O(n2757));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 displacement_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4664));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1810_3_lut (.I0(n2657), .I1(n2724_adj_4823), .I2(n2669), 
            .I3(GND_net), .O(n2756));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1810_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut_adj_1896 (.I0(n2756), .I1(n2757), .I2(n2758), .I3(GND_net), 
            .O(n36026));
    defparam i1_3_lut_adj_1896.LUT_INIT = 16'hfefe;
    SB_LUT4 displacement_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4676));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4677));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4681));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4682));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4683));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i14_4_lut_adj_1897 (.I0(n2746), .I1(n2745), .I2(n2753), .I3(n2747), 
            .O(n34_adj_5238));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i14_4_lut_adj_1897.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1339_3_lut_3_lut (.I0(n1991), .I1(n6065), .I2(n1979), 
            .I3(GND_net), .O(n2081));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1339_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_mux_3_i1_3_lut (.I0(communication_counter[0]), .I1(n33), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3360));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i1_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i5_4_lut_adj_1898 (.I0(n2743), .I1(n2754), .I2(n36026), .I3(n2755), 
            .O(n25_adj_5241));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i5_4_lut_adj_1898.LUT_INIT = 16'heaaa;
    SB_LUT4 rem_4_mux_3_i2_3_lut (.I0(communication_counter[1]), .I1(n32), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n3458));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i2_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i12_3_lut_adj_1899 (.I0(bit_ctr[9]), .I1(n40698), .I2(n4483), 
            .I3(GND_net), .O(n33589));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1899.LUT_INIT = 16'hacac;
    SB_LUT4 i12_4_lut_adj_1900 (.I0(n2739), .I1(n2741), .I2(n2740), .I3(n2742), 
            .O(n32_adj_5239));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i12_4_lut_adj_1900.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_3_lut (.I0(blink), .I1(color[12]), .I2(n25734), .I3(GND_net), 
            .O(n32167));
    defparam i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_2_lut (.I0(color_23__N_164[4]), .I1(color_23__N_164[1]), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_4744));   // verilog/TinyFPGA_B.v(54[6:36])
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1901 (.I0(color_23__N_164[5]), .I1(color_23__N_164[6]), 
            .I2(color_23__N_164[3]), .I3(color_23__N_164[0]), .O(n13_adj_5341));   // verilog/TinyFPGA_B.v(54[6:36])
    defparam i1_4_lut_adj_1901.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1902 (.I0(color_23__N_164[7]), .I1(n13_adj_5341), 
            .I2(n12_adj_4744), .I3(color_23__N_164[2]), .O(n25734));   // verilog/TinyFPGA_B.v(54[6:36])
    defparam i1_4_lut_adj_1902.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1903 (.I0(n2736), .I1(n2737), .I2(n2735), .I3(n2738), 
            .O(n31_adj_5240));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i11_4_lut_adj_1903.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1904 (.I0(color_23__N_164[2]), .I1(blink), .I2(GND_net), 
            .I3(GND_net), .O(n37725));
    defparam i1_2_lut_adj_1904.LUT_INIT = 16'h4444;
    SB_LUT4 i1_4_lut_adj_1905 (.I0(color_23__N_164[7]), .I1(n13_adj_5341), 
            .I2(n12_adj_4744), .I3(n37725), .O(n25736));
    defparam i1_4_lut_adj_1905.LUT_INIT = 16'h0100;
    SB_LUT4 i1_3_lut_adj_1906 (.I0(color[11]), .I1(n25736), .I2(n25734), 
            .I3(GND_net), .O(n18223));
    defparam i1_3_lut_adj_1906.LUT_INIT = 16'hecec;
    SB_LUT4 div_46_i1337_3_lut_3_lut (.I0(n1991), .I1(n6063), .I2(n1977), 
            .I3(GND_net), .O(n2079));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1337_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12764_4_lut (.I0(n17505), .I1(r_Clock_Count_adj_5401[2]), .I2(n319), 
            .I3(r_SM_Main_adj_5400[2]), .O(n17503));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12764_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 i15_4_lut_adj_1907 (.I0(n2751), .I1(n2748), .I2(n2750), .I3(n2749), 
            .O(n35_adj_5237));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i15_4_lut_adj_1907.LUT_INIT = 16'hfffe;
    SB_LUT4 div_46_i1341_3_lut_3_lut (.I0(n1991), .I1(n6067), .I2(n1057_adj_4736), 
            .I3(GND_net), .O(n2083));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1341_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i17_4_lut_adj_1908 (.I0(n25_adj_5241), .I1(n34_adj_5238), .I2(n2752), 
            .I3(n2744), .O(n37_adj_5236));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i17_4_lut_adj_1908.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1909 (.I0(n37_adj_5236), .I1(n35_adj_5237), .I2(n31_adj_5240), 
            .I3(n32_adj_5239), .O(n2768));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i19_4_lut_adj_1909.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_mux_3_i9_3_lut (.I0(communication_counter[8]), .I1(n25_adj_4784), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2758));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1333_3_lut_3_lut (.I0(n1991), .I1(n6059), .I2(n1973), 
            .I3(GND_net), .O(n2075));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1333_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12767_4_lut (.I0(n17505), .I1(r_Clock_Count_adj_5401[1]), .I2(n320), 
            .I3(r_SM_Main_adj_5400[2]), .O(n17506));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12767_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i1_1_lut (.I0(communication_counter[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n33_adj_5306));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1331_3_lut_3_lut (.I0(n1991), .I1(n6057), .I2(n1971), 
            .I3(GND_net), .O(n2073));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1331_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_mux_3_i8_3_lut (.I0(communication_counter[7]), .I1(n26_adj_4783), 
            .I2(communication_counter[31]), .I3(GND_net), .O(n2858));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i2_1_lut (.I0(communication_counter[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_5305));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 displacement_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4689));   // verilog/TinyFPGA_B.v(232[21:79])
    defparam displacement_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i3_1_lut (.I0(communication_counter[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_5304));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i4_1_lut (.I0(communication_counter[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_5303));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36734_1_lut (.I0(n38575), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43581));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i36734_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2287_rep_5_3_lut (.I0(n3358), .I1(n10249), .I2(n3362), 
            .I3(GND_net), .O(n38575));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2287_rep_5_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i5_1_lut (.I0(communication_counter[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_5302));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1879_3_lut (.I0(n2758), .I1(n2825), .I2(n2768), .I3(GND_net), 
            .O(n2857));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i6_1_lut (.I0(communication_counter[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_5301));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i1878_3_lut (.I0(n2757), .I1(n2824), .I2(n2768), .I3(GND_net), 
            .O(n2856));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i1878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i7_1_lut (.I0(communication_counter[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_5300));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i8_1_lut (.I0(communication_counter[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_5299));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36731_1_lut (.I0(n3456), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43578));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i36731_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2286_3_lut (.I0(n3357), .I1(n10248), .I2(n3362), .I3(GND_net), 
            .O(n3456));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2286_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i9_1_lut (.I0(communication_counter[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5298));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_3_lut_adj_1910 (.I0(n2856), .I1(n2857), .I2(n2858), .I3(GND_net), 
            .O(n36097));
    defparam i1_3_lut_adj_1910.LUT_INIT = 16'hfefe;
    SB_LUT4 i5_4_lut_adj_1911 (.I0(n2842), .I1(n2854), .I2(n36097), .I3(n2855), 
            .O(n26_adj_5260));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i5_4_lut_adj_1911.LUT_INIT = 16'heaaa;
    SB_LUT4 i12_4_lut_adj_1912 (.I0(n2836), .I1(n2838), .I2(n2837), .I3(n2839), 
            .O(n33_adj_5259));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i12_4_lut_adj_1912.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i10_1_lut (.I0(communication_counter[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5297));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i11_1_lut (.I0(communication_counter[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5296));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i12_1_lut (.I0(communication_counter[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5295));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i13_1_lut (.I0(communication_counter[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5294));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36728_1_lut (.I0(n3455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43575));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i36728_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2285_3_lut (.I0(n3356), .I1(n10247), .I2(n3362), .I3(GND_net), 
            .O(n3455));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2285_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i1_2_lut_adj_1913 (.I0(n2835), .I1(n2834), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_5261));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i1_2_lut_adj_1913.LUT_INIT = 16'heeee;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i14_1_lut (.I0(communication_counter[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5293));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i15_1_lut (.I0(communication_counter[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5292));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i16_1_lut (.I0(communication_counter[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5291));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36725_1_lut (.I0(n3454), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43572));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i36725_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2284_3_lut (.I0(n3355), .I1(n10246), .I2(n3362), .I3(GND_net), 
            .O(n3454));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2284_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i17_4_lut_adj_1914 (.I0(n33_adj_5259), .I1(n2840), .I2(n26_adj_5260), 
            .I3(n2841), .O(n38_adj_5255));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i17_4_lut_adj_1914.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i17_1_lut (.I0(communication_counter[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5290));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i18_1_lut (.I0(communication_counter[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5289));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i19_1_lut (.I0(communication_counter[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5288));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36722_1_lut (.I0(n3453), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43569));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i36722_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_i2283_3_lut (.I0(n3354), .I1(n10245), .I2(n3362), .I3(GND_net), 
            .O(n3453));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2283_3_lut.LUT_INIT = 16'h3535;
    SB_LUT4 i15_4_lut_adj_1915 (.I0(n2851), .I1(n2846), .I2(n2847), .I3(n2845), 
            .O(n36_adj_5257));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i15_4_lut_adj_1915.LUT_INIT = 16'hfffe;
    SB_LUT4 rem_4_i2206_3_lut (.I0(n3245), .I1(n3312), .I2(n3263), .I3(GND_net), 
            .O(n3344));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2205_3_lut (.I0(n3244), .I1(n3311), .I2(n3263), .I3(GND_net), 
            .O(n3343));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i16_4_lut_adj_1916 (.I0(n2850), .I1(n2853), .I2(n2849), .I3(n22_adj_5261), 
            .O(n37_adj_5256));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i16_4_lut_adj_1916.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1917 (.I0(n3246), .I1(n3343), .I2(n3313), .I3(n3263), 
            .O(n38049));
    defparam i1_4_lut_adj_1917.LUT_INIT = 16'hfcee;
    SB_LUT4 rem_4_i2208_3_lut (.I0(n3247), .I1(n3314), .I2(n3263), .I3(GND_net), 
            .O(n3346));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 rem_4_i2213_3_lut (.I0(n3252), .I1(n3319), .I2(n3263), .I3(GND_net), 
            .O(n3351));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2213_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1918 (.I0(n3249), .I1(n3351), .I2(n3316), .I3(n3263), 
            .O(n38099));
    defparam i1_4_lut_adj_1918.LUT_INIT = 16'hfcee;
    SB_LUT4 div_46_i1405_3_lut_3_lut (.I0(n2093), .I1(n6081), .I2(n2080), 
            .I3(GND_net), .O(n2179));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1405_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1406_3_lut_3_lut (.I0(n2093), .I1(n6082), .I2(n2081), 
            .I3(GND_net), .O(n2180));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1406_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1409_3_lut_3_lut (.I0(n2093), .I1(n6085), .I2(n1058_adj_4737), 
            .I3(GND_net), .O(n2183));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1409_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_4_lut_adj_1919 (.I0(n38099), .I1(n3251), .I2(n3318), .I3(n3263), 
            .O(n38101));
    defparam i1_4_lut_adj_1919.LUT_INIT = 16'hfaee;
    SB_LUT4 i1_4_lut_adj_1920 (.I0(n3242), .I1(n38101), .I2(n3309), .I3(n3263), 
            .O(n38103));
    defparam i1_4_lut_adj_1920.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1921 (.I0(n3240), .I1(n38103), .I2(n3307), .I3(n3263), 
            .O(n38105));
    defparam i1_4_lut_adj_1921.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1922 (.I0(n3239), .I1(n38105), .I2(n3306), .I3(n3263), 
            .O(n38107));
    defparam i1_4_lut_adj_1922.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_2_lut_adj_1923 (.I0(n3356), .I1(n3358), .I2(GND_net), .I3(GND_net), 
            .O(n38401));
    defparam i1_2_lut_adj_1923.LUT_INIT = 16'heeee;
    SB_LUT4 i14_4_lut_adj_1924 (.I0(n2843), .I1(n2844), .I2(n2852), .I3(n2848), 
            .O(n35_adj_5258));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i14_4_lut_adj_1924.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1925 (.I0(n3253), .I1(n3344), .I2(n3320), .I3(n3263), 
            .O(n38047));
    defparam i1_4_lut_adj_1925.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1926 (.I0(n38049), .I1(n3243), .I2(n3310), .I3(n3263), 
            .O(n38051));
    defparam i1_4_lut_adj_1926.LUT_INIT = 16'hfaee;
    SB_LUT4 div_46_i1397_3_lut_3_lut (.I0(n2093), .I1(n6073), .I2(n2072), 
            .I3(GND_net), .O(n2171));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1397_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1396_3_lut_3_lut (.I0(n2093), .I1(n6072), .I2(n2071), 
            .I3(GND_net), .O(n2170));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1396_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_i2202_3_lut (.I0(n3241), .I1(n3308), .I2(n3263), .I3(GND_net), 
            .O(n3340));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1927 (.I0(n3354), .I1(n38401), .I2(n3355), .I3(n3357), 
            .O(n36058));
    defparam i1_4_lut_adj_1927.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1928 (.I0(n36058), .I1(n3340), .I2(n38051), .I3(n38047), 
            .O(n38057));
    defparam i1_4_lut_adj_1928.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1929 (.I0(n3237), .I1(n38057), .I2(n3304), .I3(n3263), 
            .O(n38059));
    defparam i1_4_lut_adj_1929.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1930 (.I0(n3236), .I1(n38107), .I2(n3303), .I3(n3263), 
            .O(n38109));
    defparam i1_4_lut_adj_1930.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1931 (.I0(n3353), .I1(n3250), .I2(n3317), .I3(n3263), 
            .O(n38137));
    defparam i1_4_lut_adj_1931.LUT_INIT = 16'hfaee;
    SB_LUT4 i12771_4_lut (.I0(n17385), .I1(r_Bit_Index_adj_5402[2]), .I2(n4720), 
            .I3(n17256), .O(n17510));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12771_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 i3_4_lut_adj_1932 (.I0(n3248), .I1(n3346), .I2(n3315), .I3(n3263), 
            .O(n28_adj_5339));
    defparam i3_4_lut_adj_1932.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1933 (.I0(n38109), .I1(n3235), .I2(n3302), .I3(n3263), 
            .O(n46_adj_5337));
    defparam i1_4_lut_adj_1933.LUT_INIT = 16'hfaee;
    SB_LUT4 i1_4_lut_adj_1934 (.I0(n38059), .I1(n3233), .I2(n3300), .I3(n3263), 
            .O(n47_adj_5331));
    defparam i1_4_lut_adj_1934.LUT_INIT = 16'hfaee;
    SB_LUT4 rem_4_i2199_3_lut (.I0(n3238), .I1(n3305), .I2(n3263), .I3(GND_net), 
            .O(n3337));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20_4_lut_adj_1935 (.I0(n35_adj_5258), .I1(n37_adj_5256), .I2(n36_adj_5257), 
            .I3(n38_adj_5255), .O(n2867));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i20_4_lut_adj_1935.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1936 (.I0(n3234), .I1(n3337), .I2(n3301), .I3(n3263), 
            .O(n37783));
    defparam i1_4_lut_adj_1936.LUT_INIT = 16'hfcee;
    SB_LUT4 rem_4_i2192_3_lut (.I0(n3231), .I1(n3298), .I2(n3263), .I3(GND_net), 
            .O(n3330));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i2192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1937 (.I0(n47_adj_5331), .I1(n46_adj_5337), .I2(n28_adj_5339), 
            .I3(n38137), .O(n38143));
    defparam i1_4_lut_adj_1937.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1938 (.I0(n3232), .I1(n37783), .I2(n3299), .I3(n3263), 
            .O(n37785));
    defparam i1_4_lut_adj_1938.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1939 (.I0(n38464), .I1(n37785), .I2(n38143), 
            .I3(n3330), .O(n3362));
    defparam i1_4_lut_adj_1939.LUT_INIT = 16'hfffe;
    SB_LUT4 i36721_2_lut (.I0(n3362), .I1(n10244), .I2(GND_net), .I3(GND_net), 
            .O(n3452));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i36721_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 div_46_i1395_3_lut_3_lut (.I0(n2093), .I1(n6071), .I2(n2070), 
            .I3(GND_net), .O(n2169));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1395_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i20_1_lut (.I0(communication_counter[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5287));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i21_1_lut (.I0(communication_counter[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5286));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i22_1_lut (.I0(communication_counter[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5285));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i23_1_lut (.I0(communication_counter[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5284));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i24_1_lut (.I0(communication_counter[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_5283));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1398_3_lut_3_lut (.I0(n2093), .I1(n6074), .I2(n2073), 
            .I3(GND_net), .O(n2172));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1398_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i25_1_lut (.I0(communication_counter[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_5282));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1394_3_lut_3_lut (.I0(n2093), .I1(n6070), .I2(n2069), 
            .I3(GND_net), .O(n2168));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1394_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i26_1_lut (.I0(communication_counter[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_5281));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i27_1_lut (.I0(communication_counter[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_5280));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_unary_minus_4_inv_0_i1_1_lut (.I0(gearBoxRatio[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4911));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i28_1_lut (.I0(communication_counter[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_5279));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i29_1_lut (.I0(communication_counter[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_5278));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i30_1_lut (.I0(communication_counter[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_5277));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i31_1_lut (.I0(communication_counter[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_5276));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 rem_4_unary_minus_2_inv_0_i32_1_lut (.I0(communication_counter[31]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_5275));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1404_3_lut_3_lut (.I0(n2093), .I1(n6080), .I2(n2079), 
            .I3(GND_net), .O(n2178));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1404_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_unary_minus_4_inv_0_i2_1_lut (.I0(gearBoxRatio[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n24_adj_4910));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 div_46_i1408_3_lut_3_lut (.I0(n2093), .I1(n6084), .I2(n2083), 
            .I3(GND_net), .O(n2182));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1408_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1402_3_lut_3_lut (.I0(n2093), .I1(n6078), .I2(n2077), 
            .I3(GND_net), .O(n2176));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1402_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1403_3_lut_3_lut (.I0(n2093), .I1(n6079), .I2(n2078), 
            .I3(GND_net), .O(n2177));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1403_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12774_4_lut (.I0(n17385), .I1(r_Bit_Index_adj_5402[1]), .I2(r_Bit_Index_adj_5402[0]), 
            .I3(n17256), .O(n17513));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12774_4_lut.LUT_INIT = 16'h1444;
    SB_LUT4 div_46_i1400_3_lut_3_lut (.I0(n2093), .I1(n6076), .I2(n2075), 
            .I3(GND_net), .O(n2174));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1400_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13498_3_lut (.I0(setpoint[8]), .I1(n4394), .I2(n37622), .I3(GND_net), 
            .O(n18237));   // verilog/coms.v(127[12] 295[6])
    defparam i13498_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1401_3_lut_3_lut (.I0(n2093), .I1(n6077), .I2(n2076), 
            .I3(GND_net), .O(n2175));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1401_3_lut_3_lut.LUT_INIT = 16'he4e4;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(35[10] 38[2])
    coms setpoint_23__I_0 (.clk32MHz(clk32MHz), .GND_net(GND_net), .rx_data({rx_data}), 
         .\data_in_frame[20] ({\data_in_frame[20] }), .\data_in_frame[8] ({\data_in_frame[8] }), 
         .n18251(n18251), .setpoint({setpoint}), .n36556(n36556), .n18252(n18252), 
         .n18231(n18231), .n18232(n18232), .n18233(n18233), .n18234(n18234), 
         .n18235(n18235), .n18236(n18236), .n18237(n18237), .n34167(n34167), 
         .\byte_transmit_counter[7] (byte_transmit_counter[7]), .n34267(n34267), 
         .\byte_transmit_counter[4] (byte_transmit_counter[4]), .n34225(n34225), 
         .\byte_transmit_counter[5] (byte_transmit_counter[5]), .n34421(n34421), 
         .\byte_transmit_counter[2] (byte_transmit_counter[2]), .n34315(n34315), 
         .\byte_transmit_counter[3] (byte_transmit_counter[3]), .n34419(n34419), 
         .\byte_transmit_counter[1] (byte_transmit_counter[1]), .n43830(n43830), 
         .n18249(n18249), .n18250(n18250), .n18247(n18247), .n18248(n18248), 
         .n18245(n18245), .n18246(n18246), .n18243(n18243), .n18244(n18244), 
         .n18241(n18241), .n18242(n18242), .n18238(n18238), .n18239(n18239), 
         .n18240(n18240), .n18230(n18230), .n18145(n18145), .PWMLimit({PWMLimit}), 
         .n18146(n18146), .n18147(n18147), .n18148(n18148), .n18149(n18149), 
         .n18150(n18150), .n18151(n18151), .n34409(n34409), .\byte_transmit_counter[0] (byte_transmit_counter[0]), 
         .n18137(n18137), .n18138(n18138), .n18139(n18139), .n18140(n18140), 
         .n18141(n18141), .n18142(n18142), .\data_in_frame[21] ({\data_in_frame[21] }), 
         .n18155(n18155), .n18156(n18156), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .n18152(n18152), .n18153(n18153), .n18154(n18154), .n18143(n18143), 
         .n18144(n18144), .n18133(n18133), .\data_in_frame[24] ({\data_in_frame[24] }), 
         .n18134(n18134), .n18135(n18135), .n18136(n18136), .n18126(n18126), 
         .n18127(n18127), .n18128(n18128), .n18129(n18129), .n18130(n18130), 
         .n18131(n18131), .n18132(n18132), .\data_in_frame[22] ({\data_in_frame[22] }), 
         .\data_in_frame[4] ({\data_in_frame[4] }), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .\data_in_frame[12] ({\data_in_frame[12] }), .\data_in_frame[3] ({\data_in_frame[3] }), 
         .\data_in_frame[2] ({\data_in_frame[2] }), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .\data_in_frame[1] ({\data_in_frame[1] }), .\FRAME_MATCHER.state[3] (\FRAME_MATCHER.state [3]), 
         .\FRAME_MATCHER.state[1] (\FRAME_MATCHER.state [1]), .n15963(n15963), 
         .n13302(n13302), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .\data_out_frame[5] ({\data_out_frame[5] }), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .\data_out_frame[7] ({\data_out_frame[7] }), .n17934(n17934), .control_mode({control_mode}), 
         .rx_data_ready(rx_data_ready), .n17933(n17933), .n17932(n17932), 
         .n17931(n17931), .n17930(n17930), .n17929(n17929), .n17928(n17928), 
         .n17927(n17927), .n17926(n17926), .n17925(n17925), .n17924(n17924), 
         .n17923(n17923), .n17922(n17922), .n17921(n17921), .n17920(n17920), 
         .n17919(n17919), .\data_out_frame[19] ({\data_out_frame[19] }), 
         .n17918(n17918), .n17917(n17917), .n17916(n17916), .n17915(n17915), 
         .\data_in_frame[9] ({\data_in_frame[9] }), .n17914(n17914), .n17913(n17913), 
         .n17912(n17912), .n17911(n17911), .\data_out_frame[18] ({\data_out_frame[18] }), 
         .n17910(n17910), .\data_in_frame[14][1] (\data_in_frame[14] [1]), 
         .n17909(n17909), .n35644(n35644), .n17908(n17908), .\data_in_frame[10] ({\data_in_frame[10] }), 
         .n17907(n17907), .n17906(n17906), .n17905(n17905), .n40740(n40740), 
         .n34978(n34978), .n17904(n17904), .n40742(n40742), .n40743(n40743), 
         .n17903(n17903), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .n17902(n17902), .n40744(n40744), .n37132(n37132), .n16086(n16086), 
         .n17011(n17011), .n35463(n35463), .n35626(n35626), .n17901(n17901), 
         .n17900(n17900), .n40747(n40747), .n17899(n17899), .n17898(n17898), 
         .n17897(n17897), .n17896(n17896), .n17895(n17895), .\data_out_frame[16] ({\data_out_frame[16] }), 
         .n17894(n17894), .n17893(n17893), .n17892(n17892), .n17891(n17891), 
         .PIN_11_c(PIN_11_c), .n17890(n17890), .n17889(n17889), .n17888(n17888), 
         .n17887(n17887), .\data_out_frame[15] ({\data_out_frame[15] }), 
         .n17886(n17886), .n17885(n17885), .n17884(n17884), .n17883(n17883), 
         .n17882(n17882), .n17881(n17881), .n17880(n17880), .n17879(n17879), 
         .\data_out_frame[14] ({\data_out_frame[14] }), .n17878(n17878), 
         .n17877(n17877), .n17876(n17876), .n17875(n17875), .n17874(n17874), 
         .n17873(n17873), .n40746(n40746), .n17872(n17872), .n17871(n17871), 
         .\data_out_frame[13] ({\data_out_frame[13] }), .n17870(n17870), 
         .n17869(n17869), .n17868(n17868), .n17867(n17867), .n17866(n17866), 
         .n17865(n17865), .n17864(n17864), .n17863(n17863), .\data_out_frame[12] ({\data_out_frame[12] }), 
         .n17862(n17862), .n17861(n17861), .n17860(n17860), .n17859(n17859), 
         .n17858(n17858), .n17857(n17857), .n17856(n17856), .n17855(n17855), 
         .\data_out_frame[11] ({\data_out_frame[11] }), .n17854(n17854), 
         .n17853(n17853), .n17852(n17852), .n17851(n17851), .n17850(n17850), 
         .n17849(n17849), .n17848(n17848), .n17847(n17847), .\data_out_frame[10] ({\data_out_frame[10] }), 
         .n17846(n17846), .n17845(n17845), .n40745(n40745), .n17844(n17844), 
         .n17843(n17843), .n17842(n17842), .n17841(n17841), .n17840(n17840), 
         .n17839(n17839), .\data_out_frame[9] ({\data_out_frame[9] }), .n17838(n17838), 
         .n17837(n17837), .n17836(n17836), .n17835(n17835), .n17834(n17834), 
         .n17833(n17833), .n17832(n17832), .n17831(n17831), .\data_out_frame[8] ({\data_out_frame[8] }), 
         .n17830(n17830), .n17829(n17829), .n17828(n17828), .n17827(n17827), 
         .n17826(n17826), .n17825(n17825), .n17824(n17824), .n17823(n17823), 
         .n17822(n17822), .n17821(n17821), .n17820(n17820), .n17819(n17819), 
         .n17818(n17818), .n17817(n17817), .n17816(n17816), .n17815(n17815), 
         .n17814(n17814), .n17813(n17813), .n17812(n17812), .n17811(n17811), 
         .n17810(n17810), .n17809(n17809), .n17808(n17808), .n17807(n17807), 
         .n37622(n37622), .n4408(n4408), .n17806(n17806), .n17805(n17805), 
         .n17804(n17804), .n17803(n17803), .n17802(n17802), .n17801(n17801), 
         .n17800(n17800), .n17799(n17799), .\data_in[3] ({\data_in[3] }), 
         .n17798(n17798), .n17797(n17797), .n17796(n17796), .n17795(n17795), 
         .n17794(n17794), .n17793(n17793), .n17792(n17792), .n17791(n17791), 
         .\data_in[2] ({\data_in[2] }), .n17790(n17790), .n17789(n17789), 
         .n17788(n17788), .n17787(n17787), .n17786(n17786), .n17785(n17785), 
         .n17784(n17784), .n17783(n17783), .\data_in[1] ({\data_in[1] }), 
         .n17782(n17782), .n17781(n17781), .n17780(n17780), .n17779(n17779), 
         .n17778(n17778), .n17777(n17777), .n17776(n17776), .n17775(n17775), 
         .\data_in[0] ({\data_in[0] }), .n17774(n17774), .n17773(n17773), 
         .n17772(n17772), .n17771(n17771), .n17770(n17770), .n17769(n17769), 
         .n17768(n17768), .\Ki[15] (Ki[15]), .n17767(n17767), .\Ki[14] (Ki[14]), 
         .n17766(n17766), .\Ki[13] (Ki[13]), .n17765(n17765), .\Ki[12] (Ki[12]), 
         .n17764(n17764), .\Ki[11] (Ki[11]), .n17763(n17763), .\Ki[10] (Ki[10]), 
         .n17762(n17762), .\Ki[9] (Ki[9]), .n17761(n17761), .\Ki[8] (Ki[8]), 
         .n17760(n17760), .\Ki[7] (Ki[7]), .n17759(n17759), .\Ki[6] (Ki[6]), 
         .n17758(n17758), .\Ki[5] (Ki[5]), .n17757(n17757), .\Ki[4] (Ki[4]), 
         .n17756(n17756), .\Ki[3] (Ki[3]), .n17755(n17755), .\Ki[2] (Ki[2]), 
         .n17754(n17754), .\Ki[1] (Ki[1]), .n17753(n17753), .\Kp[15] (Kp[15]), 
         .n17752(n17752), .\Kp[14] (Kp[14]), .n17751(n17751), .\Kp[13] (Kp[13]), 
         .n17750(n17750), .\Kp[12] (Kp[12]), .n17749(n17749), .\Kp[11] (Kp[11]), 
         .n17748(n17748), .\Kp[10] (Kp[10]), .n17747(n17747), .\Kp[9] (Kp[9]), 
         .n17746(n17746), .\Kp[8] (Kp[8]), .n17745(n17745), .\Kp[7] (Kp[7]), 
         .n17744(n17744), .\Kp[6] (Kp[6]), .n17743(n17743), .\Kp[5] (Kp[5]), 
         .n17742(n17742), .\Kp[4] (Kp[4]), .n17741(n17741), .\Kp[3] (Kp[3]), 
         .n17740(n17740), .\Kp[2] (Kp[2]), .n17739(n17739), .\Kp[1] (Kp[1]), 
         .n17738(n17738), .gearBoxRatio({gearBoxRatio}), .n17737(n17737), 
         .n17736(n17736), .n17735(n17735), .n17734(n17734), .n17733(n17733), 
         .n17732(n17732), .n17731(n17731), .n17730(n17730), .n17729(n17729), 
         .n17728(n17728), .n17727(n17727), .n17726(n17726), .n17725(n17725), 
         .n17724(n17724), .n17723(n17723), .n17722(n17722), .n17721(n17721), 
         .n17720(n17720), .n4593(n4593), .n17719(n17719), .n17718(n17718), 
         .n17717(n17717), .n17716(n17716), .n4387(n4387), .n4397(n4397), 
         .n4396(n4396), .n17714(n17714), .IntegralLimit({IntegralLimit}), 
         .n4395(n4395), .n17713(n17713), .n17712(n17712), .n17711(n17711), 
         .n17710(n17710), .n17709(n17709), .n17708(n17708), .n17707(n17707), 
         .n17706(n17706), .n17705(n17705), .n17704(n17704), .n17703(n17703), 
         .n17702(n17702), .n17701(n17701), .n17700(n17700), .n17699(n17699), 
         .n4399(n4399), .n17698(n17698), .n17697(n17697), .n17696(n17696), 
         .n17695(n17695), .n17694(n17694), .n17693(n17693), .n17692(n17692), 
         .n63(n63_adj_4745), .n4398(n4398), .n4401(n4401), .n4400(n4400), 
         .n4403(n4403), .n4402(n4402), .n18021(n18021), .n18020(n18020), 
         .n18019(n18019), .n18018(n18018), .n18017(n18017), .n18016(n18016), 
         .n18015(n18015), .LED_c(LED_c), .n4405(n4405), .n4404(n4404), 
         .n4407(n4407), .n4406(n4406), .n18014(n18014), .n17616(n17616), 
         .n3894(n3894), .n788(n788), .n34343(n34343), .n17593(n17593), 
         .n17591(n17591), .n17590(n17590), .n17589(n17589), .\Ki[0] (Ki[0]), 
         .n17588(n17588), .\Kp[0] (Kp[0]), .n17587(n17587), .n17445(n17445), 
         .\data_in_frame[6][7] (\data_in_frame[6] [7]), .n2774(n2774), .n122(n122), 
         .n15957(n15957), .n2957(n2957_adj_4671), .n5(n5_adj_4766), .n44342(n44342), 
         .n24190(n24190), .n36526(n36526), .tx_active(tx_active), .n24918(n24918), 
         .n3(n3_adj_5329), .n4394(n4394), .n4393(n4393), .n4392(n4392), 
         .n4391(n4391), .n4390(n4390), .n4389(n4389), .\FRAME_MATCHER.state_31__N_2661[0] (\FRAME_MATCHER.state_31__N_2661 [0]), 
         .n34989(n34989), .n4388(n4388), .n15960(n15960), .n63_adj_3(n63_adj_4657), 
         .n35562(n35562), .n15994(n15994), .n4386(n4386), .n4409(n4409), 
         .n5_adj_4(n5_adj_5340), .n17500(n17500), .\r_Clock_Count[3] (r_Clock_Count_adj_5401[3]), 
         .n17497(n17497), .\r_Clock_Count[4] (r_Clock_Count_adj_5401[4]), 
         .n17494(n17494), .\r_Clock_Count[5] (r_Clock_Count_adj_5401[5]), 
         .n17491(n17491), .\r_Clock_Count[6] (r_Clock_Count_adj_5401[6]), 
         .n17488(n17488), .\r_Clock_Count[7] (r_Clock_Count_adj_5401[7]), 
         .n17485(n17485), .\r_Clock_Count[8] (r_Clock_Count_adj_5401[8]), 
         .n17513(n17513), .r_Bit_Index({r_Bit_Index_adj_5402}), .n17510(n17510), 
         .n17506(n17506), .\r_Clock_Count[1] (r_Clock_Count_adj_5401[1]), 
         .n17503(n17503), .\r_Clock_Count[2] (r_Clock_Count_adj_5401[2]), 
         .r_SM_Main({r_SM_Main_adj_5400}), .n17637(n17637), .n313(n313), 
         .n314(n314), .n315(n315), .n316(n316), .n317(n317), .n318(n318), 
         .n319(n319), .n320(n320), .VCC_net(VCC_net), .n17505(n17505), 
         .tx_o(tx_o), .tx_enable(tx_enable), .n17607(n17607), .n17606(n17606), 
         .n17605(n17605), .n19670(n19670), .n4(n4_adj_5272), .n4720(n4720), 
         .n17256(n17256), .n17385(n17385), .n3_adj_5(n3_adj_5267), .n8950(n8950), 
         .n29(n29), .n17537(n17537), .r_Bit_Index_adj_14({r_Bit_Index}), 
         .n17540(n17540), .n24794(n24794), .\r_SM_Main[1]_adj_9 (r_SM_Main[1]), 
         .r_Rx_Data(r_Rx_Data), .PIN_13_N_105(PIN_13_N_105), .\r_SM_Main[2]_adj_10 (r_SM_Main[2]), 
         .n15851(n15851), .n15740(n15740), .n17250(n17250), .n40690(n40690), 
         .n40689(n40689), .n17656(n17656), .n17623(n17623), .n17622(n17622), 
         .n17621(n17621), .n17620(n17620), .n17619(n17619), .n17618(n17618), 
         .n17598(n17598), .n17541(n17541), .n43694(n43694), .n17376(n17376), 
         .n4698(n4698), .n23989(n23989), .n4_adj_11(n4_adj_4704), .n4_adj_12(n4_adj_4715), 
         .n4_adj_13(n4)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(183[8] 205[4])
    SB_LUT4 div_46_i1399_3_lut_3_lut (.I0(n2093), .I1(n6075), .I2(n2074), 
            .I3(GND_net), .O(n2173));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1399_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12705_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n36533), .I3(GND_net), .O(n17444));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12706_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n4593), .I3(GND_net), .O(n17445));   // verilog/coms.v(127[12] 295[6])
    defparam i12706_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34509_2_lut (.I0(n24984), .I1(start), .I2(GND_net), .I3(GND_net), 
            .O(n40730));   // verilog/neopixel.v(35[12] 117[6])
    defparam i34509_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i31_4_lut (.I0(n40730), .I1(n40728), .I2(state[1]), .I3(\neo_pixel_transmitter.done ), 
            .O(n33675));   // verilog/neopixel.v(35[12] 117[6])
    defparam i31_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i12848_3_lut (.I0(gearBoxRatio[0]), .I1(\data_in_frame[22] [0]), 
            .I2(n4593), .I3(GND_net), .O(n17587));   // verilog/coms.v(127[12] 295[6])
    defparam i12848_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12849_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n36556), 
            .I3(GND_net), .O(n17588));   // verilog/coms.v(127[12] 295[6])
    defparam i12849_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12850_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n36556), 
            .I3(GND_net), .O(n17589));   // verilog/coms.v(127[12] 295[6])
    defparam i12850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13497_3_lut (.I0(setpoint[7]), .I1(n4393), .I2(n37622), .I3(GND_net), 
            .O(n18236));   // verilog/coms.v(127[12] 295[6])
    defparam i13497_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12851_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n17590));   // verilog/coms.v(127[12] 295[6])
    defparam i12851_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1407_3_lut_3_lut (.I0(n2093), .I1(n6083), .I2(n2082), 
            .I3(GND_net), .O(n2181));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1407_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13496_3_lut (.I0(setpoint[6]), .I1(n4392), .I2(n37622), .I3(GND_net), 
            .O(n18235));   // verilog/coms.v(127[12] 295[6])
    defparam i13496_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1468_3_lut_3_lut (.I0(n2192), .I1(n6097), .I2(n2177), 
            .I3(GND_net), .O(n2273));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1468_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12852_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n4593), .I3(GND_net), .O(n17591));   // verilog/coms.v(127[12] 295[6])
    defparam i12852_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13495_3_lut (.I0(setpoint[5]), .I1(n4391), .I2(n37622), .I3(GND_net), 
            .O(n18234));   // verilog/coms.v(127[12] 295[6])
    defparam i13495_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13494_3_lut (.I0(setpoint[4]), .I1(n4390), .I2(n37622), .I3(GND_net), 
            .O(n18233));   // verilog/coms.v(127[12] 295[6])
    defparam i13494_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12854_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n4593), .I3(GND_net), .O(n17593));   // verilog/coms.v(127[12] 295[6])
    defparam i12854_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1459_3_lut_3_lut (.I0(n2192), .I1(n6088), .I2(n2168), 
            .I3(GND_net), .O(n2264));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1459_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13493_3_lut (.I0(setpoint[3]), .I1(n4389), .I2(n37622), .I3(GND_net), 
            .O(n18232));   // verilog/coms.v(127[12] 295[6])
    defparam i13493_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12855_3_lut (.I0(encoder0_position[0]), .I1(n3016), .I2(count_enable), 
            .I3(GND_net), .O(n17594));   // quad.v(35[10] 41[6])
    defparam i12855_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31792_4_lut (.I0(n15960), .I1(n15957), .I2(n788), .I3(n2957_adj_4671), 
            .O(n38562));
    defparam i31792_4_lut.LUT_INIT = 16'hfac8;
    SB_LUT4 i1_4_lut_adj_1940 (.I0(n63_adj_4657), .I1(\FRAME_MATCHER.state_31__N_2661 [0]), 
            .I2(n5_adj_5340), .I3(n38562), .O(n34343));   // verilog/coms.v(127[12] 295[6])
    defparam i1_4_lut_adj_1940.LUT_INIT = 16'hd5dd;
    SB_LUT4 i12857_3_lut (.I0(encoder1_position[0]), .I1(n2966), .I2(count_enable_adj_4680), 
            .I3(GND_net), .O(n17596));   // quad.v(35[10] 41[6])
    defparam i12857_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13492_3_lut (.I0(setpoint[2]), .I1(n4388), .I2(n37622), .I3(GND_net), 
            .O(n18231));   // verilog/coms.v(127[12] 295[6])
    defparam i13492_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1469_3_lut_3_lut (.I0(n2192), .I1(n6098), .I2(n2178), 
            .I3(GND_net), .O(n2274));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1469_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1473_3_lut_3_lut (.I0(n2192), .I1(n6102), .I2(n2182), 
            .I3(GND_net), .O(n2278));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1473_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1472_3_lut_3_lut (.I0(n2192), .I1(n6101), .I2(n2181), 
            .I3(GND_net), .O(n2277));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1472_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1475_3_lut_3_lut (.I0(n2192), .I1(n6104), .I2(n1059), 
            .I3(GND_net), .O(n2280));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1475_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12858_3_lut (.I0(quadB_debounced), .I1(reg_B[0]), .I2(n36518), 
            .I3(GND_net), .O(n17597));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i12858_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12859_2_lut (.I0(r_SM_Main[2]), .I1(n43694), .I2(GND_net), 
            .I3(GND_net), .O(n17598));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12859_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 div_46_i1463_3_lut_3_lut (.I0(n2192), .I1(n6092), .I2(n2172), 
            .I3(GND_net), .O(n2268));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1463_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1462_3_lut_3_lut (.I0(n2192), .I1(n6091), .I2(n2171), 
            .I3(GND_net), .O(n2267));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1462_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1461_3_lut_3_lut (.I0(n2192), .I1(n6090), .I2(n2170), 
            .I3(GND_net), .O(n2266));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1461_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12746_4_lut (.I0(n17505), .I1(r_Clock_Count_adj_5401[8]), .I2(n313), 
            .I3(r_SM_Main_adj_5400[2]), .O(n17485));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12746_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 div_46_i1464_3_lut_3_lut (.I0(n2192), .I1(n6093), .I2(n2173), 
            .I3(GND_net), .O(n2269));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1464_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12749_4_lut (.I0(n17505), .I1(r_Clock_Count_adj_5401[7]), .I2(n314), 
            .I3(r_SM_Main_adj_5400[2]), .O(n17488));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12749_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 div_46_i1460_3_lut_3_lut (.I0(n2192), .I1(n6089), .I2(n2169), 
            .I3(GND_net), .O(n2265));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1460_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12752_4_lut (.I0(n17505), .I1(r_Clock_Count_adj_5401[6]), .I2(n315), 
            .I3(r_SM_Main_adj_5400[2]), .O(n17491));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12752_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 div_46_i1470_3_lut_3_lut (.I0(n2192), .I1(n6099), .I2(n2179), 
            .I3(GND_net), .O(n2275));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1470_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12755_4_lut (.I0(n17505), .I1(r_Clock_Count_adj_5401[5]), .I2(n316), 
            .I3(r_SM_Main_adj_5400[2]), .O(n17494));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12755_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 div_46_i1471_3_lut_3_lut (.I0(n2192), .I1(n6100), .I2(n2180), 
            .I3(GND_net), .O(n2276));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1471_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1474_3_lut_3_lut (.I0(n2192), .I1(n6103), .I2(n2183), 
            .I3(GND_net), .O(n2279));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1474_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1467_3_lut_3_lut (.I0(n2192), .I1(n6096), .I2(n2176), 
            .I3(GND_net), .O(n2272));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1467_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1465_3_lut_3_lut (.I0(n2192), .I1(n6094), .I2(n2174), 
            .I3(GND_net), .O(n2270));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1465_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i21120_3_lut (.I0(bit_ctr[1]), .I1(n40620), .I2(n4483), .I3(GND_net), 
            .O(n18307));
    defparam i21120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1466_3_lut_3_lut (.I0(n2192), .I1(n6095), .I2(n2175), 
            .I3(GND_net), .O(n2271));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1466_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1533_3_lut_3_lut (.I0(n2288), .I1(n6118), .I2(n2275), 
            .I3(GND_net), .O(n2368));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1533_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1522_3_lut_3_lut (.I0(n2288), .I1(n6107), .I2(n2264), 
            .I3(GND_net), .O(n2357));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1522_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1523_3_lut_3_lut (.I0(n2288), .I1(n6108), .I2(n2265), 
            .I3(GND_net), .O(n2358));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1523_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12866_3_lut (.I0(tx_o), .I1(n3_adj_5267), .I2(r_SM_Main_adj_5400[2]), 
            .I3(GND_net), .O(n17605));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12866_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12867_4_lut (.I0(tx_active), .I1(r_SM_Main_adj_5400[1]), .I2(n8950), 
            .I3(n4_adj_5272), .O(n17606));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12867_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 div_46_i1525_3_lut_3_lut (.I0(n2288), .I1(n6110), .I2(n2267), 
            .I3(GND_net), .O(n2360));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1525_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1526_3_lut_3_lut (.I0(n2288), .I1(n6111), .I2(n2268), 
            .I3(GND_net), .O(n2361));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1526_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1535_3_lut_3_lut (.I0(n2288), .I1(n6120), .I2(n2277), 
            .I3(GND_net), .O(n2370));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1535_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12868_4_lut (.I0(r_SM_Main_adj_5400[2]), .I1(n29), .I2(n19670), 
            .I3(r_SM_Main_adj_5400[0]), .O(n17607));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12868_4_lut.LUT_INIT = 16'h0544;
    SB_LUT4 i12869_3_lut (.I0(quadB_debounced_adj_4679), .I1(reg_B_adj_5411[0]), 
            .I2(n36342), .I3(GND_net), .O(n17608));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    defparam i12869_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36718_1_lut_2_lut (.I0(n3362), .I1(n10244), .I2(GND_net), 
            .I3(GND_net), .O(n43565));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i36718_1_lut_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 div_46_i1532_3_lut_3_lut (.I0(n2288), .I1(n6117), .I2(n2274), 
            .I3(GND_net), .O(n2367));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1532_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1531_3_lut_3_lut (.I0(n2288), .I1(n6116), .I2(n2273), 
            .I3(GND_net), .O(n2366));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1531_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1530_3_lut_3_lut (.I0(n2288), .I1(n6115), .I2(n2272), 
            .I3(GND_net), .O(n2365));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1530_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1529_3_lut_3_lut (.I0(n2288), .I1(n6114), .I2(n2271), 
            .I3(GND_net), .O(n2364));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1529_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i21123_3_lut (.I0(bit_ctr[2]), .I1(n40619), .I2(n4483), .I3(GND_net), 
            .O(n17458));
    defparam i21123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12877_3_lut (.I0(setpoint[0]), .I1(n4386), .I2(n37622), .I3(GND_net), 
            .O(n17616));   // verilog/coms.v(127[12] 295[6])
    defparam i12877_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i107_1_lut_4_lut (.I0(n99), .I1(n16003), .I2(n224), 
            .I3(n558), .O(n249));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i107_1_lut_4_lut.LUT_INIT = 16'h2220;
    SB_LUT4 div_46_i1528_3_lut_3_lut (.I0(n2288), .I1(n6113), .I2(n2270), 
            .I3(GND_net), .O(n2363));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1528_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut (.I0(n98), .I1(n97), .I2(n96), .I3(n15971), 
            .O(n16003));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hff7f;
    SB_LUT4 i12878_3_lut (.I0(\half_duty[0] [0]), .I1(half_duty_new[0]), 
            .I2(n1170), .I3(GND_net), .O(n17617));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i12878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 div_46_i1524_3_lut_3_lut (.I0(n2288), .I1(n6109), .I2(n2266), 
            .I3(GND_net), .O(n2359));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1524_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut_adj_1941 (.I0(n97), .I1(n96), .I2(n15971), 
            .I3(GND_net), .O(n15996));
    defparam i1_2_lut_3_lut_adj_1941.LUT_INIT = 16'hf7f7;
    SB_LUT4 i12879_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n15740), 
            .I3(n23989), .O(n17618));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12879_4_lut.LUT_INIT = 16'hcacc;
    SB_LUT4 div_46_i1539_3_lut_3_lut (.I0(n2288), .I1(n6124), .I2(n1060), 
            .I3(GND_net), .O(n2374));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1539_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12880_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_4704), 
            .I3(n15851), .O(n17619));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12880_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_adj_1942 (.I0(n95), .I1(n94), .I2(n93), .I3(n15877), 
            .O(n15971));
    defparam i1_2_lut_4_lut_adj_1942.LUT_INIT = 16'hff7f;
    SB_LUT4 div_46_i1534_3_lut_3_lut (.I0(n2288), .I1(n6119), .I2(n2276), 
            .I3(GND_net), .O(n2369));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1534_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut_adj_1943 (.I0(n94), .I1(n93), .I2(n15877), 
            .I3(GND_net), .O(n15864));
    defparam i1_2_lut_3_lut_adj_1943.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_46_i1527_3_lut_3_lut (.I0(n2288), .I1(n6112), .I2(n2269), 
            .I3(GND_net), .O(n2362));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1527_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12881_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n15740), 
            .I3(n4_adj_4704), .O(n17620));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12881_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i1_2_lut_4_lut_adj_1944 (.I0(n92), .I1(n91), .I2(n90), .I3(n15974), 
            .O(n15877));
    defparam i1_2_lut_4_lut_adj_1944.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1945 (.I0(n91), .I1(n90), .I2(n15974), 
            .I3(GND_net), .O(n15880));
    defparam i1_2_lut_3_lut_adj_1945.LUT_INIT = 16'hf7f7;
    SB_LUT4 i12882_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_4715), 
            .I3(n15851), .O(n17621));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12882_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12883_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n15740), 
            .I3(n4_adj_4715), .O(n17622));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12883_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 div_46_i1538_3_lut_3_lut (.I0(n2288), .I1(n6123), .I2(n2280), 
            .I3(GND_net), .O(n2373));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1538_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i13513_3_lut (.I0(setpoint[23]), .I1(n4409), .I2(n37622), 
            .I3(GND_net), .O(n18252));   // verilog/coms.v(127[12] 295[6])
    defparam i13513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_4_lut_adj_1946 (.I0(n89), .I1(n88), .I2(n87), .I3(n15893), 
            .O(n15974));
    defparam i1_2_lut_4_lut_adj_1946.LUT_INIT = 16'hff7f;
    SB_LUT4 div_46_i1537_3_lut_3_lut (.I0(n2288), .I1(n6122), .I2(n2279), 
            .I3(GND_net), .O(n2372));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1537_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut_adj_1947 (.I0(n88), .I1(n87), .I2(n15893), 
            .I3(GND_net), .O(n15889));
    defparam i1_2_lut_3_lut_adj_1947.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1948 (.I0(n86), .I1(n85), .I2(n84), .I3(n15901), 
            .O(n15893));
    defparam i1_2_lut_4_lut_adj_1948.LUT_INIT = 16'hff7f;
    SB_LUT4 div_46_i1536_3_lut_3_lut (.I0(n2288), .I1(n6121), .I2(n2278), 
            .I3(GND_net), .O(n2371));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1536_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1595_3_lut_3_lut (.I0(n2381), .I1(n6139), .I2(n2369), 
            .I3(GND_net), .O(n2459));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1595_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1583_3_lut_3_lut (.I0(n2381), .I1(n6127), .I2(n2357), 
            .I3(GND_net), .O(n2447));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1583_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut_adj_1949 (.I0(n85), .I1(n84), .I2(n15901), 
            .I3(GND_net), .O(n15980));
    defparam i1_2_lut_3_lut_adj_1949.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_46_i1584_3_lut_3_lut (.I0(n2381), .I1(n6128), .I2(n2358), 
            .I3(GND_net), .O(n2448));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1584_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1587_3_lut_3_lut (.I0(n2381), .I1(n6131), .I2(n2361), 
            .I3(GND_net), .O(n2451));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1587_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i20253_4_lut (.I0(n954), .I1(n953), .I2(n35948), .I3(n955), 
            .O(n986));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i20253_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 div_46_i1588_3_lut_3_lut (.I0(n2381), .I1(n6132), .I2(n2362), 
            .I3(GND_net), .O(n2452));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1588_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut_adj_1950 (.I0(n83), .I1(n82), .I2(n81), .I3(n15987), 
            .O(n15901));
    defparam i1_2_lut_4_lut_adj_1950.LUT_INIT = 16'hff7f;
    SB_LUT4 i1_2_lut_3_lut_adj_1951 (.I0(n82), .I1(n81), .I2(n15987), 
            .I3(GND_net), .O(n16000));
    defparam i1_2_lut_3_lut_adj_1951.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_46_i1585_3_lut_3_lut (.I0(n2381), .I1(n6129), .I2(n2359), 
            .I3(GND_net), .O(n2449));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1585_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1586_3_lut_3_lut (.I0(n2381), .I1(n6130), .I2(n2360), 
            .I3(GND_net), .O(n2450));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1586_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut_adj_1952 (.I0(n80), .I1(n79), .I2(n78), .I3(n77), 
            .O(n15987));
    defparam i1_2_lut_4_lut_adj_1952.LUT_INIT = 16'hff7f;
    SB_LUT4 div_46_i1601_3_lut_3_lut (.I0(n2381), .I1(n6145), .I2(n1061), 
            .I3(GND_net), .O(n2465));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1601_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1597_3_lut_3_lut (.I0(n2381), .I1(n6141), .I2(n2371), 
            .I3(GND_net), .O(n2461));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1597_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1598_3_lut_3_lut (.I0(n2381), .I1(n6142), .I2(n2372), 
            .I3(GND_net), .O(n2462));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1598_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1594_3_lut_3_lut (.I0(n2381), .I1(n6138), .I2(n2368), 
            .I3(GND_net), .O(n2458));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1594_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1593_3_lut_3_lut (.I0(n2381), .I1(n6137), .I2(n2367), 
            .I3(GND_net), .O(n2457));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1593_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_3_lut_adj_1953 (.I0(n79), .I1(n78), .I2(n77), .I3(GND_net), 
            .O(n15904));
    defparam i1_2_lut_3_lut_adj_1953.LUT_INIT = 16'hf7f7;
    SB_LUT4 div_46_i1592_3_lut_3_lut (.I0(n2381), .I1(n6136), .I2(n2366), 
            .I3(GND_net), .O(n2456));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1592_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1591_3_lut_3_lut (.I0(n2381), .I1(n6135), .I2(n2365), 
            .I3(GND_net), .O(n2455));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1591_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1590_3_lut_3_lut (.I0(n2381), .I1(n6134), .I2(n2364), 
            .I3(GND_net), .O(n2454));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1590_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i1_2_lut_4_lut_adj_1954 (.I0(\FRAME_MATCHER.state [1]), .I1(n24190), 
            .I2(\FRAME_MATCHER.state [3]), .I3(n15963), .O(n34978));   // verilog/coms.v(127[12] 295[6])
    defparam i1_2_lut_4_lut_adj_1954.LUT_INIT = 16'h0008;
    SB_LUT4 div_46_i1596_3_lut_3_lut (.I0(n2381), .I1(n6140), .I2(n2370), 
            .I3(GND_net), .O(n2460));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1596_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1589_3_lut_3_lut (.I0(n2381), .I1(n6133), .I2(n2363), 
            .I3(GND_net), .O(n2453));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1589_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1600_3_lut_3_lut (.I0(n2381), .I1(n6144), .I2(n2374), 
            .I3(GND_net), .O(n2464));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1600_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1599_3_lut_3_lut (.I0(n2381), .I1(n6143), .I2(n2373), 
            .I3(GND_net), .O(n2463));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1599_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i22771_3_lut_4_lut (.I0(n510), .I1(n99), .I2(n511), .I3(n558), 
            .O(n4_adj_5252));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i22771_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i22739_3_lut_4_lut (.I0(n649), .I1(n99), .I2(n650), .I3(n558), 
            .O(n4_adj_5269));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i22739_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i22699_3_lut_4_lut (.I0(n785), .I1(n99), .I2(n786), .I3(n558), 
            .O(n4_adj_4672));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam i22699_3_lut_4_lut.LUT_INIT = 16'heee8;
    SB_LUT4 i13275_3_lut (.I0(\data_in_frame[10] [0]), .I1(rx_data[0]), 
            .I2(n34989), .I3(GND_net), .O(n18014));   // verilog/coms.v(127[12] 295[6])
    defparam i13275_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21099_3_lut (.I0(color[10]), .I1(color[11]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n5_adj_4675));   // verilog/neopixel.v(18[12:19])
    defparam i21099_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34_4_lut (.I0(color[12]), .I1(bit_ctr[0]), .I2(bit_ctr[2]), 
            .I3(color[9]), .O(n29_adj_4674));   // verilog/neopixel.v(18[12:19])
    defparam i34_4_lut.LUT_INIT = 16'h2c20;
    SB_LUT4 i50_4_lut (.I0(n29_adj_4674), .I1(n5_adj_4675), .I2(bit_ctr[1]), 
            .I3(bit_ctr[2]), .O(n35));
    defparam i50_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31748_4_lut (.I0(state_3__N_362[1]), .I1(n3209_adj_5249), .I2(bit_ctr[3]), 
            .I3(n24824), .O(n38513));
    defparam i31748_4_lut.LUT_INIT = 16'hbeee;
    SB_LUT4 i3_4_lut_adj_1955 (.I0(n38513), .I1(n35), .I2(bit_ctr[3]), 
            .I3(n24824), .O(state_3__N_362[0]));
    defparam i3_4_lut_adj_1955.LUT_INIT = 16'h0440;
    SB_LUT4 i12884_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4), .I3(n15851), 
            .O(n17623));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12884_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12886_4_lut (.I0(n35833), .I1(state[1]), .I2(state_3__N_362[1]), 
            .I3(n17203), .O(n17625));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12886_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 div_46_LessThan_985_i32_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1536), 
            .I3(GND_net), .O(n32_adj_4962));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_985_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33972_2_lut_4_lut (.I0(n1531), .I1(n92), .I2(n1535), .I3(n96), 
            .O(n40818));
    defparam i33972_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_985_i34_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1531), 
            .I3(GND_net), .O(n34_adj_4964));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_985_i34_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_4_lut_4_lut (.I0(n15960), .I1(n63_adj_4745), .I2(n788), 
            .I3(n3_adj_5329), .O(n5_adj_5338));   // verilog/coms.v(127[12] 295[6])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hcc04;
    SB_LUT4 div_46_LessThan_1062_i30_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1651), 
            .I3(GND_net), .O(n30_adj_4974));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1062_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33948_2_lut_4_lut (.I0(n1646), .I1(n92), .I2(n1650), .I3(n96), 
            .O(n40794));
    defparam i33948_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1062_i32_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1646), 
            .I3(GND_net), .O(n32_adj_4976));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1062_i32_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1137_i28_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1763), 
            .I3(GND_net), .O(n28_adj_4987));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1137_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33922_2_lut_4_lut (.I0(n1758), .I1(n92), .I2(n1762), .I3(n96), 
            .O(n40768));
    defparam i33922_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1137_i30_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1758), 
            .I3(GND_net), .O(n30_adj_4989));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1137_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34599_2_lut_4_lut (.I0(n1869), .I1(n94), .I2(n1870), .I3(n95), 
            .O(n41446));
    defparam i34599_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1210_i30_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1869), 
            .I3(GND_net), .O(n30_adj_5003));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1210_i30_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1210_i26_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1872), 
            .I3(GND_net), .O(n26_adj_4999));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1210_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34583_2_lut_4_lut (.I0(n1867), .I1(n92), .I2(n1871), .I3(n96), 
            .O(n41430));
    defparam i34583_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1210_i28_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1867), 
            .I3(GND_net), .O(n28_adj_5001));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1210_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1281_i24_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n1978), 
            .I3(GND_net), .O(n24_adj_5013));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1281_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34521_2_lut_4_lut (.I0(n1973), .I1(n92), .I2(n1977), .I3(n96), 
            .O(n41368));
    defparam i34521_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1281_i26_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n1973), 
            .I3(GND_net), .O(n26_adj_5015));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1281_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34538_2_lut_4_lut (.I0(n1975), .I1(n94), .I2(n1976), .I3(n95), 
            .O(n41385));
    defparam i34538_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1281_i28_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n1975), 
            .I3(GND_net), .O(n28_adj_5017));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1281_i28_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_2_lut_3_lut_adj_1956 (.I0(n852), .I1(n6_adj_4668), .I2(n746), 
            .I3(GND_net), .O(n884));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i1_2_lut_3_lut_adj_1956.LUT_INIT = 16'h8080;
    SB_LUT4 div_46_LessThan_1350_i22_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2081), 
            .I3(GND_net), .O(n22_adj_5031));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1350_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i28927_2_lut_3_lut (.I0(n852), .I1(n6_adj_4668), .I2(n746), 
            .I3(GND_net), .O(n953));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i28927_2_lut_3_lut.LUT_INIT = 16'h7070;
    SB_LUT4 i34467_2_lut_4_lut (.I0(n2076), .I1(n92), .I2(n2080), .I3(n96), 
            .O(n41314));
    defparam i34467_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1350_i24_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2076), 
            .I3(GND_net), .O(n24_adj_5033));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1350_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34477_2_lut_4_lut (.I0(n2078), .I1(n94), .I2(n2079), .I3(n95), 
            .O(n41324));
    defparam i34477_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1350_i26_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2078), 
            .I3(GND_net), .O(n26_adj_5035));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1350_i26_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 rem_4_i585_3_lut_4_lut (.I0(n749), .I1(n855), .I2(n884), .I3(n748), 
            .O(n955));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam rem_4_i585_3_lut_4_lut.LUT_INIT = 16'hef10;
    SB_LUT4 i23008_2_lut_3_lut (.I0(n749), .I1(n855), .I2(n748), .I3(GND_net), 
            .O(n6_adj_4668));   // verilog/TinyFPGA_B.v(54[6:33])
    defparam i23008_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 div_46_LessThan_1417_i20_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2181), 
            .I3(GND_net), .O(n20_adj_5048));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34411_2_lut_4_lut (.I0(n2176), .I1(n92), .I2(n2180), .I3(n96), 
            .O(n41258));
    defparam i34411_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1417_i22_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2176), 
            .I3(GND_net), .O(n22_adj_5050));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1417_i24_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2178), 
            .I3(GND_net), .O(n24_adj_5052));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1417_i24_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34425_2_lut_4_lut (.I0(n2178), .I1(n94), .I2(n2179), .I3(n95), 
            .O(n41272));
    defparam i34425_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1482_i18_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2278), 
            .I3(GND_net), .O(n18_adj_5068));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34365_2_lut_4_lut (.I0(n2273), .I1(n92), .I2(n2277), .I3(n96), 
            .O(n41212));
    defparam i34365_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1482_i20_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2273), 
            .I3(GND_net), .O(n20_adj_5070));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1482_i22_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2275), 
            .I3(GND_net), .O(n22_adj_5072));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1482_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34375_2_lut_4_lut (.I0(n2275), .I1(n94), .I2(n2276), .I3(n95), 
            .O(n41222));
    defparam i34375_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1545_i16_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2372), 
            .I3(GND_net), .O(n16_adj_5086));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34275_2_lut_4_lut (.I0(n2367), .I1(n92), .I2(n2371), .I3(n96), 
            .O(n41122));
    defparam i34275_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1545_i18_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2367), 
            .I3(GND_net), .O(n18_adj_5088));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1545_i20_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2369), 
            .I3(GND_net), .O(n20_adj_5090));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i13276_3_lut (.I0(\data_in_frame[10] [1]), .I1(rx_data[1]), 
            .I2(n34989), .I3(GND_net), .O(n18015));   // verilog/coms.v(127[12] 295[6])
    defparam i13276_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i34207_2_lut_4_lut (.I0(n2359), .I1(n84), .I2(n2368), .I3(n93), 
            .O(n41053));
    defparam i34207_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1545_i22_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2359), 
            .I3(GND_net), .O(n22_adj_5092));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1545_i22_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1606_i14_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2463), 
            .I3(GND_net), .O(n14_adj_5108));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34172_2_lut_4_lut (.I0(n2458), .I1(n92), .I2(n2462), .I3(n96), 
            .O(n41018));
    defparam i34172_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_i1659_3_lut_3_lut (.I0(n2471), .I1(n6165), .I2(n2464), 
            .I3(GND_net), .O(n2551));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1659_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1606_i16_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2458), 
            .I3(GND_net), .O(n16_adj_5110));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i1642_3_lut_3_lut (.I0(n2471), .I1(n6148), .I2(n2447), 
            .I3(GND_net), .O(n2534));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1642_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1643_3_lut_3_lut (.I0(n2471), .I1(n6149), .I2(n2448), 
            .I3(GND_net), .O(n2535));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1643_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1644_3_lut_3_lut (.I0(n2471), .I1(n6150), .I2(n2449), 
            .I3(GND_net), .O(n2536));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1644_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1606_i18_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2460), 
            .I3(GND_net), .O(n18_adj_5112));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_i1645_3_lut_3_lut (.I0(n2471), .I1(n6151), .I2(n2450), 
            .I3(GND_net), .O(n2537));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1645_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1647_3_lut_3_lut (.I0(n2471), .I1(n6153), .I2(n2452), 
            .I3(GND_net), .O(n2539));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1647_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i34111_2_lut_4_lut (.I0(n2450), .I1(n84), .I2(n2459), .I3(n93), 
            .O(n40957));
    defparam i34111_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1606_i20_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2450), 
            .I3(GND_net), .O(n20_adj_5114));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1606_i20_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i1_3_lut_4_lut_adj_1957 (.I0(n855), .I1(n884), .I2(n956), 
            .I3(n958), .O(n35948));
    defparam i1_3_lut_4_lut_adj_1957.LUT_INIT = 16'hfff6;
    SB_LUT4 div_46_i1648_3_lut_3_lut (.I0(n2471), .I1(n6154), .I2(n2453), 
            .I3(GND_net), .O(n2540));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1648_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1661_3_lut_3_lut (.I0(n2471), .I1(n6167), .I2(n1062), 
            .I3(GND_net), .O(n2553));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1661_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1646_3_lut_3_lut (.I0(n2471), .I1(n6152), .I2(n2451), 
            .I3(GND_net), .O(n2538));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1646_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1650_3_lut_3_lut (.I0(n2471), .I1(n6156), .I2(n2455), 
            .I3(GND_net), .O(n2542));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1650_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1651_3_lut_3_lut (.I0(n2471), .I1(n6157), .I2(n2456), 
            .I3(GND_net), .O(n2543));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1651_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1660_3_lut_3_lut (.I0(n2471), .I1(n6166), .I2(n2465), 
            .I3(GND_net), .O(n2552));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1660_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1655_3_lut_3_lut (.I0(n2471), .I1(n6161), .I2(n2460), 
            .I3(GND_net), .O(n2547));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1655_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1656_3_lut_3_lut (.I0(n2471), .I1(n6162), .I2(n2461), 
            .I3(GND_net), .O(n2548));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1656_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1654_3_lut_3_lut (.I0(n2471), .I1(n6160), .I2(n2459), 
            .I3(GND_net), .O(n2546));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1654_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1653_3_lut_3_lut (.I0(n2471), .I1(n6159), .I2(n2458), 
            .I3(GND_net), .O(n2545));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1653_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1652_3_lut_3_lut (.I0(n2471), .I1(n6158), .I2(n2457), 
            .I3(GND_net), .O(n2544));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1652_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1658_3_lut_3_lut (.I0(n2471), .I1(n6164), .I2(n2463), 
            .I3(GND_net), .O(n2550));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1658_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1657_3_lut_3_lut (.I0(n2471), .I1(n6163), .I2(n2462), 
            .I3(GND_net), .O(n2549));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1657_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1649_3_lut_3_lut (.I0(n2471), .I1(n6155), .I2(n2454), 
            .I3(GND_net), .O(n2541));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1649_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_LessThan_1665_i12_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2551), 
            .I3(GND_net), .O(n12_adj_5130));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34082_2_lut_4_lut (.I0(n2546), .I1(n92), .I2(n2550), .I3(n96), 
            .O(n40928));
    defparam i34082_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1665_i14_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2546), 
            .I3(GND_net), .O(n14_adj_5132));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1665_i16_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2548), 
            .I3(GND_net), .O(n16_adj_5134));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34041_2_lut_4_lut (.I0(n2538), .I1(n84), .I2(n2547), .I3(n93), 
            .O(n40887));
    defparam i34041_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1665_i18_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2538), 
            .I3(GND_net), .O(n18_adj_5136));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1665_i18_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1722_i12_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2631), 
            .I3(GND_net), .O(n12_adj_5154));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1722_i10_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2636), 
            .I3(GND_net), .O(n10_adj_5152));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1722_i14_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2633), 
            .I3(GND_net), .O(n14_adj_5156));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33969_2_lut_4_lut (.I0(n2623), .I1(n84), .I2(n2632), .I3(n93), 
            .O(n40815));
    defparam i33969_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1722_i16_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2623), 
            .I3(GND_net), .O(n16_adj_5158));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1722_i16_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34010_2_lut_4_lut (.I0(n2631), .I1(n92), .I2(n2635), .I3(n96), 
            .O(n40856));
    defparam i34010_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i13277_3_lut (.I0(\data_in_frame[10] [2]), .I1(rx_data[2]), 
            .I2(n34989), .I3(GND_net), .O(n18016));   // verilog/coms.v(127[12] 295[6])
    defparam i13277_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_LessThan_1777_i8_3_lut_3_lut (.I0(n98), .I1(n97), .I2(n2718), 
            .I3(GND_net), .O(n8_adj_5178));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i8_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1777_i12_3_lut_3_lut (.I0(n95), .I1(n94), .I2(n2715), 
            .I3(GND_net), .O(n12_adj_5182));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i12_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i34579_2_lut_4_lut (.I0(n2705), .I1(n84), .I2(n2714), .I3(n93), 
            .O(n41426));
    defparam i34579_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 div_46_LessThan_1777_i14_3_lut_3_lut (.I0(n93), .I1(n84), .I2(n2705), 
            .I3(GND_net), .O(n14_adj_5184));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i14_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 div_46_LessThan_1777_i10_3_lut_3_lut (.I0(n96), .I1(n92), .I2(n2713), 
            .I3(GND_net), .O(n10_adj_5180));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_LessThan_1777_i10_3_lut_3_lut.LUT_INIT = 16'h1717;
    SB_LUT4 i33924_2_lut_4_lut (.I0(n2713), .I1(n92), .I2(n2717), .I3(n96), 
            .O(n40770));
    defparam i33924_2_lut_4_lut.LUT_INIT = 16'hf99f;
    SB_LUT4 i13278_3_lut (.I0(\data_in_frame[10] [3]), .I1(rx_data[3]), 
            .I2(n34989), .I3(GND_net), .O(n18017));   // verilog/coms.v(127[12] 295[6])
    defparam i13278_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13279_3_lut (.I0(\data_in_frame[10] [4]), .I1(rx_data[4]), 
            .I2(n34989), .I3(GND_net), .O(n18018));   // verilog/coms.v(127[12] 295[6])
    defparam i13279_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13280_3_lut (.I0(\data_in_frame[10] [5]), .I1(rx_data[5]), 
            .I2(n34989), .I3(GND_net), .O(n18019));   // verilog/coms.v(127[12] 295[6])
    defparam i13280_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13281_3_lut (.I0(\data_in_frame[10] [6]), .I1(rx_data[6]), 
            .I2(n34989), .I3(GND_net), .O(n18020));   // verilog/coms.v(127[12] 295[6])
    defparam i13281_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13282_3_lut (.I0(\data_in_frame[10] [7]), .I1(rx_data[7]), 
            .I2(n34989), .I3(GND_net), .O(n18021));   // verilog/coms.v(127[12] 295[6])
    defparam i13282_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12917_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n15740), 
            .I3(n4), .O(n17656));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12917_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i12918_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n36533), .I3(GND_net), .O(n17657));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12918_3_lut.LUT_INIT = 16'hacac;
    \quad(DEBOUNCE_TICKS=100)  quad_counter1 (.encoder1_position({encoder1_position}), 
            .GND_net(GND_net), .n18184(n18184), .clk32MHz(clk32MHz), .n18185(n18185), 
            .n18186(n18186), .n18187(n18187), .n18188(n18188), .n18189(n18189), 
            .n18190(n18190), .n18181(n18181), .n18202(n18202), .n18203(n18203), 
            .n18200(n18200), .n18201(n18201), .n18198(n18198), .n18199(n18199), 
            .n18196(n18196), .n18197(n18197), .n18194(n18194), .n18195(n18195), 
            .n18191(n18191), .n18192(n18192), .n18193(n18193), .n18182(n18182), 
            .n18183(n18183), .data_o({quadA_debounced_adj_4678, quadB_debounced_adj_4679}), 
            .n17596(n17596), .n2942({n2943, n2944, n2945, n2946, n2947, 
            n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, 
            n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, 
            n2964, n2965, n2966}), .count_enable(count_enable_adj_4680), 
            .n18229(n18229), .reg_B({reg_B_adj_5411}), .n36342(n36342), 
            .PIN_6_c_1(PIN_6_c_1), .PIN_7_c_0(PIN_7_c_0), .n17608(n17608)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(244[15] 249[4])
    SB_LUT4 i12919_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n36533), .I3(GND_net), .O(n17658));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1716_3_lut_3_lut (.I0(n2558), .I1(n6187), .I2(n2551), 
            .I3(GND_net), .O(n2635));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1716_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1699_3_lut_3_lut (.I0(n2558), .I1(n6170), .I2(n2534), 
            .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1699_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12920_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n36533), .I3(GND_net), .O(n17659));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12920_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1700_3_lut_3_lut (.I0(n2558), .I1(n6171), .I2(n2535), 
            .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1700_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1701_3_lut_3_lut (.I0(n2558), .I1(n6172), .I2(n2536), 
            .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1701_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1702_3_lut_3_lut (.I0(n2558), .I1(n6173), .I2(n2537), 
            .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1702_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12921_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n36533), .I3(GND_net), .O(n17660));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1719_3_lut_3_lut (.I0(n2558), .I1(n6190), .I2(n1063), 
            .I3(GND_net), .O(n2638));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1719_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1705_3_lut_3_lut (.I0(n2558), .I1(n6176), .I2(n2540), 
            .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1705_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1706_3_lut_3_lut (.I0(n2558), .I1(n6177), .I2(n2541), 
            .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1706_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12922_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n36533), .I3(GND_net), .O(n17661));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12922_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12923_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n36533), .I3(GND_net), .O(n17662));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12923_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12924_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n36533), .I3(GND_net), .O(n17663));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12925_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n36533), .I3(GND_net), .O(n17664));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1708_3_lut_3_lut (.I0(n2558), .I1(n6179), .I2(n2543), 
            .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1708_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1709_3_lut_3_lut (.I0(n2558), .I1(n6180), .I2(n2544), 
            .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1709_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1710_3_lut_3_lut (.I0(n2558), .I1(n6181), .I2(n2545), 
            .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1710_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12926_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n36533), .I3(GND_net), .O(n17665));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12927_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n36533), .I3(GND_net), .O(n17666));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12928_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n36533), .I3(GND_net), .O(n17667));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12929_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n36533), .I3(GND_net), .O(n17668));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12930_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n36533), .I3(GND_net), .O(n17669));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12931_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n36533), .I3(GND_net), .O(n17670));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12932_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n36533), .I3(GND_net), .O(n17671));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12932_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1711_3_lut_3_lut (.I0(n2558), .I1(n6182), .I2(n2546), 
            .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1711_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12933_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n36533), .I3(GND_net), .O(n17672));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1717_3_lut_3_lut (.I0(n2558), .I1(n6188), .I2(n2552), 
            .I3(GND_net), .O(n2636));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1717_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12934_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n36533), .I3(GND_net), .O(n17673));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12934_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12935_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n36533), .I3(GND_net), .O(n17674));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12935_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1718_3_lut_3_lut (.I0(n2558), .I1(n6189), .I2(n2553), 
            .I3(GND_net), .O(n2637));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1718_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1712_3_lut_3_lut (.I0(n2558), .I1(n6183), .I2(n2547), 
            .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1712_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12936_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n36533), .I3(GND_net), .O(n17675));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12936_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12937_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n36533), .I3(GND_net), .O(n17676));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12937_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12938_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n36533), .I3(GND_net), .O(n17677));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12938_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12939_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n36533), .I3(GND_net), .O(n17678));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12939_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1707_3_lut_3_lut (.I0(n2558), .I1(n6178), .I2(n2542), 
            .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1707_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12940_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n36533), .I3(GND_net), .O(n17679));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12940_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1714_3_lut_3_lut (.I0(n2558), .I1(n6185), .I2(n2549), 
            .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1714_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12941_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n36533), .I3(GND_net), .O(n17680));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12941_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1704_3_lut_3_lut (.I0(n2558), .I1(n6175), .I2(n2539), 
            .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1704_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12942_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n36533), .I3(GND_net), .O(n17681));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12942_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12943_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n36533), .I3(GND_net), .O(n17682));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12943_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12944_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n36533), .I3(GND_net), .O(n17683));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12944_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12945_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n36533), .I3(GND_net), .O(n17684));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12945_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12946_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n36533), .I3(GND_net), .O(n17685));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12946_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i12947_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n36533), .I3(GND_net), .O(n17686));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12947_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 div_46_i1703_3_lut_3_lut (.I0(n2558), .I1(n6174), .I2(n2538), 
            .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1703_3_lut_3_lut.LUT_INIT = 16'he4e4;
    motorControl control (.GND_net(GND_net), .\Kp[2] (Kp[2]), .\Kp[3] (Kp[3]), 
            .duty({duty}), .IntegralLimit({IntegralLimit}), .\Kp[1] (Kp[1]), 
            .\Kp[0] (Kp[0]), .\Kp[4] (Kp[4]), .\Kp[5] (Kp[5]), .\Kp[6] (Kp[6]), 
            .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), .PWMLimit({PWMLimit}), .\Kp[9] (Kp[9]), 
            .\Kp[10] (Kp[10]), .\Kp[11] (Kp[11]), .\Kp[12] (Kp[12]), .\Kp[13] (Kp[13]), 
            .\Kp[14] (Kp[14]), .\Kp[15] (Kp[15]), .clk32MHz(clk32MHz), 
            .VCC_net(VCC_net), .n25(n25), .\Ki[0] (Ki[0]), .\Ki[3] (Ki[3]), 
            .\Ki[2] (Ki[2]), .\Ki[1] (Ki[1]), .motor_state({motor_state}), 
            .\Ki[4] (Ki[4]), .\Ki[5] (Ki[5]), .\Ki[6] (Ki[6]), .\Ki[7] (Ki[7]), 
            .\Ki[8] (Ki[8]), .\Ki[9] (Ki[9]), .\Ki[10] (Ki[10]), .\Ki[11] (Ki[11]), 
            .\Ki[12] (Ki[12]), .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), 
            .n43653(n43653), .setpoint({setpoint})) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(216[16] 229[4])
    SB_LUT4 div_46_i1715_3_lut_3_lut (.I0(n2558), .I1(n6186), .I2(n2550), 
            .I3(GND_net), .O(n2634));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1715_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 div_46_i1713_3_lut_3_lut (.I0(n2558), .I1(n6184), .I2(n2548), 
            .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(232[21:53])
    defparam div_46_i1713_3_lut_3_lut.LUT_INIT = 16'he4e4;
    SB_LUT4 i12948_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n36533), .I3(GND_net), .O(n17687));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12948_3_lut.LUT_INIT = 16'hacac;
    \quad(DEBOUNCE_TICKS=100)_U1  quad_counter0 (.n18176(n18176), .encoder0_position({encoder0_position}), 
            .clk32MHz(clk32MHz), .n18177(n18177), .n18178(n18178), .n18179(n18179), 
            .n18165(n18165), .n18166(n18166), .n18167(n18167), .n18168(n18168), 
            .n18169(n18169), .n18170(n18170), .n18171(n18171), .n18172(n18172), 
            .n18173(n18173), .n18174(n18174), .n18175(n18175), .n18163(n18163), 
            .n18164(n18164), .n18161(n18161), .n18162(n18162), .n18159(n18159), 
            .n18160(n18160), .n18157(n18157), .n18158(n18158), .data_o({quadA_debounced, 
            quadB_debounced}), .GND_net(GND_net), .n2992({n2993, n2994, 
            n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, 
            n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, 
            n3011, n3012, n3013, n3014, n3015, n3016}), .n17594(n17594), 
            .count_enable(count_enable), .n18213(n18213), .reg_B({reg_B}), 
            .n36518(n36518), .PIN_2_c_0(PIN_2_c_0), .PIN_1_c_1(PIN_1_c_1), 
            .n17597(n17597)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(236[15] 241[4])
    SB_LUT4 i12_3_lut_adj_1958 (.I0(bit_ctr[3]), .I1(n40705), .I2(n4483), 
            .I3(GND_net), .O(n33629));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1958.LUT_INIT = 16'hacac;
    SB_LUT4 i12_3_lut_adj_1959 (.I0(bit_ctr[6]), .I1(n40701), .I2(n4483), 
            .I3(GND_net), .O(n33617));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1959.LUT_INIT = 16'hacac;
    SB_LUT4 i12953_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n4593), .I3(GND_net), .O(n17692));   // verilog/coms.v(127[12] 295[6])
    defparam i12953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12954_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n4593), .I3(GND_net), .O(n17693));   // verilog/coms.v(127[12] 295[6])
    defparam i12954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12955_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n4593), .I3(GND_net), .O(n17694));   // verilog/coms.v(127[12] 295[6])
    defparam i12955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12956_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n4593), .I3(GND_net), .O(n17695));   // verilog/coms.v(127[12] 295[6])
    defparam i12956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12957_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n4593), .I3(GND_net), .O(n17696));   // verilog/coms.v(127[12] 295[6])
    defparam i12957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12958_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n4593), .I3(GND_net), .O(n17697));   // verilog/coms.v(127[12] 295[6])
    defparam i12958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12959_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n4593), .I3(GND_net), .O(n17698));   // verilog/coms.v(127[12] 295[6])
    defparam i12959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12960_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n4593), .I3(GND_net), .O(n17699));   // verilog/coms.v(127[12] 295[6])
    defparam i12960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12961_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n4593), .I3(GND_net), .O(n17700));   // verilog/coms.v(127[12] 295[6])
    defparam i12961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12962_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n4593), .I3(GND_net), .O(n17701));   // verilog/coms.v(127[12] 295[6])
    defparam i12962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12963_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n4593), .I3(GND_net), .O(n17702));   // verilog/coms.v(127[12] 295[6])
    defparam i12963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12964_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n4593), .I3(GND_net), .O(n17703));   // verilog/coms.v(127[12] 295[6])
    defparam i12964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12965_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n4593), .I3(GND_net), .O(n17704));   // verilog/coms.v(127[12] 295[6])
    defparam i12965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12966_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n4593), .I3(GND_net), .O(n17705));   // verilog/coms.v(127[12] 295[6])
    defparam i12966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12967_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n4593), .I3(GND_net), .O(n17706));   // verilog/coms.v(127[12] 295[6])
    defparam i12967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12968_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n4593), .I3(GND_net), .O(n17707));   // verilog/coms.v(127[12] 295[6])
    defparam i12968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12969_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n4593), .I3(GND_net), .O(n17708));   // verilog/coms.v(127[12] 295[6])
    defparam i12969_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12970_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n4593), .I3(GND_net), .O(n17709));   // verilog/coms.v(127[12] 295[6])
    defparam i12970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12971_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n4593), .I3(GND_net), .O(n17710));   // verilog/coms.v(127[12] 295[6])
    defparam i12971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12972_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n4593), .I3(GND_net), .O(n17711));   // verilog/coms.v(127[12] 295[6])
    defparam i12972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12973_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n4593), .I3(GND_net), .O(n17712));   // verilog/coms.v(127[12] 295[6])
    defparam i12973_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12974_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n4593), .I3(GND_net), .O(n17713));   // verilog/coms.v(127[12] 295[6])
    defparam i12974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12975_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n4593), .I3(GND_net), .O(n17714));   // verilog/coms.v(127[12] 295[6])
    defparam i12975_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_3_lut_adj_1960 (.I0(n40702), .I1(bit_ctr[12]), .I2(n4483), 
            .I3(GND_net), .O(n33619));   // verilog/neopixel.v(35[12] 117[6])
    defparam i12_3_lut_adj_1960.LUT_INIT = 16'hcaca;
    SB_LUT4 i12977_3_lut (.I0(gearBoxRatio[1]), .I1(\data_in_frame[22] [1]), 
            .I2(n4593), .I3(GND_net), .O(n17716));   // verilog/coms.v(127[12] 295[6])
    defparam i12977_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12978_3_lut (.I0(gearBoxRatio[2]), .I1(\data_in_frame[22] [2]), 
            .I2(n4593), .I3(GND_net), .O(n17717));   // verilog/coms.v(127[12] 295[6])
    defparam i12978_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12979_3_lut (.I0(gearBoxRatio[3]), .I1(\data_in_frame[22] [3]), 
            .I2(n4593), .I3(GND_net), .O(n17718));   // verilog/coms.v(127[12] 295[6])
    defparam i12979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12980_3_lut (.I0(gearBoxRatio[4]), .I1(\data_in_frame[22] [4]), 
            .I2(n4593), .I3(GND_net), .O(n17719));   // verilog/coms.v(127[12] 295[6])
    defparam i12980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12981_3_lut (.I0(gearBoxRatio[5]), .I1(\data_in_frame[22] [5]), 
            .I2(n4593), .I3(GND_net), .O(n17720));   // verilog/coms.v(127[12] 295[6])
    defparam i12981_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12982_3_lut (.I0(gearBoxRatio[6]), .I1(\data_in_frame[22] [6]), 
            .I2(n4593), .I3(GND_net), .O(n17721));   // verilog/coms.v(127[12] 295[6])
    defparam i12982_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12983_3_lut (.I0(gearBoxRatio[7]), .I1(\data_in_frame[22] [7]), 
            .I2(n4593), .I3(GND_net), .O(n17722));   // verilog/coms.v(127[12] 295[6])
    defparam i12983_3_lut.LUT_INIT = 16'hcaca;
    \pwm(32000000,20000,32000000,23,1)  PWM (.GND_net(GND_net), .VCC_net(VCC_net), 
            .\half_duty_new[0] (half_duty_new[0]), .CLK_c(CLK_c), .PIN_19_c_0(PIN_19_c_0), 
            .pwm_setpoint({pwm_setpoint}), .n18253(n18253), .\half_duty[0][1] (\half_duty[0] [1]), 
            .n18254(n18254), .\half_duty[0][2] (\half_duty[0] [2]), .n18255(n18255), 
            .\half_duty[0][3] (\half_duty[0] [3]), .n18256(n18256), .\half_duty[0][4] (\half_duty[0] [4]), 
            .n18258(n18258), .\half_duty[0][6] (\half_duty[0] [6]), .n18259(n18259), 
            .\half_duty[0][7] (\half_duty[0] [7]), .\half_duty[0][0] (\half_duty[0] [0]), 
            .n1170(n1170), .\half_duty_new[1] (half_duty_new[1]), .\half_duty_new[2] (half_duty_new[2]), 
            .\half_duty_new[3] (half_duty_new[3]), .\half_duty_new[4] (half_duty_new[4]), 
            .\half_duty_new[6] (half_duty_new[6]), .\half_duty_new[7] (half_duty_new[7]), 
            .n17617(n17617)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // verilog/TinyFPGA_B.v(131[43] 137[3])
    SB_LUT4 i12984_3_lut (.I0(gearBoxRatio[8]), .I1(\data_in_frame[21] [0]), 
            .I2(n4593), .I3(GND_net), .O(n17723));   // verilog/coms.v(127[12] 295[6])
    defparam i12984_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12985_3_lut (.I0(gearBoxRatio[9]), .I1(\data_in_frame[21] [1]), 
            .I2(n4593), .I3(GND_net), .O(n17724));   // verilog/coms.v(127[12] 295[6])
    defparam i12985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12986_3_lut (.I0(gearBoxRatio[10]), .I1(\data_in_frame[21] [2]), 
            .I2(n4593), .I3(GND_net), .O(n17725));   // verilog/coms.v(127[12] 295[6])
    defparam i12986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12987_3_lut (.I0(gearBoxRatio[11]), .I1(\data_in_frame[21] [3]), 
            .I2(n4593), .I3(GND_net), .O(n17726));   // verilog/coms.v(127[12] 295[6])
    defparam i12987_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12988_3_lut (.I0(gearBoxRatio[12]), .I1(\data_in_frame[21] [4]), 
            .I2(n4593), .I3(GND_net), .O(n17727));   // verilog/coms.v(127[12] 295[6])
    defparam i12988_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12989_3_lut (.I0(gearBoxRatio[13]), .I1(\data_in_frame[21] [5]), 
            .I2(n4593), .I3(GND_net), .O(n17728));   // verilog/coms.v(127[12] 295[6])
    defparam i12989_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12990_3_lut (.I0(gearBoxRatio[14]), .I1(\data_in_frame[21] [6]), 
            .I2(n4593), .I3(GND_net), .O(n17729));   // verilog/coms.v(127[12] 295[6])
    defparam i12990_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12991_3_lut (.I0(gearBoxRatio[15]), .I1(\data_in_frame[21] [7]), 
            .I2(n4593), .I3(GND_net), .O(n17730));   // verilog/coms.v(127[12] 295[6])
    defparam i12991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12992_3_lut (.I0(gearBoxRatio[16]), .I1(\data_in_frame[20] [0]), 
            .I2(n4593), .I3(GND_net), .O(n17731));   // verilog/coms.v(127[12] 295[6])
    defparam i12992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12993_3_lut (.I0(gearBoxRatio[17]), .I1(\data_in_frame[20] [1]), 
            .I2(n4593), .I3(GND_net), .O(n17732));   // verilog/coms.v(127[12] 295[6])
    defparam i12993_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12994_3_lut (.I0(gearBoxRatio[18]), .I1(\data_in_frame[20] [2]), 
            .I2(n4593), .I3(GND_net), .O(n17733));   // verilog/coms.v(127[12] 295[6])
    defparam i12994_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12995_3_lut (.I0(gearBoxRatio[19]), .I1(\data_in_frame[20] [3]), 
            .I2(n4593), .I3(GND_net), .O(n17734));   // verilog/coms.v(127[12] 295[6])
    defparam i12995_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12996_3_lut (.I0(gearBoxRatio[20]), .I1(\data_in_frame[20] [4]), 
            .I2(n4593), .I3(GND_net), .O(n17735));   // verilog/coms.v(127[12] 295[6])
    defparam i12996_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12997_3_lut (.I0(gearBoxRatio[21]), .I1(\data_in_frame[20] [5]), 
            .I2(n4593), .I3(GND_net), .O(n17736));   // verilog/coms.v(127[12] 295[6])
    defparam i12997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12998_3_lut (.I0(gearBoxRatio[22]), .I1(\data_in_frame[20] [6]), 
            .I2(n4593), .I3(GND_net), .O(n17737));   // verilog/coms.v(127[12] 295[6])
    defparam i12998_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12999_3_lut (.I0(gearBoxRatio[23]), .I1(\data_in_frame[20] [7]), 
            .I2(n4593), .I3(GND_net), .O(n17738));   // verilog/coms.v(127[12] 295[6])
    defparam i12999_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13000_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n36556), 
            .I3(GND_net), .O(n17739));   // verilog/coms.v(127[12] 295[6])
    defparam i13000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13_3_lut (.I0(n3252), .I1(n3231), .I2(n3230), .I3(GND_net), 
            .O(n38_adj_5312));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i13001_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n36556), 
            .I3(GND_net), .O(n17740));   // verilog/coms.v(127[12] 295[6])
    defparam i13001_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13002_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n36556), 
            .I3(GND_net), .O(n17741));   // verilog/coms.v(127[12] 295[6])
    defparam i13002_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13003_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n36556), 
            .I3(GND_net), .O(n17742));   // verilog/coms.v(127[12] 295[6])
    defparam i13003_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13004_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n36556), 
            .I3(GND_net), .O(n17743));   // verilog/coms.v(127[12] 295[6])
    defparam i13004_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13005_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n36556), 
            .I3(GND_net), .O(n17744));   // verilog/coms.v(127[12] 295[6])
    defparam i13005_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13006_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n36556), 
            .I3(GND_net), .O(n17745));   // verilog/coms.v(127[12] 295[6])
    defparam i13006_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13007_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n36556), 
            .I3(GND_net), .O(n17746));   // verilog/coms.v(127[12] 295[6])
    defparam i13007_3_lut.LUT_INIT = 16'hacac;
    
endmodule
//
// Verilog Description of module neopixel
//

module neopixel (\neo_pixel_transmitter.done , clk32MHz, \state_3__N_362[1] , 
            \state[1] , n40674, GND_net, bit_ctr, VCC_net, n33653, 
            n33655, n33657, n33659, n33661, n33663, n33665, n33635, 
            n33639, n33641, n33643, n33645, n33647, n18307, n33589, 
            n33673, n33623, n33667, n33669, n33671, n33649, n33651, 
            n33631, n33633, n33595, n18212, n33601, n33621, timer, 
            n40726, n25779, n40725, n40724, n40723, n40722, n40721, 
            n40720, n40719, n3209, n40718, n40717, n40716, n40715, 
            n40714, n40713, n33619, n33617, n33629, n17687, \neo_pixel_transmitter.t0 , 
            n17686, n17685, n17684, n17683, n17682, n17681, n17680, 
            n17679, n17678, n17677, n17676, n17675, n17674, n17673, 
            n17672, n17671, n17670, n17669, n17668, n17667, n17666, 
            n17665, n17664, n17663, n17662, n17661, n17660, n17659, 
            n17658, n17657, start, \one_wire_N_513[9] , \one_wire_N_513[10] , 
            \one_wire_N_513[6] , \one_wire_N_513[8] , n11, \one_wire_N_513[11] , 
            n4451, n1164, \state[0] , n4483, n40712, n35873, n40709, 
            n40708, n17625, \state_3__N_362[0] , n17203, n35833, n40704, 
            n40703, n17458, PIN_8_c, n37483, n40702, n40700, n33675, 
            n17444, n40699, n40698, n40707, n40706, n40701, n40711, 
            n40710, n40705, n40619, n40620, n40616, n24984, n24782, 
            n24824, n36533) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output \neo_pixel_transmitter.done ;
    input clk32MHz;
    output \state_3__N_362[1] ;
    output \state[1] ;
    output n40674;
    input GND_net;
    output [31:0]bit_ctr;
    input VCC_net;
    input n33653;
    input n33655;
    input n33657;
    input n33659;
    input n33661;
    input n33663;
    input n33665;
    input n33635;
    input n33639;
    input n33641;
    input n33643;
    input n33645;
    input n33647;
    input n18307;
    input n33589;
    input n33673;
    input n33623;
    input n33667;
    input n33669;
    input n33671;
    input n33649;
    input n33651;
    input n33631;
    input n33633;
    input n33595;
    input n18212;
    input n33601;
    input n33621;
    output [31:0]timer;
    output n40726;
    input n25779;
    output n40725;
    output n40724;
    output n40723;
    output n40722;
    output n40721;
    output n40720;
    output n40719;
    output n3209;
    output n40718;
    output n40717;
    output n40716;
    output n40715;
    output n40714;
    output n40713;
    input n33619;
    input n33617;
    input n33629;
    input n17687;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input n17686;
    input n17685;
    input n17684;
    input n17683;
    input n17682;
    input n17681;
    input n17680;
    input n17679;
    input n17678;
    input n17677;
    input n17676;
    input n17675;
    input n17674;
    input n17673;
    input n17672;
    input n17671;
    input n17670;
    input n17669;
    input n17668;
    input n17667;
    input n17666;
    input n17665;
    input n17664;
    input n17663;
    input n17662;
    input n17661;
    input n17660;
    input n17659;
    input n17658;
    input n17657;
    output start;
    output \one_wire_N_513[9] ;
    output \one_wire_N_513[10] ;
    output \one_wire_N_513[6] ;
    output \one_wire_N_513[8] ;
    output n11;
    output \one_wire_N_513[11] ;
    output n4451;
    output n1164;
    output \state[0] ;
    output n4483;
    output n40712;
    input n35873;
    output n40709;
    output n40708;
    input n17625;
    input \state_3__N_362[0] ;
    output n17203;
    output n35833;
    output n40704;
    output n40703;
    input n17458;
    output PIN_8_c;
    input n37483;
    output n40702;
    output n40700;
    input n33675;
    input n17444;
    output n40699;
    output n40698;
    output n40707;
    output n40706;
    output n40701;
    output n40711;
    output n40710;
    output n40705;
    output n40619;
    output n40620;
    output n40616;
    output n24984;
    output n24782;
    output n24824;
    output n36533;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n29235, n2603, n2621, n29236, n2703, n2604, n29234, \neo_pixel_transmitter.done_N_570 , 
        n37672, n2704, n2605, n29233, n2705, n2606, n29232, n2706, 
        n2607, n29231, n1598, n1499, n1532, n27952, n2707, n2608, 
        n29230, n2708, n2609, n43630, n29229, n2709, n1599, n1500, 
        n27951, n2588, n2489, n2522, n29228, n1600, n1501, n27950, 
        n2589, n2490, n29227, n2590, n2491, n29226, n1601, n1502, 
        n27949, n2907, n2909, n33, n2900, n2891, n2897, n2888, 
        n41, n2906, n2887, n2892, n38, n2896, n2885, n2905, 
        n2902, n43, n1602, n1503, n27948, n2899, n2890, n2898, 
        n2908, n40, n2889, n2901, n46, n2886, n2894, n2895, 
        n2903, n39, n2904, n2893, n47, n2918, n1603, n1504, 
        n27947, n2401, n2409, n27, n2390, n2391, n2397, n2407, 
        n33_adj_4527, n2405, n2394, n2400, n2399, n32, n2406, 
        n2396, n2403, n2402, n31, n2393, n2392, n2408, n2398, 
        n35, n2404, n2395, n37, n2423, n2591, n2492, n29225, 
        n2302, n2292, n22, n1604, n1505, n27946, n2299, n2309, 
        n30, n43632, n3017, n43639, n2294, n2306, n2297, n34, 
        n2301, n2307, n2291, n2305, n32_adj_4528, n2592, n2493, 
        n29224, n2298, n2295, n2304, n2300, n33_adj_4529, n2593, 
        n2494, n29223, n2308, n2296, n2303, n2293, n31_adj_4530, 
        n2324, n2594, n2495, n29222, n43633, n1605, n1506, n27945, 
        n1606, n1507, n27944, n2595, n2496, n29221, n1607, n1508, 
        n27943, n2596, n2497, n29220, n2597, n2498, n29219, n2598, 
        n2499, n29218, n1608, n1509, n43631, n27942, n2599, n2500, 
        n29217, n2600, n2501, n29216, n2601, n2502, n29215, n2602, 
        n2503, n29214, n2504, n29213, n1609;
    wire [31:0]n133;
    
    wire n28601, n2505, n29212, n28600, n2506, n29211, n2507, 
        n29210, n28599, n28598, n2508, n29209, n28597, n28596, 
        n28595, n28594, n28593, n28592, n2509, n29208, n28591, 
        n28590, n28589, n28588, n28587, n28586, n28585, n28584, 
        n28583, n28582, n28581, n28580, n29207, n29206, n29205, 
        n28579, n28578, n28577, n29204, n28576, n28575, n29203, 
        n28574, n28573, n28572, n29202, n28571, n29201, n29200, 
        n29199, n29198, n29197, n29196, n27871, n27870, n29195, 
        n29194, n29193, n29192, n27869, n29191, n29190, n29189, 
        n29188, n27868, n29187, n29186, n29185, n29184, n29183, 
        n29182, n29181, n29180, n27867, n29179, n29178, n29177, 
        n29176, n29175, n3182, n3083, n3116, n29375, n27866, n29174, 
        n3183, n3084, n29374, n29173, n3184, n3085, n29373, n29172, 
        n3185, n3086, n29372, n29171, n3186, n3087, n29371, n3187, 
        n3088, n29370, n3188, n3089, n29369, n29170, n3189, n3090, 
        n29368, n43634, n29169, n3190, n3091, n29367, n3191, n3092, 
        n29366, n3192, n3093, n29365, n2192, n2225, n29168, n2193, 
        n29167, n27865, n1998, n2004, n18, n2003, n1999, n1996, 
        n2007, n28, n1997, n2005, n2000, n2002, n26, n2001, 
        n2008, n1994, n1995, n27_adj_4531, n2006, n2009, n25, 
        n3193, n3094, n29364, n2194, n29166, n2027, n2195, n29165, 
        n27864, n3194, n3095, n29363, n2196, n29164, n2197, n29163, 
        n3195, n3096, n29362, n2198, n29162, n2199, n29161, n3196, 
        n3097, n29361, n2200, n29160, n3197, n3098, n29360, n2201, 
        n29159, n2202, n29158, n2203, n29157, n3198, n3099, n29359, 
        n2204, n29156, n2205, n29155, n3199, n3100, n29358, n2206, 
        n29154, n3200, n3101, n29357, n2207, n29153, n3201, n3102, 
        n29356, n2208, n29152, n3202, n3103, n29355, n3203, n3104, 
        n29354, n2209, n43637, n29151, n3204, n3105, n29353, n3205, 
        n3106, n29352, n2093, n2126, n29150, n3206, n3107, n29351, 
        n2094, n29149, n3207, n3108, n29350, n2095, n29148, n2096, 
        n29147, n3208, n3109, n43636, n29349, n2097, n29146, n2984, 
        n29348, n2098, n29145, n2985, n29347, n2099, n29144, n2986, 
        n29346, n2100, n29143, n2987, n29345, n2988, n29344, n2101, 
        n29142, n2102, n29141, n2103, n29140, n2989, n29343, n2990, 
        n29342, n2991, n29341, n2992, n29340, n2104, n29139, n2993, 
        n29339, n2105, n29138, n27863, n2106, n29137, n2994, n29338, 
        n2107, n29136, n2108, n29135, n2995, n29337, n2996, n29336, 
        n27862, n2109, n43638, n29134, n2997, n29335, n2998, n29334, 
        n2999, n29333, n3000, n29332, n3001, n29331, n3002, n29330, 
        n29133, n29132, n27861, n27860, n3003, n29329, n3004, 
        n29328, n3005, n29327, n29131, n3006, n29326, n27859, 
        n3007, n29325, n29130, n3008, n29324, n3009, n29323, n29129, 
        n29322, n29128, n29321, n27858, n29127, n14, n13, n14_adj_4532, 
        n15, n16, n22_adj_4533, n37594, n20, n24, n15841;
    wire [31:0]one_wire_N_513;
    
    wire n30047, n24922, n4, n13_adj_4534, n15961, n15776, n24962, 
        n24_adj_4535, n34_adj_4536, n22_adj_4537, n38_adj_4538, n36, 
        n37_adj_4539, n35_adj_4540, n18_adj_4541, n17, n19, n27857, 
        n21, n23, n22_adj_4542, n24_adj_4543, n36_adj_4544, n25_adj_4545, 
        n27_adj_4546, n26_adj_4547, n28_adj_4548, n37_adj_4549, n29, 
        n30_adj_4550, n34976, n35738, n30206, n24698, n35021, n116, 
        n29320, n29126, n27856, n29319, n29125, n29318, n29124, 
        n29317, n29123, n29122, n29316, n29121, n29315, n29120, 
        n29314, n29119, n29313, n43640, n29118, n29312, n29311, 
        n1895, n1928, n29117, n29310, n1896, n29116, n29309, n1897, 
        n29115, n29308, n1898, n29114, n1899, n29113, n27855, 
        n29307, n29306, n1900, n29112, n29305, n29304, n36_adj_4551, 
        n1901, n29111, n29303, n29302, n1902, n29110, n25_adj_4552, 
        n1903, n29109, n29301, n1904, n29108, n29300, n1905, n29107, 
        n27854, n34_adj_4553, n40_adj_4554, n29299, n1906, n29106, 
        n27853, n35682, n14452, n807, n838, n35829, n1907, n29105, 
        n24982, n35706, n24488, n43641, n29298, \neo_pixel_transmitter.done_N_576 , 
        n17155, n1908, n29104, n1909, n43642, n29103, n27852, 
        n2786, n2819, n29297, n2787, n29296, n1796, n1829, n29102, 
        n1797, n29101, n2788, n29295, n1798, n29100, n2789, n29294, 
        n1799, n29099, n2790, n29293, n1800, n29098, n2791, n29292, 
        n40_adj_4555, n44, n42, n1801, n29097, n43_adj_4556, n41_adj_4557, 
        n38_adj_4558, n46_adj_4559, n50, n37_adj_4560, n38_adj_4561, 
        n1802, n29096, n39_adj_4562, n37_adj_4563, n1803, n29095, 
        n2792, n29291, n2793, n29290, n1804, n29094;
    wire [31:0]n971;
    
    wire n905, n28245, n906, n28244, n28243, n17296, n28242, n14450, 
        n28241, n1103, n4_adj_4564, n1037, n28240, n1104, n1005, 
        n28239, n2794, n29289, n1805, n29093, n1105, n1006, n28238, 
        n2795, n29288, n1806, n29092, n1106, n1007, n28237, n1807, 
        n29091, n1107, n1008, n28236, n1108, n1009, n43645, n28235, 
        n1109, n2796, n29287, n1808, n29090, n2797, n29286, n1809, 
        n43644, n29089, n1202, n1136, n28234, n1203, n28233, n1204, 
        n28232, n1205, n28231, n1206, n28230, n1207, n28229, n2798, 
        n29285, n1697, n1730, n29088, n1208, n43646, n28228, n1698, 
        n29087, n1209, n2799, n29284, n1699, n29086, n27851, n1301, 
        n1235, n28221, n1302, n28220, n1303, n28219, n1304, n28218, 
        n1305, n28217, n1306, n28216, n1307, n28215, n2800, n29283, 
        n1308, n43648, n28214, n27850, n1309, n1700, n29085, n2801, 
        n29282, n1701, n29084, n2802, n29281, n1702, n29083, n1703, 
        n29082, n2803, n29280, n2804, n29279, n1704, n29081, n2805, 
        n29278, n1705, n29080, n27849, n2806, n29277, n1706, n29079, 
        n1707, n29078, n2807, n29276, n27848, n1708, n29077, n27847, 
        n2808, n29275, n1709, n43647, n29076, n18_adj_4565, n24876, 
        n1400, n1334, n28204, n2809, n43643, n29274, n27846, n1631, 
        n29075, n1401, n28203, n1402, n28202, n29074, n30_adj_4566, 
        n27845, n27844, n2687, n2720, n29273, n29073, n1403, n28201, 
        n28_adj_4567, n2688, n29272, n29072, n27843, n1404, n28200, 
        n2689, n29271, n1405, n28199, n29071, n2690, n29270, n1406, 
        n28198, n29070, n29069, n27842, n2691, n29269, n2692, 
        n29268, n29068, n1407, n28197, n27841, n2693, n29267, 
        n29_adj_4568, n1408, n43649, n28196, n1409, n29067, n29066, 
        n2694, n29266, n29065, n2695, n29265, n43650, n29064, 
        n2696, n29264, n27_adj_4569, n2697, n29263, n2698, n29262, 
        n2699, n29261, n2700, n29260, n2701, n29259, n2702, n29258, 
        n29257, n29256, n29255, n29254, n1433, n28132, n28131, 
        n28130, n28129, n29253, n28128, n28127, n28126, n28125, 
        n29252, n28124, n43652, n28123, n43651, n29251, n29250, 
        n29249;
    wire [31:0]n1;
    
    wire n28100, n28099, n28098, n29248, n28097, n28096, n28095, 
        n28094, n29247, n28093, n28092, n28091, n28090, n28089, 
        n28088, n28087, n28086, n28085, n28084, n29246, n28083, 
        n28082, n29245, n28081, n28080, n28079, n28078, n28077, 
        n28076, n28075, n29244, n28074, n28073, n29243, n28072, 
        n28071, n28070, n4_adj_4592, n29242, n29241, n29240, n29239, 
        n29238, n29237, n28_adj_4594, n32_adj_4595, n30_adj_4596, 
        n31_adj_4597, n29_adj_4598, n36198, n35720, n36_adj_4599, 
        n46_adj_4600, n42_adj_4601, n34_adj_4602, n43_adj_4603, n50_adj_4604, 
        n48, n49, n47_adj_4605, n24567, n16_adj_4606, n17_adj_4607, 
        n708, n28_adj_4608, n38_adj_4609, n24904, n36_adj_4610, n42_adj_4611, 
        n40_adj_4612, n41_adj_4613, n39_adj_4614, n20_adj_4615, n13_adj_4616, 
        n18_adj_4617, n22_adj_4618, n10_adj_4619, n12_adj_4620, n16_adj_4621, 
        n14_adj_4622, n9_adj_4623, n17_adj_4624, n21_adj_4625, n20_adj_4626, 
        n24_adj_4627, n24800, n12_adj_4628, n31409, n38528, n38573, 
        n6_adj_4629, n60, n608, n35702, n13425, n24840, n18_adj_4630, 
        n24_adj_4631, n22_adj_4632, n26_adj_4633, n40_adj_4634, n38_adj_4635, 
        n39_adj_4636, n35879, n37_adj_4637, n34_adj_4638, n42_adj_4639, 
        n46_adj_4640, n33_adj_4641, n35847, n24747, n103, n34897, 
        n24770, n28_adj_4642, n26_adj_4643, n27_adj_4644, n25_adj_4645, 
        n20_adj_4646, n19_adj_4647, n37402, n21_adj_4648, n1167, n26_adj_4649, 
        n19_adj_4650, n16_adj_4651, n24_adj_4652, n28_adj_4653, n36438;
    
    SB_CARRY mod_5_add_1808_9 (.CI(n29235), .I0(n2603), .I1(n2621), .CO(n29236));
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n29234), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(clk32MHz), .E(n37672), .D(\neo_pixel_transmitter.done_N_570 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i34214_2_lut (.I0(\state_3__N_362[1] ), .I1(\state[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n40674));
    defparam i34214_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mod_5_add_1808_8 (.CI(n29234), .I0(n2604), .I1(n2621), .CO(n29235));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n29233), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_7 (.CI(n29233), .I0(n2605), .I1(n2621), .CO(n29234));
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n29232), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_6 (.CI(n29232), .I0(n2606), .I1(n2621), .CO(n29233));
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n29231), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1499), .I1(n1499), .I2(n1532), 
            .I3(n27952), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_5 (.CI(n29231), .I0(n2607), .I1(n2621), .CO(n29232));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n29230), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_4 (.CI(n29230), .I0(n2608), .I1(n2621), .CO(n29231));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n43630), 
            .I3(n29229), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_3 (.CI(n29229), .I0(n2609), .I1(n43630), .CO(n29230));
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n43630), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1071_12_lut (.I0(n1500), .I1(n1500), .I2(n1532), 
            .I3(n27951), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_12 (.CI(n27951), .I0(n1500), .I1(n1532), .CO(n27952));
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n43630), 
            .CO(n29229));
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2489), .I1(n2489), .I2(n2522), 
            .I3(n29228), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_11_lut (.I0(n1501), .I1(n1501), .I2(n1532), 
            .I3(n27950), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(n2490), .I1(n2490), .I2(n2522), 
            .I3(n29227), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_22 (.CI(n29227), .I0(n2490), .I1(n2522), .CO(n29228));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(n2491), .I1(n2491), .I2(n2522), 
            .I3(n29226), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_21 (.CI(n29226), .I0(n2491), .I1(n2522), .CO(n29227));
    SB_CARRY mod_5_add_1071_11 (.CI(n27950), .I0(n1501), .I1(n1532), .CO(n27951));
    SB_LUT4 mod_5_add_1071_10_lut (.I0(n1502), .I1(n1502), .I2(n1532), 
            .I3(n27949), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_10 (.CI(n27949), .I0(n1502), .I1(n1532), .CO(n27950));
    SB_DFF bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(clk32MHz), .D(n33653));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(clk32MHz), .D(n33655));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(clk32MHz), .D(n33657));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(clk32MHz), .D(n33659));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(clk32MHz), .D(n33661));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(clk32MHz), .D(n33663));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(clk32MHz), .D(n33665));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(clk32MHz), .D(n33635));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(clk32MHz), .D(n33639));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(clk32MHz), .D(n33641));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(clk32MHz), .D(n33643));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(clk32MHz), .D(n33645));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(clk32MHz), .D(n33647));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(clk32MHz), .D(n18307));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(clk32MHz), .E(VCC_net), 
            .D(n33589));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(clk32MHz), .D(n33673));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(clk32MHz), .D(n33623));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(clk32MHz), .D(n33667));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(clk32MHz), .D(n33669));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(clk32MHz), .D(n33671));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(clk32MHz), .D(n33649));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(clk32MHz), .D(n33651));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(clk32MHz), .D(n33631));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(clk32MHz), .D(n33633));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(clk32MHz), .E(VCC_net), 
            .D(n33595));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(clk32MHz), .D(n18212));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(clk32MHz), .E(VCC_net), 
            .D(n33601));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(clk32MHz), .D(n33621));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i8_3_lut (.I0(bit_ctr[6]), .I1(n2907), .I2(n2909), .I3(GND_net), 
            .O(n33));
    defparam i8_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i16_4_lut (.I0(n2900), .I1(n2891), .I2(n2897), .I3(n2888), 
            .O(n41));
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n2906), .I1(n2887), .I2(n2892), .I3(GND_net), 
            .O(n38));
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut (.I0(n2896), .I1(n2885), .I2(n2905), .I3(n2902), 
            .O(n43));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1071_9_lut (.I0(n1503), .I1(n1503), .I2(n1532), 
            .I3(n27948), .O(n1602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i15_4_lut (.I0(n2899), .I1(n2890), .I2(n2898), .I3(n2908), 
            .O(n40));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut (.I0(n41), .I1(n33), .I2(n2889), .I3(n2901), .O(n46));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n2886), .I1(n2894), .I2(n2895), .I3(n2903), 
            .O(n39));
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut (.I0(n43), .I1(n2904), .I2(n38), .I3(n2893), .O(n47));
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n47), .I1(n39), .I2(n46), .I3(n40), .O(n2918));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1071_9 (.CI(n27948), .I0(n1503), .I1(n1532), .CO(n27949));
    SB_LUT4 mod_5_add_1071_8_lut (.I0(n1504), .I1(n1504), .I2(n1532), 
            .I3(n27947), .O(n1603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i7_3_lut (.I0(bit_ctr[11]), .I1(n2401), .I2(n2409), .I3(GND_net), 
            .O(n27));
    defparam i7_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i13_4_lut (.I0(n2390), .I1(n2391), .I2(n2397), .I3(n2407), 
            .O(n33_adj_4527));
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(n2405), .I1(n2394), .I2(n2400), .I3(n2399), 
            .O(n32));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n2406), .I1(n2396), .I2(n2403), .I3(n2402), 
            .O(n31));
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1600 (.I0(n2393), .I1(n2392), .I2(n2408), .I3(n2398), 
            .O(n35));
    defparam i15_4_lut_adj_1600.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(n33_adj_4527), .I1(n27), .I2(n2404), .I3(n2395), 
            .O(n37));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(n37), .I1(n35), .I2(n31), .I3(n32), .O(n2423));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1741_20_lut (.I0(n2492), .I1(n2492), .I2(n2522), 
            .I3(n29225), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i3_2_lut (.I0(n2302), .I1(n2292), .I2(GND_net), .I3(GND_net), 
            .O(n22));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY mod_5_add_1071_8 (.CI(n27947), .I0(n1504), .I1(n1532), .CO(n27948));
    SB_LUT4 mod_5_add_1071_7_lut (.I0(n1505), .I1(n1505), .I2(n1532), 
            .I3(n27946), .O(n1604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i11_4_lut_adj_1601 (.I0(bit_ctr[12]), .I1(n22), .I2(n2299), 
            .I3(n2309), .O(n30));
    defparam i11_4_lut_adj_1601.LUT_INIT = 16'hfefc;
    SB_LUT4 i36787_1_lut (.I0(n2522), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43632));
    defparam i36787_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36794_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43639));
    defparam i36794_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15_4_lut_adj_1602 (.I0(n2294), .I1(n30), .I2(n2306), .I3(n2297), 
            .O(n34));
    defparam i15_4_lut_adj_1602.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1603 (.I0(n2301), .I1(n2307), .I2(n2291), .I3(n2305), 
            .O(n32_adj_4528));
    defparam i13_4_lut_adj_1603.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1741_20 (.CI(n29225), .I0(n2492), .I1(n2522), .CO(n29226));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(n2493), .I1(n2493), .I2(n2522), 
            .I3(n29224), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i14_4_lut_adj_1604 (.I0(n2298), .I1(n2295), .I2(n2304), .I3(n2300), 
            .O(n33_adj_4529));
    defparam i14_4_lut_adj_1604.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1741_19 (.CI(n29224), .I0(n2493), .I1(n2522), .CO(n29225));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(n2494), .I1(n2494), .I2(n2522), 
            .I3(n29223), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i12_4_lut_adj_1605 (.I0(n2308), .I1(n2296), .I2(n2303), .I3(n2293), 
            .O(n31_adj_4530));
    defparam i12_4_lut_adj_1605.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1606 (.I0(n31_adj_4530), .I1(n33_adj_4529), .I2(n32_adj_4528), 
            .I3(n34), .O(n2324));
    defparam i18_4_lut_adj_1606.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1741_18 (.CI(n29223), .I0(n2494), .I1(n2522), .CO(n29224));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(n2495), .I1(n2495), .I2(n2522), 
            .I3(n29222), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_17 (.CI(n29222), .I0(n2495), .I1(n2522), .CO(n29223));
    SB_CARRY mod_5_add_1071_7 (.CI(n27946), .I0(n1505), .I1(n1532), .CO(n27947));
    SB_LUT4 i36788_1_lut (.I0(n2423), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43633));
    defparam i36788_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1071_6_lut (.I0(n1506), .I1(n1506), .I2(n1532), 
            .I3(n27945), .O(n1605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_6 (.CI(n27945), .I0(n1506), .I1(n1532), .CO(n27946));
    SB_LUT4 mod_5_add_1071_5_lut (.I0(n1507), .I1(n1507), .I2(n1532), 
            .I3(n27944), .O(n1606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_5 (.CI(n27944), .I0(n1507), .I1(n1532), .CO(n27945));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(n2496), .I1(n2496), .I2(n2522), 
            .I3(n29221), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_4_lut (.I0(n1508), .I1(n1508), .I2(n1532), 
            .I3(n27943), .O(n1607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_4 (.CI(n27943), .I0(n1508), .I1(n1532), .CO(n27944));
    SB_CARRY mod_5_add_1741_16 (.CI(n29221), .I0(n2496), .I1(n2522), .CO(n29222));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(n2497), .I1(n2497), .I2(n2522), 
            .I3(n29220), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_15 (.CI(n29220), .I0(n2497), .I1(n2522), .CO(n29221));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(n2498), .I1(n2498), .I2(n2522), 
            .I3(n29219), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_14 (.CI(n29219), .I0(n2498), .I1(n2522), .CO(n29220));
    SB_LUT4 mod_5_add_1741_13_lut (.I0(n2499), .I1(n2499), .I2(n2522), 
            .I3(n29218), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_3_lut (.I0(n1509), .I1(n1509), .I2(n43631), 
            .I3(n27942), .O(n1608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1741_13 (.CI(n29218), .I0(n2499), .I1(n2522), .CO(n29219));
    SB_CARRY mod_5_add_1071_3 (.CI(n27942), .I0(n1509), .I1(n43631), .CO(n27943));
    SB_LUT4 mod_5_add_1741_12_lut (.I0(n2500), .I1(n2500), .I2(n2522), 
            .I3(n29217), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_12 (.CI(n29217), .I0(n2500), .I1(n2522), .CO(n29218));
    SB_LUT4 mod_5_add_1741_11_lut (.I0(n2501), .I1(n2501), .I2(n2522), 
            .I3(n29216), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_11 (.CI(n29216), .I0(n2501), .I1(n2522), .CO(n29217));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(n2502), .I1(n2502), .I2(n2522), 
            .I3(n29215), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_10 (.CI(n29215), .I0(n2502), .I1(n2522), .CO(n29216));
    SB_LUT4 mod_5_add_1741_9_lut (.I0(n2503), .I1(n2503), .I2(n2522), 
            .I3(n29214), .O(n2602)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_9 (.CI(n29214), .I0(n2503), .I1(n2522), .CO(n29215));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(n2504), .I1(n2504), .I2(n2522), 
            .I3(n29213), .O(n2603)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1741_8 (.CI(n29213), .I0(n2504), .I1(n2522), .CO(n29214));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(bit_ctr[20]), .I1(bit_ctr[20]), .I2(n43631), 
            .I3(VCC_net), .O(n1609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 timer_1223_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n28601), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(n43631), 
            .CO(n27942));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(n2505), .I1(n2505), .I2(n2522), 
            .I3(n29212), .O(n2604)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1223_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n28600), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_7 (.CI(n29212), .I0(n2505), .I1(n2522), .CO(n29213));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(n2506), .I1(n2506), .I2(n2522), 
            .I3(n29211), .O(n2605)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1223_add_4_32 (.CI(n28600), .I0(GND_net), .I1(timer[30]), 
            .CO(n28601));
    SB_CARRY mod_5_add_1741_6 (.CI(n29211), .I0(n2506), .I1(n2522), .CO(n29212));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(n2507), .I1(n2507), .I2(n2522), 
            .I3(n29210), .O(n2606)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1223_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n28599), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_5 (.CI(n29210), .I0(n2507), .I1(n2522), .CO(n29211));
    SB_CARRY timer_1223_add_4_31 (.CI(n28599), .I0(GND_net), .I1(timer[29]), 
            .CO(n28600));
    SB_LUT4 timer_1223_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n28598), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_4_lut (.I0(n2508), .I1(n2508), .I2(n2522), 
            .I3(n29209), .O(n2607)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1223_add_4_30 (.CI(n28598), .I0(GND_net), .I1(timer[28]), 
            .CO(n28599));
    SB_LUT4 timer_1223_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n28597), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_29 (.CI(n28597), .I0(GND_net), .I1(timer[27]), 
            .CO(n28598));
    SB_LUT4 timer_1223_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n28596), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_28 (.CI(n28596), .I0(GND_net), .I1(timer[26]), 
            .CO(n28597));
    SB_LUT4 timer_1223_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n28595), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_27 (.CI(n28595), .I0(GND_net), .I1(timer[25]), 
            .CO(n28596));
    SB_CARRY mod_5_add_1741_4 (.CI(n29209), .I0(n2508), .I1(n2522), .CO(n29210));
    SB_LUT4 timer_1223_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n28594), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_26 (.CI(n28594), .I0(GND_net), .I1(timer[24]), 
            .CO(n28595));
    SB_LUT4 timer_1223_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n28593), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_25 (.CI(n28593), .I0(GND_net), .I1(timer[23]), 
            .CO(n28594));
    SB_LUT4 timer_1223_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n28592), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_3_lut (.I0(n2509), .I1(n2509), .I2(n43632), 
            .I3(n29208), .O(n2608)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY timer_1223_add_4_24 (.CI(n28592), .I0(GND_net), .I1(timer[22]), 
            .CO(n28593));
    SB_LUT4 timer_1223_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n28591), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_23 (.CI(n28591), .I0(GND_net), .I1(timer[21]), 
            .CO(n28592));
    SB_LUT4 timer_1223_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n28590), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_22 (.CI(n28590), .I0(GND_net), .I1(timer[20]), 
            .CO(n28591));
    SB_LUT4 timer_1223_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n28589), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_21 (.CI(n28589), .I0(GND_net), .I1(timer[19]), 
            .CO(n28590));
    SB_CARRY mod_5_add_1741_3 (.CI(n29208), .I0(n2509), .I1(n43632), .CO(n29209));
    SB_LUT4 timer_1223_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n28588), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_20 (.CI(n28588), .I0(GND_net), .I1(timer[18]), 
            .CO(n28589));
    SB_LUT4 timer_1223_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n28587), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_19 (.CI(n28587), .I0(GND_net), .I1(timer[17]), 
            .CO(n28588));
    SB_LUT4 timer_1223_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n28586), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_18 (.CI(n28586), .I0(GND_net), .I1(timer[16]), 
            .CO(n28587));
    SB_LUT4 timer_1223_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n28585), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_17 (.CI(n28585), .I0(GND_net), .I1(timer[15]), 
            .CO(n28586));
    SB_LUT4 timer_1223_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n28584), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_16 (.CI(n28584), .I0(GND_net), .I1(timer[14]), 
            .CO(n28585));
    SB_LUT4 timer_1223_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n28583), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_2_lut (.I0(bit_ctr[10]), .I1(bit_ctr[10]), .I2(n43632), 
            .I3(VCC_net), .O(n2609)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY timer_1223_add_4_15 (.CI(n28583), .I0(GND_net), .I1(timer[13]), 
            .CO(n28584));
    SB_LUT4 timer_1223_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n28582), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_14 (.CI(n28582), .I0(GND_net), .I1(timer[12]), 
            .CO(n28583));
    SB_LUT4 timer_1223_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n28581), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_13 (.CI(n28581), .I0(GND_net), .I1(timer[11]), 
            .CO(n28582));
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(n43632), 
            .CO(n29208));
    SB_LUT4 timer_1223_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n28580), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2390), .I1(n2390), .I2(n2423), 
            .I3(n29207), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1223_add_4_12 (.CI(n28580), .I0(GND_net), .I1(timer[10]), 
            .CO(n28581));
    SB_LUT4 mod_5_add_1674_21_lut (.I0(n2391), .I1(n2391), .I2(n2423), 
            .I3(n29206), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_21 (.CI(n29206), .I0(n2391), .I1(n2423), .CO(n29207));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(n2392), .I1(n2392), .I2(n2423), 
            .I3(n29205), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1223_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n28579), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_11 (.CI(n28579), .I0(GND_net), .I1(timer[9]), 
            .CO(n28580));
    SB_LUT4 timer_1223_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n28578), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_20 (.CI(n29205), .I0(n2392), .I1(n2423), .CO(n29206));
    SB_CARRY timer_1223_add_4_10 (.CI(n28578), .I0(GND_net), .I1(timer[8]), 
            .CO(n28579));
    SB_LUT4 timer_1223_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n28577), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_19_lut (.I0(n2393), .I1(n2393), .I2(n2423), 
            .I3(n29204), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_19 (.CI(n29204), .I0(n2393), .I1(n2423), .CO(n29205));
    SB_CARRY timer_1223_add_4_9 (.CI(n28577), .I0(GND_net), .I1(timer[7]), 
            .CO(n28578));
    SB_LUT4 timer_1223_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n28576), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_8 (.CI(n28576), .I0(GND_net), .I1(timer[6]), 
            .CO(n28577));
    SB_LUT4 timer_1223_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n28575), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_18_lut (.I0(n2394), .I1(n2394), .I2(n2423), 
            .I3(n29203), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1223_add_4_7 (.CI(n28575), .I0(GND_net), .I1(timer[5]), 
            .CO(n28576));
    SB_CARRY mod_5_add_1674_18 (.CI(n29203), .I0(n2394), .I1(n2423), .CO(n29204));
    SB_LUT4 timer_1223_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n28574), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_6 (.CI(n28574), .I0(GND_net), .I1(timer[4]), 
            .CO(n28575));
    SB_LUT4 timer_1223_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n28573), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_5 (.CI(n28573), .I0(GND_net), .I1(timer[3]), 
            .CO(n28574));
    SB_LUT4 timer_1223_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n28572), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1674_17_lut (.I0(n2395), .I1(n2395), .I2(n2423), 
            .I3(n29202), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1223_add_4_4 (.CI(n28572), .I0(GND_net), .I1(timer[2]), 
            .CO(n28573));
    SB_CARRY mod_5_add_1674_17 (.CI(n29202), .I0(n2395), .I1(n2423), .CO(n29203));
    SB_LUT4 timer_1223_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n28571), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36786_1_lut (.I0(n1532), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43631));
    defparam i36786_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1674_16_lut (.I0(n2396), .I1(n2396), .I2(n2423), 
            .I3(n29201), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY timer_1223_add_4_3 (.CI(n28571), .I0(GND_net), .I1(timer[1]), 
            .CO(n28572));
    SB_LUT4 timer_1223_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1223_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1223_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n28571));
    SB_CARRY mod_5_add_1674_16 (.CI(n29201), .I0(n2396), .I1(n2423), .CO(n29202));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(n2397), .I1(n2397), .I2(n2423), 
            .I3(n29200), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_15 (.CI(n29200), .I0(n2397), .I1(n2423), .CO(n29201));
    SB_LUT4 mod_5_add_1674_14_lut (.I0(n2398), .I1(n2398), .I2(n2423), 
            .I3(n29199), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_14 (.CI(n29199), .I0(n2398), .I1(n2423), .CO(n29200));
    SB_LUT4 mod_5_add_1674_13_lut (.I0(n2399), .I1(n2399), .I2(n2423), 
            .I3(n29198), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_13 (.CI(n29198), .I0(n2399), .I1(n2423), .CO(n29199));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(n2400), .I1(n2400), .I2(n2423), 
            .I3(n29197), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_12 (.CI(n29197), .I0(n2400), .I1(n2423), .CO(n29198));
    SB_LUT4 mod_5_add_1674_11_lut (.I0(n2401), .I1(n2401), .I2(n2423), 
            .I3(n29196), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_11 (.CI(n29196), .I0(n2401), .I1(n2423), .CO(n29197));
    SB_LUT4 add_21_33_lut (.I0(n25779), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(n27871), .O(n40726)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_32_lut (.I0(n25779), .I1(bit_ctr[30]), .I2(GND_net), 
            .I3(n27870), .O(n40725)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1674_10_lut (.I0(n2402), .I1(n2402), .I2(n2423), 
            .I3(n29195), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_32 (.CI(n27870), .I0(bit_ctr[30]), .I1(GND_net), .CO(n27871));
    SB_CARRY mod_5_add_1674_10 (.CI(n29195), .I0(n2402), .I1(n2423), .CO(n29196));
    SB_LUT4 mod_5_add_1674_9_lut (.I0(n2403), .I1(n2403), .I2(n2423), 
            .I3(n29194), .O(n2502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_9 (.CI(n29194), .I0(n2403), .I1(n2423), .CO(n29195));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(n2404), .I1(n2404), .I2(n2423), 
            .I3(n29193), .O(n2503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_8 (.CI(n29193), .I0(n2404), .I1(n2423), .CO(n29194));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(n2405), .I1(n2405), .I2(n2423), 
            .I3(n29192), .O(n2504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_7 (.CI(n29192), .I0(n2405), .I1(n2423), .CO(n29193));
    SB_LUT4 add_21_31_lut (.I0(n25779), .I1(bit_ctr[29]), .I2(GND_net), 
            .I3(n27869), .O(n40724)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1674_6_lut (.I0(n2406), .I1(n2406), .I2(n2423), 
            .I3(n29191), .O(n2505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_6 (.CI(n29191), .I0(n2406), .I1(n2423), .CO(n29192));
    SB_LUT4 mod_5_add_1674_5_lut (.I0(n2407), .I1(n2407), .I2(n2423), 
            .I3(n29190), .O(n2506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_5 (.CI(n29190), .I0(n2407), .I1(n2423), .CO(n29191));
    SB_LUT4 mod_5_add_1674_4_lut (.I0(n2408), .I1(n2408), .I2(n2423), 
            .I3(n29189), .O(n2507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_31 (.CI(n27869), .I0(bit_ctr[29]), .I1(GND_net), .CO(n27870));
    SB_CARRY mod_5_add_1674_4 (.CI(n29189), .I0(n2408), .I1(n2423), .CO(n29190));
    SB_LUT4 mod_5_add_1674_3_lut (.I0(n2409), .I1(n2409), .I2(n43633), 
            .I3(n29188), .O(n2508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_30_lut (.I0(n25779), .I1(bit_ctr[28]), .I2(GND_net), 
            .I3(n27868), .O(n40723)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1674_3 (.CI(n29188), .I0(n2409), .I1(n43633), .CO(n29189));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(bit_ctr[11]), .I1(bit_ctr[11]), .I2(n43633), 
            .I3(VCC_net), .O(n2509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(n43633), 
            .CO(n29188));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2291), .I1(n2291), .I2(n2324), 
            .I3(n29187), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(n2292), .I1(n2292), .I2(n2324), 
            .I3(n29186), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_30 (.CI(n27868), .I0(bit_ctr[28]), .I1(GND_net), .CO(n27869));
    SB_CARRY mod_5_add_1607_20 (.CI(n29186), .I0(n2292), .I1(n2324), .CO(n29187));
    SB_LUT4 mod_5_add_1607_19_lut (.I0(n2293), .I1(n2293), .I2(n2324), 
            .I3(n29185), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_19 (.CI(n29185), .I0(n2293), .I1(n2324), .CO(n29186));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(n2294), .I1(n2294), .I2(n2324), 
            .I3(n29184), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_18 (.CI(n29184), .I0(n2294), .I1(n2324), .CO(n29185));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(n2295), .I1(n2295), .I2(n2324), 
            .I3(n29183), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_17 (.CI(n29183), .I0(n2295), .I1(n2324), .CO(n29184));
    SB_LUT4 mod_5_add_1607_16_lut (.I0(n2296), .I1(n2296), .I2(n2324), 
            .I3(n29182), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_16 (.CI(n29182), .I0(n2296), .I1(n2324), .CO(n29183));
    SB_LUT4 mod_5_add_1607_15_lut (.I0(n2297), .I1(n2297), .I2(n2324), 
            .I3(n29181), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_15 (.CI(n29181), .I0(n2297), .I1(n2324), .CO(n29182));
    SB_LUT4 mod_5_add_1607_14_lut (.I0(n2298), .I1(n2298), .I2(n2324), 
            .I3(n29180), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_14 (.CI(n29180), .I0(n2298), .I1(n2324), .CO(n29181));
    SB_LUT4 add_21_29_lut (.I0(n25779), .I1(bit_ctr[27]), .I2(GND_net), 
            .I3(n27867), .O(n40722)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1607_13_lut (.I0(n2299), .I1(n2299), .I2(n2324), 
            .I3(n29179), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_13 (.CI(n29179), .I0(n2299), .I1(n2324), .CO(n29180));
    SB_LUT4 mod_5_add_1607_12_lut (.I0(n2300), .I1(n2300), .I2(n2324), 
            .I3(n29178), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_12 (.CI(n29178), .I0(n2300), .I1(n2324), .CO(n29179));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(n2301), .I1(n2301), .I2(n2324), 
            .I3(n29177), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_29 (.CI(n27867), .I0(bit_ctr[27]), .I1(GND_net), .CO(n27868));
    SB_CARRY mod_5_add_1607_11 (.CI(n29177), .I0(n2301), .I1(n2324), .CO(n29178));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(n2302), .I1(n2302), .I2(n2324), 
            .I3(n29176), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_10 (.CI(n29176), .I0(n2302), .I1(n2324), .CO(n29177));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(n2303), .I1(n2303), .I2(n2324), 
            .I3(n29175), .O(n2402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_9 (.CI(n29175), .I0(n2303), .I1(n2324), .CO(n29176));
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3083), .I1(n3083), .I2(n3116), 
            .I3(n29375), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_28_lut (.I0(n25779), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(n27866), .O(n40721)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1607_8_lut (.I0(n2304), .I1(n2304), .I2(n2324), 
            .I3(n29174), .O(n2403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(n3084), .I1(n3084), .I2(n3116), 
            .I3(n29374), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_8 (.CI(n29174), .I0(n2304), .I1(n2324), .CO(n29175));
    SB_LUT4 mod_5_add_1607_7_lut (.I0(n2305), .I1(n2305), .I2(n2324), 
            .I3(n29173), .O(n2404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_28 (.CI(n29374), .I0(n3084), .I1(n3116), .CO(n29375));
    SB_CARRY mod_5_add_1607_7 (.CI(n29173), .I0(n2305), .I1(n2324), .CO(n29174));
    SB_LUT4 mod_5_add_2143_27_lut (.I0(n3085), .I1(n3085), .I2(n3116), 
            .I3(n29373), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_27 (.CI(n29373), .I0(n3085), .I1(n3116), .CO(n29374));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(n2306), .I1(n2306), .I2(n2324), 
            .I3(n29172), .O(n2405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_26_lut (.I0(n3086), .I1(n3086), .I2(n3116), 
            .I3(n29372), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_26 (.CI(n29372), .I0(n3086), .I1(n3116), .CO(n29373));
    SB_CARRY add_21_28 (.CI(n27866), .I0(bit_ctr[26]), .I1(GND_net), .CO(n27867));
    SB_CARRY mod_5_add_1607_6 (.CI(n29172), .I0(n2306), .I1(n2324), .CO(n29173));
    SB_LUT4 mod_5_add_1607_5_lut (.I0(n2307), .I1(n2307), .I2(n2324), 
            .I3(n29171), .O(n2406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_25_lut (.I0(n3087), .I1(n3087), .I2(n3116), 
            .I3(n29371), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_5 (.CI(n29171), .I0(n2307), .I1(n2324), .CO(n29172));
    SB_CARRY mod_5_add_2143_25 (.CI(n29371), .I0(n3087), .I1(n3116), .CO(n29372));
    SB_LUT4 mod_5_add_2143_24_lut (.I0(n3088), .I1(n3088), .I2(n3116), 
            .I3(n29370), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_24 (.CI(n29370), .I0(n3088), .I1(n3116), .CO(n29371));
    SB_LUT4 mod_5_add_2143_23_lut (.I0(n3089), .I1(n3089), .I2(n3116), 
            .I3(n29369), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_4_lut (.I0(n2308), .I1(n2308), .I2(n2324), 
            .I3(n29170), .O(n2407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_23 (.CI(n29369), .I0(n3089), .I1(n3116), .CO(n29370));
    SB_CARRY mod_5_add_1607_4 (.CI(n29170), .I0(n2308), .I1(n2324), .CO(n29171));
    SB_LUT4 mod_5_add_2143_22_lut (.I0(n3090), .I1(n3090), .I2(n3116), 
            .I3(n29368), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_3_lut (.I0(n2309), .I1(n2309), .I2(n43634), 
            .I3(n29169), .O(n2408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_22 (.CI(n29368), .I0(n3090), .I1(n3116), .CO(n29369));
    SB_LUT4 mod_5_add_2143_21_lut (.I0(n3091), .I1(n3091), .I2(n3116), 
            .I3(n29367), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_3 (.CI(n29169), .I0(n2309), .I1(n43634), .CO(n29170));
    SB_LUT4 mod_5_add_1607_2_lut (.I0(bit_ctr[12]), .I1(bit_ctr[12]), .I2(n43634), 
            .I3(VCC_net), .O(n2409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_21 (.CI(n29367), .I0(n3091), .I1(n3116), .CO(n29368));
    SB_LUT4 mod_5_add_2143_20_lut (.I0(n3092), .I1(n3092), .I2(n3116), 
            .I3(n29366), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(n43634), 
            .CO(n29169));
    SB_CARRY mod_5_add_2143_20 (.CI(n29366), .I0(n3092), .I1(n3116), .CO(n29367));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(n3093), .I1(n3093), .I2(n3116), 
            .I3(n29365), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2192), .I1(n2192), .I2(n2225), 
            .I3(n29168), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_19 (.CI(n29365), .I0(n3093), .I1(n3116), .CO(n29366));
    SB_LUT4 mod_5_add_1540_19_lut (.I0(n2193), .I1(n2193), .I2(n2225), 
            .I3(n29167), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_27_lut (.I0(n25779), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(n27865), .O(n40720)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_27 (.CI(n27865), .I0(bit_ctr[25]), .I1(GND_net), .CO(n27866));
    SB_LUT4 i2_2_lut (.I0(n1998), .I1(n2004), .I2(GND_net), .I3(GND_net), 
            .O(n18));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1607 (.I0(n2003), .I1(n1999), .I2(n1996), .I3(n2007), 
            .O(n28));
    defparam i12_4_lut_adj_1607.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(n1997), .I1(n2005), .I2(n2000), .I3(n2002), 
            .O(n26));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1540_19 (.CI(n29167), .I0(n2193), .I1(n2225), .CO(n29168));
    SB_LUT4 i11_4_lut_adj_1608 (.I0(n2001), .I1(n2008), .I2(n1994), .I3(n1995), 
            .O(n27_adj_4531));
    defparam i11_4_lut_adj_1608.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(bit_ctr[15]), .I1(n18), .I2(n2006), .I3(n2009), 
            .O(n25));
    defparam i9_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 mod_5_add_2143_18_lut (.I0(n3094), .I1(n3094), .I2(n3116), 
            .I3(n29364), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_18_lut (.I0(n2194), .I1(n2194), .I2(n2225), 
            .I3(n29166), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_18 (.CI(n29364), .I0(n3094), .I1(n3116), .CO(n29365));
    SB_CARRY mod_5_add_1540_18 (.CI(n29166), .I0(n2194), .I1(n2225), .CO(n29167));
    SB_LUT4 i15_4_lut_adj_1609 (.I0(n25), .I1(n27_adj_4531), .I2(n26), 
            .I3(n28), .O(n2027));
    defparam i15_4_lut_adj_1609.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_17_lut (.I0(n2195), .I1(n2195), .I2(n2225), 
            .I3(n29165), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_26_lut (.I0(n25779), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(n27864), .O(n40719)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2143_17_lut (.I0(n3095), .I1(n3095), .I2(n3116), 
            .I3(n29363), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_17 (.CI(n29165), .I0(n2195), .I1(n2225), .CO(n29166));
    SB_LUT4 mod_5_add_1540_16_lut (.I0(n2196), .I1(n2196), .I2(n2225), 
            .I3(n29164), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_17 (.CI(n29363), .I0(n3095), .I1(n3116), .CO(n29364));
    SB_CARRY mod_5_add_1540_16 (.CI(n29164), .I0(n2196), .I1(n2225), .CO(n29165));
    SB_LUT4 mod_5_add_1540_15_lut (.I0(n2197), .I1(n2197), .I2(n2225), 
            .I3(n29163), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_15 (.CI(n29163), .I0(n2197), .I1(n2225), .CO(n29164));
    SB_LUT4 mod_5_add_2143_16_lut (.I0(n3096), .I1(n3096), .I2(n3116), 
            .I3(n29362), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_14_lut (.I0(n2198), .I1(n2198), .I2(n2225), 
            .I3(n29162), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_14 (.CI(n29162), .I0(n2198), .I1(n2225), .CO(n29163));
    SB_CARRY mod_5_add_2143_16 (.CI(n29362), .I0(n3096), .I1(n3116), .CO(n29363));
    SB_LUT4 mod_5_add_1540_13_lut (.I0(n2199), .I1(n2199), .I2(n2225), 
            .I3(n29161), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_15_lut (.I0(n3097), .I1(n3097), .I2(n3116), 
            .I3(n29361), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_13 (.CI(n29161), .I0(n2199), .I1(n2225), .CO(n29162));
    SB_CARRY mod_5_add_2143_15 (.CI(n29361), .I0(n3097), .I1(n3116), .CO(n29362));
    SB_LUT4 mod_5_add_1540_12_lut (.I0(n2200), .I1(n2200), .I2(n2225), 
            .I3(n29160), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_12 (.CI(n29160), .I0(n2200), .I1(n2225), .CO(n29161));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(n3098), .I1(n3098), .I2(n3116), 
            .I3(n29360), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_11_lut (.I0(n2201), .I1(n2201), .I2(n2225), 
            .I3(n29159), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_11 (.CI(n29159), .I0(n2201), .I1(n2225), .CO(n29160));
    SB_CARRY mod_5_add_2143_14 (.CI(n29360), .I0(n3098), .I1(n3116), .CO(n29361));
    SB_LUT4 mod_5_add_1540_10_lut (.I0(n2202), .I1(n2202), .I2(n2225), 
            .I3(n29158), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_10 (.CI(n29158), .I0(n2202), .I1(n2225), .CO(n29159));
    SB_LUT4 mod_5_add_1540_9_lut (.I0(n2203), .I1(n2203), .I2(n2225), 
            .I3(n29157), .O(n2302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_13_lut (.I0(n3099), .I1(n3099), .I2(n3116), 
            .I3(n29359), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_9 (.CI(n29157), .I0(n2203), .I1(n2225), .CO(n29158));
    SB_LUT4 mod_5_add_1540_8_lut (.I0(n2204), .I1(n2204), .I2(n2225), 
            .I3(n29156), .O(n2303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_13 (.CI(n29359), .I0(n3099), .I1(n3116), .CO(n29360));
    SB_CARRY mod_5_add_1540_8 (.CI(n29156), .I0(n2204), .I1(n2225), .CO(n29157));
    SB_LUT4 mod_5_add_1540_7_lut (.I0(n2205), .I1(n2205), .I2(n2225), 
            .I3(n29155), .O(n2304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_12_lut (.I0(n3100), .I1(n3100), .I2(n3116), 
            .I3(n29358), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_7 (.CI(n29155), .I0(n2205), .I1(n2225), .CO(n29156));
    SB_CARRY mod_5_add_2143_12 (.CI(n29358), .I0(n3100), .I1(n3116), .CO(n29359));
    SB_LUT4 mod_5_add_1540_6_lut (.I0(n2206), .I1(n2206), .I2(n2225), 
            .I3(n29154), .O(n2305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_11_lut (.I0(n3101), .I1(n3101), .I2(n3116), 
            .I3(n29357), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_6 (.CI(n29154), .I0(n2206), .I1(n2225), .CO(n29155));
    SB_LUT4 mod_5_add_1540_5_lut (.I0(n2207), .I1(n2207), .I2(n2225), 
            .I3(n29153), .O(n2306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_11 (.CI(n29357), .I0(n3101), .I1(n3116), .CO(n29358));
    SB_LUT4 mod_5_add_2143_10_lut (.I0(n3102), .I1(n3102), .I2(n3116), 
            .I3(n29356), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_10 (.CI(n29356), .I0(n3102), .I1(n3116), .CO(n29357));
    SB_CARRY mod_5_add_1540_5 (.CI(n29153), .I0(n2207), .I1(n2225), .CO(n29154));
    SB_LUT4 mod_5_add_1540_4_lut (.I0(n2208), .I1(n2208), .I2(n2225), 
            .I3(n29152), .O(n2307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2143_9_lut (.I0(n3103), .I1(n3103), .I2(n3116), 
            .I3(n29355), .O(n3202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1540_4 (.CI(n29152), .I0(n2208), .I1(n2225), .CO(n29153));
    SB_CARRY mod_5_add_2143_9 (.CI(n29355), .I0(n3103), .I1(n3116), .CO(n29356));
    SB_LUT4 mod_5_add_2143_8_lut (.I0(n3104), .I1(n3104), .I2(n3116), 
            .I3(n29354), .O(n3203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_3_lut (.I0(n2209), .I1(n2209), .I2(n43637), 
            .I3(n29151), .O(n2308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_8 (.CI(n29354), .I0(n3104), .I1(n3116), .CO(n29355));
    SB_CARRY mod_5_add_1540_3 (.CI(n29151), .I0(n2209), .I1(n43637), .CO(n29152));
    SB_LUT4 mod_5_add_2143_7_lut (.I0(n3105), .I1(n3105), .I2(n3116), 
            .I3(n29353), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_2_lut (.I0(bit_ctr[13]), .I1(bit_ctr[13]), .I2(n43637), 
            .I3(VCC_net), .O(n2309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_7 (.CI(n29353), .I0(n3105), .I1(n3116), .CO(n29354));
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(n43637), 
            .CO(n29151));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(n3106), .I1(n3106), .I2(n3116), 
            .I3(n29352), .O(n3205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2093), .I1(n2093), .I2(n2126), 
            .I3(n29150), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_6 (.CI(n29352), .I0(n3106), .I1(n3116), .CO(n29353));
    SB_LUT4 mod_5_add_2143_5_lut (.I0(n3107), .I1(n3107), .I2(n3116), 
            .I3(n29351), .O(n3206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_18_lut (.I0(n2094), .I1(n2094), .I2(n2126), 
            .I3(n29149), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_18 (.CI(n29149), .I0(n2094), .I1(n2126), .CO(n29150));
    SB_CARRY mod_5_add_2143_5 (.CI(n29351), .I0(n3107), .I1(n3116), .CO(n29352));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(n3108), .I1(n3108), .I2(n3116), 
            .I3(n29350), .O(n3207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_4 (.CI(n29350), .I0(n3108), .I1(n3116), .CO(n29351));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(n2095), .I1(n2095), .I2(n2126), 
            .I3(n29148), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_17 (.CI(n29148), .I0(n2095), .I1(n2126), .CO(n29149));
    SB_LUT4 mod_5_add_1473_16_lut (.I0(n2096), .I1(n2096), .I2(n2126), 
            .I3(n29147), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_16 (.CI(n29147), .I0(n2096), .I1(n2126), .CO(n29148));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(n3109), .I1(n3109), .I2(n43636), 
            .I3(n29349), .O(n3208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1473_15_lut (.I0(n2097), .I1(n2097), .I2(n2126), 
            .I3(n29146), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2143_3 (.CI(n29349), .I0(n3109), .I1(n43636), .CO(n29350));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(bit_ctr[4]), .I1(bit_ctr[4]), .I2(n43636), 
            .I3(VCC_net), .O(n3209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(n43636), 
            .CO(n29349));
    SB_CARRY mod_5_add_1473_15 (.CI(n29146), .I0(n2097), .I1(n2126), .CO(n29147));
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n29348), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_14_lut (.I0(n2098), .I1(n2098), .I2(n2126), 
            .I3(n29145), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_14 (.CI(n29145), .I0(n2098), .I1(n2126), .CO(n29146));
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n29347), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_13_lut (.I0(n2099), .I1(n2099), .I2(n2126), 
            .I3(n29144), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_27 (.CI(n29347), .I0(n2985), .I1(n3017), .CO(n29348));
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n29346), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_13 (.CI(n29144), .I0(n2099), .I1(n2126), .CO(n29145));
    SB_LUT4 mod_5_add_1473_12_lut (.I0(n2100), .I1(n2100), .I2(n2126), 
            .I3(n29143), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_26 (.CI(n29346), .I0(n2986), .I1(n3017), .CO(n29347));
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n29345), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_12 (.CI(n29143), .I0(n2100), .I1(n2126), .CO(n29144));
    SB_CARRY mod_5_add_2076_25 (.CI(n29345), .I0(n2987), .I1(n3017), .CO(n29346));
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n29344), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_11_lut (.I0(n2101), .I1(n2101), .I2(n2126), 
            .I3(n29142), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_11 (.CI(n29142), .I0(n2101), .I1(n2126), .CO(n29143));
    SB_LUT4 mod_5_add_1473_10_lut (.I0(n2102), .I1(n2102), .I2(n2126), 
            .I3(n29141), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_10 (.CI(n29141), .I0(n2102), .I1(n2126), .CO(n29142));
    SB_LUT4 mod_5_add_1473_9_lut (.I0(n2103), .I1(n2103), .I2(n2126), 
            .I3(n29140), .O(n2202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_24 (.CI(n29344), .I0(n2988), .I1(n3017), .CO(n29345));
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n29343), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_23 (.CI(n29343), .I0(n2989), .I1(n3017), .CO(n29344));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n29342), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_22 (.CI(n29342), .I0(n2990), .I1(n3017), .CO(n29343));
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n29341), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_9 (.CI(n29140), .I0(n2103), .I1(n2126), .CO(n29141));
    SB_CARRY mod_5_add_2076_21 (.CI(n29341), .I0(n2991), .I1(n3017), .CO(n29342));
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n29340), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_8_lut (.I0(n2104), .I1(n2104), .I2(n2126), 
            .I3(n29139), .O(n2203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_26 (.CI(n27864), .I0(bit_ctr[24]), .I1(GND_net), .CO(n27865));
    SB_CARRY mod_5_add_2076_20 (.CI(n29340), .I0(n2992), .I1(n3017), .CO(n29341));
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n29339), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_8 (.CI(n29139), .I0(n2104), .I1(n2126), .CO(n29140));
    SB_CARRY mod_5_add_2076_19 (.CI(n29339), .I0(n2993), .I1(n3017), .CO(n29340));
    SB_LUT4 mod_5_add_1473_7_lut (.I0(n2105), .I1(n2105), .I2(n2126), 
            .I3(n29138), .O(n2204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_25_lut (.I0(n25779), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(n27863), .O(n40718)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1473_7 (.CI(n29138), .I0(n2105), .I1(n2126), .CO(n29139));
    SB_LUT4 mod_5_add_1473_6_lut (.I0(n2106), .I1(n2106), .I2(n2126), 
            .I3(n29137), .O(n2205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n29338), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_18 (.CI(n29338), .I0(n2994), .I1(n3017), .CO(n29339));
    SB_CARRY mod_5_add_1473_6 (.CI(n29137), .I0(n2106), .I1(n2126), .CO(n29138));
    SB_CARRY add_21_25 (.CI(n27863), .I0(bit_ctr[23]), .I1(GND_net), .CO(n27864));
    SB_LUT4 mod_5_add_1473_5_lut (.I0(n2107), .I1(n2107), .I2(n2126), 
            .I3(n29136), .O(n2206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_5 (.CI(n29136), .I0(n2107), .I1(n2126), .CO(n29137));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(n2108), .I1(n2108), .I2(n2126), 
            .I3(n29135), .O(n2207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n29337), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1473_4 (.CI(n29135), .I0(n2108), .I1(n2126), .CO(n29136));
    SB_CARRY mod_5_add_2076_17 (.CI(n29337), .I0(n2995), .I1(n3017), .CO(n29338));
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n29336), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_24_lut (.I0(n25779), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(n27862), .O(n40717)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_2076_16 (.CI(n29336), .I0(n2996), .I1(n3017), .CO(n29337));
    SB_LUT4 mod_5_add_1473_3_lut (.I0(n2109), .I1(n2109), .I2(n43638), 
            .I3(n29134), .O(n2208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n29335), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_15 (.CI(n29335), .I0(n2997), .I1(n3017), .CO(n29336));
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n29334), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_14 (.CI(n29334), .I0(n2998), .I1(n3017), .CO(n29335));
    SB_CARRY mod_5_add_1473_3 (.CI(n29134), .I0(n2109), .I1(n43638), .CO(n29135));
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n29333), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_13 (.CI(n29333), .I0(n2999), .I1(n3017), .CO(n29334));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n29332), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_2_lut (.I0(bit_ctr[14]), .I1(bit_ctr[14]), .I2(n43638), 
            .I3(VCC_net), .O(n2209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_12 (.CI(n29332), .I0(n3000), .I1(n3017), .CO(n29333));
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n29331), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_24 (.CI(n27862), .I0(bit_ctr[22]), .I1(GND_net), .CO(n27863));
    SB_CARRY mod_5_add_2076_11 (.CI(n29331), .I0(n3001), .I1(n3017), .CO(n29332));
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(n43638), 
            .CO(n29134));
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n29330), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n1994), .I1(n1994), .I2(n2027), 
            .I3(n29133), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_17_lut (.I0(n1995), .I1(n1995), .I2(n2027), 
            .I3(n29132), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_23_lut (.I0(n25779), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(n27861), .O(n40716)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_2076_10 (.CI(n29330), .I0(n3002), .I1(n3017), .CO(n29331));
    SB_CARRY mod_5_add_1406_17 (.CI(n29132), .I0(n1995), .I1(n2027), .CO(n29133));
    SB_CARRY add_21_23 (.CI(n27861), .I0(bit_ctr[21]), .I1(GND_net), .CO(n27862));
    SB_LUT4 add_21_22_lut (.I0(n25779), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(n27860), .O(n40715)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n29329), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_9 (.CI(n29329), .I0(n3003), .I1(n3017), .CO(n29330));
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n29328), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_8 (.CI(n29328), .I0(n3004), .I1(n3017), .CO(n29329));
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n29327), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_16_lut (.I0(n1996), .I1(n1996), .I2(n2027), 
            .I3(n29131), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_16 (.CI(n29131), .I0(n1996), .I1(n2027), .CO(n29132));
    SB_CARRY mod_5_add_2076_7 (.CI(n29327), .I0(n3005), .I1(n3017), .CO(n29328));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n29326), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_6 (.CI(n29326), .I0(n3006), .I1(n3017), .CO(n29327));
    SB_DFF timer_1223__i0 (.Q(timer[0]), .C(clk32MHz), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY add_21_22 (.CI(n27860), .I0(bit_ctr[20]), .I1(GND_net), .CO(n27861));
    SB_LUT4 add_21_21_lut (.I0(n25779), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(n27859), .O(n40714)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n29325), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_15_lut (.I0(n1997), .I1(n1997), .I2(n2027), 
            .I3(n29130), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_5 (.CI(n29325), .I0(n3007), .I1(n3017), .CO(n29326));
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n29324), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_15 (.CI(n29130), .I0(n1997), .I1(n2027), .CO(n29131));
    SB_CARRY mod_5_add_2076_4 (.CI(n29324), .I0(n3008), .I1(n3017), .CO(n29325));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n3009), .I1(n3009), .I2(n43639), 
            .I3(n29323), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_3 (.CI(n29323), .I0(n3009), .I1(n43639), .CO(n29324));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n43639), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n43639), 
            .CO(n29323));
    SB_LUT4 mod_5_add_1406_14_lut (.I0(n1998), .I1(n1998), .I2(n2027), 
            .I3(n29129), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_14 (.CI(n29129), .I0(n1998), .I1(n2027), .CO(n29130));
    SB_CARRY add_21_21 (.CI(n27859), .I0(bit_ctr[19]), .I1(GND_net), .CO(n27860));
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2885), .I1(n2885), .I2(n2918), 
            .I3(n29322), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_13_lut (.I0(n1999), .I1(n1999), .I2(n2027), 
            .I3(n29128), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(n2886), .I1(n2886), .I2(n2918), 
            .I3(n29321), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_13 (.CI(n29128), .I0(n1999), .I1(n2027), .CO(n29129));
    SB_LUT4 add_21_20_lut (.I0(n25779), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(n27858), .O(n40713)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_2009_26 (.CI(n29321), .I0(n2886), .I1(n2918), .CO(n29322));
    SB_LUT4 mod_5_add_1406_12_lut (.I0(n2000), .I1(n2000), .I2(n2027), 
            .I3(n29127), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hCA3A;
    SB_DFF bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(clk32MHz), .D(n33619));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFE bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(clk32MHz), .E(VCC_net), 
            .D(n33617));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(clk32MHz), .D(n33629));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(clk32MHz), .D(n17687));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(clk32MHz), .D(n17686));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(clk32MHz), .D(n17685));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(clk32MHz), .D(n17684));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(clk32MHz), .D(n17683));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(clk32MHz), .D(n17682));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(clk32MHz), .D(n17681));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(clk32MHz), .D(n17680));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(clk32MHz), .D(n17679));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(clk32MHz), .D(n17678));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(clk32MHz), .D(n17677));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(clk32MHz), .D(n17676));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(clk32MHz), .D(n17675));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(clk32MHz), .D(n17674));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(clk32MHz), .D(n17673));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(clk32MHz), .D(n17672));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(clk32MHz), .D(n17671));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(clk32MHz), .D(n17670));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(clk32MHz), .D(n17669));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(clk32MHz), .D(n17668));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(clk32MHz), .D(n17667));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(clk32MHz), .D(n17666));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(clk32MHz), .D(n17665));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(clk32MHz), .D(n17664));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(clk32MHz), .D(n17663));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(clk32MHz), .D(n17662));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(clk32MHz), .D(n17661));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(clk32MHz), .D(n17660));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(clk32MHz), .D(n17659));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(clk32MHz), .D(n17658));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(clk32MHz), .D(n17657));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i6_4_lut (.I0(bit_ctr[12]), .I1(bit_ctr[23]), .I2(bit_ctr[21]), 
            .I3(bit_ctr[20]), .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut (.I0(bit_ctr[17]), .I1(bit_ctr[31]), .I2(bit_ctr[28]), 
            .I3(bit_ctr[29]), .O(n13));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_4_lut_adj_1610 (.I0(bit_ctr[16]), .I1(bit_ctr[22]), .I2(n13), 
            .I3(n14), .O(n14_adj_4532));
    defparam i5_4_lut_adj_1610.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1611 (.I0(bit_ctr[5]), .I1(bit_ctr[7]), .I2(bit_ctr[14]), 
            .I3(bit_ctr[25]), .O(n15));
    defparam i6_4_lut_adj_1611.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_2_lut_adj_1612 (.I0(bit_ctr[19]), .I1(bit_ctr[27]), .I2(GND_net), 
            .I3(GND_net), .O(n16));
    defparam i3_2_lut_adj_1612.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1613 (.I0(bit_ctr[6]), .I1(bit_ctr[10]), .I2(bit_ctr[15]), 
            .I3(bit_ctr[9]), .O(n22_adj_4533));
    defparam i9_4_lut_adj_1613.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n15), .I1(bit_ctr[30]), .I2(n14_adj_4532), .I3(bit_ctr[24]), 
            .O(n37594));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(bit_ctr[26]), .I1(bit_ctr[3]), .I2(bit_ctr[13]), 
            .I3(bit_ctr[4]), .O(n20));
    defparam i7_4_lut.LUT_INIT = 16'hfefa;
    SB_LUT4 i11_4_lut_adj_1614 (.I0(n37594), .I1(n22_adj_4533), .I2(n16), 
            .I3(bit_ctr[11]), .O(n24));
    defparam i11_4_lut_adj_1614.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1615 (.I0(bit_ctr[18]), .I1(n24), .I2(n20), 
            .I3(bit_ctr[8]), .O(\state_3__N_362[1] ));
    defparam i12_4_lut_adj_1615.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), .I2(GND_net), 
            .I3(GND_net), .O(n15841));   // verilog/neopixel.v(79[18] 99[12])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_3_lut (.I0(one_wire_N_513[3]), .I1(one_wire_N_513[4]), .I2(one_wire_N_513[2]), 
            .I3(GND_net), .O(n30047));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_1616 (.I0(n24922), .I1(one_wire_N_513[4]), .I2(GND_net), 
            .I3(GND_net), .O(n4));
    defparam i1_2_lut_adj_1616.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut_adj_1617 (.I0(\one_wire_N_513[9] ), .I1(\one_wire_N_513[10] ), 
            .I2(\one_wire_N_513[6] ), .I3(\one_wire_N_513[8] ), .O(n13_adj_4534));   // verilog/neopixel.v(104[14:39])
    defparam i5_4_lut_adj_1617.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1618 (.I0(n13_adj_4534), .I1(n11), .I2(\one_wire_N_513[11] ), 
            .I3(n15961), .O(n15776));   // verilog/neopixel.v(104[14:39])
    defparam i7_4_lut_adj_1618.LUT_INIT = 16'hfffe;
    SB_LUT4 i2103_4_lut (.I0(n24962), .I1(\state_3__N_362[1] ), .I2(\state[1] ), 
            .I3(n15841), .O(n4451));
    defparam i2103_4_lut.LUT_INIT = 16'h3f35;
    SB_LUT4 i2_4_lut (.I0(\state[1] ), .I1(n1164), .I2(\state[0] ), .I3(n4451), 
            .O(n4483));
    defparam i2_4_lut.LUT_INIT = 16'hfe0e;
    SB_CARRY add_21_20 (.CI(n27858), .I0(bit_ctr[18]), .I1(GND_net), .CO(n27859));
    SB_LUT4 i3_2_lut_adj_1619 (.I0(n2491), .I1(n2504), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_4535));
    defparam i3_2_lut_adj_1619.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut_adj_1620 (.I0(n2496), .I1(n2505), .I2(n2500), .I3(n2499), 
            .O(n34_adj_4536));
    defparam i13_4_lut_adj_1620.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut (.I0(bit_ctr[10]), .I1(n2497), .I2(n2509), .I3(GND_net), 
            .O(n22_adj_4537));
    defparam i1_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i17_4_lut_adj_1621 (.I0(n2490), .I1(n34_adj_4536), .I2(n24_adj_4535), 
            .I3(n2494), .O(n38_adj_4538));
    defparam i17_4_lut_adj_1621.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1622 (.I0(n2501), .I1(n2502), .I2(n2506), .I3(n2492), 
            .O(n36));
    defparam i15_4_lut_adj_1622.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1623 (.I0(n2495), .I1(n2498), .I2(n2493), .I3(n22_adj_4537), 
            .O(n37_adj_4539));
    defparam i16_4_lut_adj_1623.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1624 (.I0(n2507), .I1(n2508), .I2(n2503), .I3(n2489), 
            .O(n35_adj_4540));
    defparam i14_4_lut_adj_1624.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut (.I0(n35_adj_4540), .I1(n37_adj_4539), .I2(n36), 
            .I3(n38_adj_4538), .O(n2522));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36785_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43630));
    defparam i36785_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i7_4_lut_adj_1625 (.I0(n1505), .I1(n1508), .I2(n1503), .I3(n1499), 
            .O(n18_adj_4541));
    defparam i7_4_lut_adj_1625.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1626 (.I0(bit_ctr[20]), .I1(n1504), .I2(n1509), 
            .I3(n1507), .O(n17));
    defparam i6_4_lut_adj_1626.LUT_INIT = 16'hffec;
    SB_LUT4 i8_4_lut_adj_1627 (.I0(n1502), .I1(n1506), .I2(n1501), .I3(n1500), 
            .O(n19));
    defparam i8_4_lut_adj_1627.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_3_lut (.I0(n19), .I1(n17), .I2(n18_adj_4541), .I3(GND_net), 
            .O(n1532));
    defparam i10_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i36793_1_lut (.I0(n2126), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43638));
    defparam i36793_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_21_19_lut (.I0(n25779), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(n27857), .O(n40712)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_19 (.CI(n27857), .I0(bit_ctr[17]), .I1(GND_net), .CO(n27858));
    SB_LUT4 i16_4_lut_adj_1628 (.I0(n21), .I1(n23), .I2(n22_adj_4542), 
            .I3(n24_adj_4543), .O(n36_adj_4544));   // verilog/neopixel.v(104[14:39])
    defparam i16_4_lut_adj_1628.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1629 (.I0(n25_adj_4545), .I1(n27_adj_4546), .I2(n26_adj_4547), 
            .I3(n28_adj_4548), .O(n37_adj_4549));   // verilog/neopixel.v(104[14:39])
    defparam i17_4_lut_adj_1629.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1630 (.I0(n37_adj_4549), .I1(n29), .I2(n36_adj_4544), 
            .I3(n30_adj_4550), .O(n15961));   // verilog/neopixel.v(104[14:39])
    defparam i19_4_lut_adj_1630.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1631 (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n34976));
    defparam i1_2_lut_adj_1631.LUT_INIT = 16'h2222;
    SB_LUT4 i28984_2_lut (.I0(one_wire_N_513[3]), .I1(one_wire_N_513[2]), 
            .I2(GND_net), .I3(GND_net), .O(n35738));
    defparam i28984_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20201_2_lut (.I0(n30206), .I1(one_wire_N_513[3]), .I2(GND_net), 
            .I3(GND_net), .O(n24922));
    defparam i20201_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19977_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(GND_net), .I3(GND_net), .O(n24698));
    defparam i19977_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(one_wire_N_513[4]), .I1(n35021), .I2(n24922), 
            .I3(n35738), .O(n116));
    defparam i1_4_lut.LUT_INIT = 16'h45cd;
    SB_LUT4 i36757_3_lut (.I0(n35873), .I1(n116), .I2(n15961), .I3(GND_net), 
            .O(n37672));
    defparam i36757_3_lut.LUT_INIT = 16'hfbfb;
    SB_CARRY mod_5_add_1406_12 (.CI(n29127), .I0(n2000), .I1(n2027), .CO(n29128));
    SB_LUT4 mod_5_add_2009_25_lut (.I0(n2887), .I1(n2887), .I2(n2918), 
            .I3(n29320), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_11_lut (.I0(n2001), .I1(n2001), .I2(n2027), 
            .I3(n29126), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_18_lut (.I0(n25779), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(n27856), .O(n40709)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_2009_25 (.CI(n29320), .I0(n2887), .I1(n2918), .CO(n29321));
    SB_CARRY mod_5_add_1406_11 (.CI(n29126), .I0(n2001), .I1(n2027), .CO(n29127));
    SB_LUT4 mod_5_add_2009_24_lut (.I0(n2888), .I1(n2888), .I2(n2918), 
            .I3(n29319), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_10_lut (.I0(n2002), .I1(n2002), .I2(n2027), 
            .I3(n29125), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_24 (.CI(n29319), .I0(n2888), .I1(n2918), .CO(n29320));
    SB_CARRY mod_5_add_1406_10 (.CI(n29125), .I0(n2002), .I1(n2027), .CO(n29126));
    SB_LUT4 mod_5_add_2009_23_lut (.I0(n2889), .I1(n2889), .I2(n2918), 
            .I3(n29318), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_9_lut (.I0(n2003), .I1(n2003), .I2(n2027), 
            .I3(n29124), .O(n2102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_18 (.CI(n27856), .I0(bit_ctr[16]), .I1(GND_net), .CO(n27857));
    SB_CARRY mod_5_add_2009_23 (.CI(n29318), .I0(n2889), .I1(n2918), .CO(n29319));
    SB_CARRY mod_5_add_1406_9 (.CI(n29124), .I0(n2003), .I1(n2027), .CO(n29125));
    SB_LUT4 mod_5_add_2009_22_lut (.I0(n2890), .I1(n2890), .I2(n2918), 
            .I3(n29317), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1406_8_lut (.I0(n2004), .I1(n2004), .I2(n2027), 
            .I3(n29123), .O(n2103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_22 (.CI(n29317), .I0(n2890), .I1(n2918), .CO(n29318));
    SB_CARRY mod_5_add_1406_8 (.CI(n29123), .I0(n2004), .I1(n2027), .CO(n29124));
    SB_LUT4 mod_5_add_1406_7_lut (.I0(n2005), .I1(n2005), .I2(n2027), 
            .I3(n29122), .O(n2104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_21_lut (.I0(n2891), .I1(n2891), .I2(n2918), 
            .I3(n29316), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_7 (.CI(n29122), .I0(n2005), .I1(n2027), .CO(n29123));
    SB_CARRY mod_5_add_2009_21 (.CI(n29316), .I0(n2891), .I1(n2918), .CO(n29317));
    SB_LUT4 mod_5_add_1406_6_lut (.I0(n2006), .I1(n2006), .I2(n2027), 
            .I3(n29121), .O(n2105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_20_lut (.I0(n2892), .I1(n2892), .I2(n2918), 
            .I3(n29315), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_6 (.CI(n29121), .I0(n2006), .I1(n2027), .CO(n29122));
    SB_CARRY mod_5_add_2009_20 (.CI(n29315), .I0(n2892), .I1(n2918), .CO(n29316));
    SB_LUT4 mod_5_add_1406_5_lut (.I0(n2007), .I1(n2007), .I2(n2027), 
            .I3(n29120), .O(n2106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_19_lut (.I0(n2893), .I1(n2893), .I2(n2918), 
            .I3(n29314), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_5 (.CI(n29120), .I0(n2007), .I1(n2027), .CO(n29121));
    SB_CARRY mod_5_add_2009_19 (.CI(n29314), .I0(n2893), .I1(n2918), .CO(n29315));
    SB_LUT4 mod_5_add_1406_4_lut (.I0(n2008), .I1(n2008), .I2(n2027), 
            .I3(n29119), .O(n2107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_18_lut (.I0(n2894), .I1(n2894), .I2(n2918), 
            .I3(n29313), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_4 (.CI(n29119), .I0(n2008), .I1(n2027), .CO(n29120));
    SB_CARRY mod_5_add_2009_18 (.CI(n29313), .I0(n2894), .I1(n2918), .CO(n29314));
    SB_LUT4 mod_5_add_1406_3_lut (.I0(n2009), .I1(n2009), .I2(n43640), 
            .I3(n29118), .O(n2108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2009_17_lut (.I0(n2895), .I1(n2895), .I2(n2918), 
            .I3(n29312), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_3 (.CI(n29118), .I0(n2009), .I1(n43640), .CO(n29119));
    SB_CARRY mod_5_add_2009_17 (.CI(n29312), .I0(n2895), .I1(n2918), .CO(n29313));
    SB_LUT4 mod_5_add_1406_2_lut (.I0(bit_ctr[15]), .I1(bit_ctr[15]), .I2(n43640), 
            .I3(VCC_net), .O(n2109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_2009_16_lut (.I0(n2896), .I1(n2896), .I2(n2918), 
            .I3(n29311), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(n43640), 
            .CO(n29118));
    SB_CARRY mod_5_add_2009_16 (.CI(n29311), .I0(n2896), .I1(n2918), .CO(n29312));
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1895), .I1(n1895), .I2(n1928), 
            .I3(n29117), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_15_lut (.I0(n2897), .I1(n2897), .I2(n2918), 
            .I3(n29310), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_16_lut (.I0(n1896), .I1(n1896), .I2(n1928), 
            .I3(n29116), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_15 (.CI(n29310), .I0(n2897), .I1(n2918), .CO(n29311));
    SB_CARRY mod_5_add_1339_16 (.CI(n29116), .I0(n1896), .I1(n1928), .CO(n29117));
    SB_LUT4 mod_5_add_2009_14_lut (.I0(n2898), .I1(n2898), .I2(n2918), 
            .I3(n29309), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_15_lut (.I0(n1897), .I1(n1897), .I2(n1928), 
            .I3(n29115), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_14 (.CI(n29309), .I0(n2898), .I1(n2918), .CO(n29310));
    SB_CARRY mod_5_add_1339_15 (.CI(n29115), .I0(n1897), .I1(n1928), .CO(n29116));
    SB_LUT4 mod_5_add_2009_13_lut (.I0(n2899), .I1(n2899), .I2(n2918), 
            .I3(n29308), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_14_lut (.I0(n1898), .I1(n1898), .I2(n1928), 
            .I3(n29114), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_13 (.CI(n29308), .I0(n2899), .I1(n2918), .CO(n29309));
    SB_CARRY mod_5_add_1339_14 (.CI(n29114), .I0(n1898), .I1(n1928), .CO(n29115));
    SB_LUT4 mod_5_add_1339_13_lut (.I0(n1899), .I1(n1899), .I2(n1928), 
            .I3(n29113), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_17_lut (.I0(n25779), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(n27855), .O(n40708)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2009_12_lut (.I0(n2900), .I1(n2900), .I2(n2918), 
            .I3(n29307), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_12 (.CI(n29307), .I0(n2900), .I1(n2918), .CO(n29308));
    SB_CARRY mod_5_add_1339_13 (.CI(n29113), .I0(n1899), .I1(n1928), .CO(n29114));
    SB_DFFE state_i1 (.Q(\state[1] ), .C(clk32MHz), .E(VCC_net), .D(n17625));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2009_11_lut (.I0(n2901), .I1(n2901), .I2(n2918), 
            .I3(n29306), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_12_lut (.I0(n1900), .I1(n1900), .I2(n1928), 
            .I3(n29112), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_11 (.CI(n29306), .I0(n2901), .I1(n2918), .CO(n29307));
    SB_LUT4 mod_5_add_2009_10_lut (.I0(n2902), .I1(n2902), .I2(n2918), 
            .I3(n29305), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_10 (.CI(n29305), .I0(n2902), .I1(n2918), .CO(n29306));
    SB_LUT4 mod_5_add_2009_9_lut (.I0(n2903), .I1(n2903), .I2(n2918), 
            .I3(n29304), .O(n3002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i14_4_lut_adj_1632 (.I0(n2591), .I1(n2608), .I2(n2601), .I3(n2605), 
            .O(n36_adj_4551));
    defparam i14_4_lut_adj_1632.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1339_12 (.CI(n29112), .I0(n1900), .I1(n1928), .CO(n29113));
    SB_CARRY mod_5_add_2009_9 (.CI(n29304), .I0(n2903), .I1(n2918), .CO(n29305));
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(clk32MHz), .E(n17203), .D(\state_3__N_362[0] ), 
            .S(n35833));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1339_11_lut (.I0(n1901), .I1(n1901), .I2(n1928), 
            .I3(n29111), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2009_8_lut (.I0(n2904), .I1(n2904), .I2(n2918), 
            .I3(n29303), .O(n3003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_8 (.CI(n29303), .I0(n2904), .I1(n2918), .CO(n29304));
    SB_CARRY mod_5_add_1339_11 (.CI(n29111), .I0(n1901), .I1(n1928), .CO(n29112));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(n2905), .I1(n2905), .I2(n2918), 
            .I3(n29302), .O(n3004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_10_lut (.I0(n1902), .I1(n1902), .I2(n1928), 
            .I3(n29110), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_7 (.CI(n29302), .I0(n2905), .I1(n2918), .CO(n29303));
    SB_CARRY mod_5_add_1339_10 (.CI(n29110), .I0(n1902), .I1(n1928), .CO(n29111));
    SB_LUT4 i3_3_lut (.I0(n2606), .I1(bit_ctr[9]), .I2(n2609), .I3(GND_net), 
            .O(n25_adj_4552));
    defparam i3_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 mod_5_add_1339_9_lut (.I0(n1903), .I1(n1903), .I2(n1928), 
            .I3(n29109), .O(n2002)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_9 (.CI(n29109), .I0(n1903), .I1(n1928), .CO(n29110));
    SB_LUT4 mod_5_add_2009_6_lut (.I0(n2906), .I1(n2906), .I2(n2918), 
            .I3(n29301), .O(n3005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_8_lut (.I0(n1904), .I1(n1904), .I2(n1928), 
            .I3(n29108), .O(n2003)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2009_6 (.CI(n29301), .I0(n2906), .I1(n2918), .CO(n29302));
    SB_CARRY mod_5_add_1339_8 (.CI(n29108), .I0(n1904), .I1(n1928), .CO(n29109));
    SB_CARRY add_21_17 (.CI(n27855), .I0(bit_ctr[15]), .I1(GND_net), .CO(n27856));
    SB_LUT4 mod_5_add_2009_5_lut (.I0(n2907), .I1(n2907), .I2(n2918), 
            .I3(n29300), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_7_lut (.I0(n1905), .I1(n1905), .I2(n1928), 
            .I3(n29107), .O(n2004)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_16_lut (.I0(n25779), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(n27854), .O(n40704)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_16 (.CI(n27854), .I0(bit_ctr[14]), .I1(GND_net), .CO(n27855));
    SB_LUT4 i12_4_lut_adj_1633 (.I0(n2593), .I1(n2596), .I2(n2600), .I3(n2590), 
            .O(n34_adj_4553));
    defparam i12_4_lut_adj_1633.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1634 (.I0(n25_adj_4552), .I1(n36_adj_4551), .I2(n2594), 
            .I3(n2589), .O(n40_adj_4554));
    defparam i18_4_lut_adj_1634.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2009_5 (.CI(n29300), .I0(n2907), .I1(n2918), .CO(n29301));
    SB_CARRY mod_5_add_1339_7 (.CI(n29107), .I0(n1905), .I1(n1928), .CO(n29108));
    SB_LUT4 mod_5_add_2009_4_lut (.I0(n2908), .I1(n2908), .I2(n2918), 
            .I3(n29299), .O(n3007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_6_lut (.I0(n1906), .I1(n1906), .I2(n1928), 
            .I3(n29106), .O(n2005)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_15_lut (.I0(n25779), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(n27853), .O(n40703)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_4_lut (.I0(n35682), .I1(n14452), .I2(n807), .I3(bit_ctr[27]), 
            .O(n838));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0405;
    SB_LUT4 mod_5_i606_3_lut_4_lut (.I0(n14452), .I1(bit_ctr[27]), .I2(n838), 
            .I3(n35682), .O(n35829));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i606_3_lut_4_lut.LUT_INIT = 16'hf40b;
    SB_CARRY mod_5_add_2009_4 (.CI(n29299), .I0(n2908), .I1(n2918), .CO(n29300));
    SB_CARRY mod_5_add_1339_6 (.CI(n29106), .I0(n1906), .I1(n1928), .CO(n29107));
    SB_LUT4 mod_5_add_1339_5_lut (.I0(n1907), .I1(n1907), .I2(n1928), 
            .I3(n29105), .O(n2006)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i34513_3_lut_4_lut (.I0(bit_ctr[29]), .I1(n24982), .I2(n35706), 
            .I3(bit_ctr[28]), .O(n35682));
    defparam i34513_3_lut_4_lut.LUT_INIT = 16'h9666;
    SB_DFF bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(clk32MHz), .D(n17458));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i19769_2_lut_3_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(bit_ctr[29]), 
            .I3(GND_net), .O(n24488));   // verilog/neopixel.v(22[26:36])
    defparam i19769_2_lut_3_lut.LUT_INIT = 16'h2020;
    SB_LUT4 mod_5_add_2009_3_lut (.I0(n2909), .I1(n2909), .I2(n43641), 
            .I3(n29298), .O(n3008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2009_3 (.CI(n29298), .I0(n2909), .I1(n43641), .CO(n29299));
    SB_CARRY mod_5_add_1339_5 (.CI(n29105), .I0(n1907), .I1(n1928), .CO(n29106));
    SB_LUT4 mod_5_add_2009_2_lut (.I0(bit_ctr[6]), .I1(bit_ctr[6]), .I2(n43641), 
            .I3(VCC_net), .O(n3009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hA3AC;
    SB_DFFESR one_wire_108 (.Q(PIN_8_c), .C(clk32MHz), .E(n17155), .D(\neo_pixel_transmitter.done_N_576 ), 
            .R(n37483));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1339_4_lut (.I0(n1908), .I1(n1908), .I2(n1928), 
            .I3(n29104), .O(n2007)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_4 (.CI(n29104), .I0(n1908), .I1(n1928), .CO(n29105));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(n1909), .I1(n1909), .I2(n43642), 
            .I3(n29103), .O(n2008)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY add_21_15 (.CI(n27853), .I0(bit_ctr[13]), .I1(GND_net), .CO(n27854));
    SB_LUT4 add_21_14_lut (.I0(n25779), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(n27852), .O(n40702)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1339_3 (.CI(n29103), .I0(n1909), .I1(n43642), .CO(n29104));
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(n43641), 
            .CO(n29298));
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2786), .I1(n2786), .I2(n2819), 
            .I3(n29297), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1339_2_lut (.I0(bit_ctr[16]), .I1(bit_ctr[16]), .I2(n43642), 
            .I3(VCC_net), .O(n2009)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(n2787), .I1(n2787), .I2(n2819), 
            .I3(n29296), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(n43642), 
            .CO(n29103));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1796), .I1(n1796), .I2(n1829), 
            .I3(n29102), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(n1797), .I1(n1797), .I2(n1829), 
            .I3(n29101), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_25 (.CI(n29296), .I0(n2787), .I1(n2819), .CO(n29297));
    SB_CARRY mod_5_add_1272_15 (.CI(n29101), .I0(n1797), .I1(n1829), .CO(n29102));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(n2788), .I1(n2788), .I2(n2819), 
            .I3(n29295), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_14_lut (.I0(n1798), .I1(n1798), .I2(n1829), 
            .I3(n29100), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_24 (.CI(n29295), .I0(n2788), .I1(n2819), .CO(n29296));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(n2789), .I1(n2789), .I2(n2819), 
            .I3(n29294), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_14 (.CI(n29100), .I0(n1798), .I1(n1829), .CO(n29101));
    SB_CARRY mod_5_add_1942_23 (.CI(n29294), .I0(n2789), .I1(n2819), .CO(n29295));
    SB_LUT4 mod_5_add_1272_13_lut (.I0(n1799), .I1(n1799), .I2(n1829), 
            .I3(n29099), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_22_lut (.I0(n2790), .I1(n2790), .I2(n2819), 
            .I3(n29293), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_13 (.CI(n29099), .I0(n1799), .I1(n1829), .CO(n29100));
    SB_CARRY mod_5_add_1942_22 (.CI(n29293), .I0(n2790), .I1(n2819), .CO(n29294));
    SB_LUT4 mod_5_add_1272_12_lut (.I0(n1800), .I1(n1800), .I2(n1829), 
            .I3(n29098), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_21_lut (.I0(n2791), .I1(n2791), .I2(n2819), 
            .I3(n29292), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_12 (.CI(n29098), .I0(n1800), .I1(n1829), .CO(n29099));
    SB_LUT4 i14_4_lut_adj_1635 (.I0(n3004), .I1(n2989), .I2(n2990), .I3(n3007), 
            .O(n40_adj_4555));
    defparam i14_4_lut_adj_1635.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1636 (.I0(n3006), .I1(n2984), .I2(n2988), .I3(n2986), 
            .O(n44));
    defparam i18_4_lut_adj_1636.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1637 (.I0(n3008), .I1(n3003), .I2(n2994), .I3(n3002), 
            .O(n42));
    defparam i16_4_lut_adj_1637.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1272_11_lut (.I0(n1801), .I1(n1801), .I2(n1829), 
            .I3(n29097), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i17_4_lut_adj_1638 (.I0(n2999), .I1(n3000), .I2(n2992), .I3(n2997), 
            .O(n43_adj_4556));
    defparam i17_4_lut_adj_1638.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1639 (.I0(n2996), .I1(n2985), .I2(n2995), .I3(n2987), 
            .O(n41_adj_4557));
    defparam i15_4_lut_adj_1639.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_2_lut (.I0(n3001), .I1(n2993), .I2(GND_net), .I3(GND_net), 
            .O(n38_adj_4558));
    defparam i12_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20_3_lut (.I0(n2998), .I1(n40_adj_4555), .I2(n2991), .I3(GND_net), 
            .O(n46_adj_4559));
    defparam i20_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i24_4_lut_adj_1640 (.I0(n41_adj_4557), .I1(n43_adj_4556), .I2(n42), 
            .I3(n44), .O(n50));
    defparam i24_4_lut_adj_1640.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_3_lut (.I0(n3005), .I1(bit_ctr[5]), .I2(n3009), .I3(GND_net), 
            .O(n37_adj_4560));
    defparam i11_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i25_4_lut (.I0(n37_adj_4560), .I1(n50), .I2(n46_adj_4559), 
            .I3(n38_adj_4558), .O(n3017));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36791_1_lut (.I0(n3116), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43636));
    defparam i36791_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1942_21 (.CI(n29292), .I0(n2791), .I1(n2819), .CO(n29293));
    SB_LUT4 i16_4_lut_adj_1641 (.I0(n2602), .I1(n2588), .I2(n2604), .I3(n2607), 
            .O(n38_adj_4561));
    defparam i16_4_lut_adj_1641.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1272_11 (.CI(n29097), .I0(n1801), .I1(n1829), .CO(n29098));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(n1802), .I1(n1802), .I2(n1829), 
            .I3(n29096), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i17_3_lut (.I0(n2598), .I1(n34_adj_4553), .I2(n2603), .I3(GND_net), 
            .O(n39_adj_4562));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i15_4_lut_adj_1642 (.I0(n2592), .I1(n2597), .I2(n2595), .I3(n2599), 
            .O(n37_adj_4563));
    defparam i15_4_lut_adj_1642.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1643 (.I0(n37_adj_4563), .I1(n39_adj_4562), .I2(n38_adj_4561), 
            .I3(n40_adj_4554), .O(n2621));
    defparam i21_4_lut_adj_1643.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1272_10 (.CI(n29096), .I0(n1802), .I1(n1829), .CO(n29097));
    SB_LUT4 mod_5_add_1272_9_lut (.I0(n1803), .I1(n1803), .I2(n1829), 
            .I3(n29095), .O(n1902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_20_lut (.I0(n2792), .I1(n2792), .I2(n2819), 
            .I3(n29291), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_20 (.CI(n29291), .I0(n2792), .I1(n2819), .CO(n29292));
    SB_CARRY mod_5_add_1272_9 (.CI(n29095), .I0(n1803), .I1(n1829), .CO(n29096));
    SB_LUT4 mod_5_add_1942_19_lut (.I0(n2793), .I1(n2793), .I2(n2819), 
            .I3(n29290), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_8_lut (.I0(n1804), .I1(n1804), .I2(n1829), 
            .I3(n29094), .O(n1903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(n905), .I2(VCC_net), 
            .I3(n28245), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(n906), .I2(VCC_net), 
            .I3(n28244), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_6 (.CI(n28244), .I0(n906), .I1(VCC_net), .CO(n28245));
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n35829), .I2(VCC_net), 
            .I3(n28243), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_5 (.CI(n28243), .I0(n35829), .I1(VCC_net), 
            .CO(n28244));
    SB_CARRY mod_5_add_1942_19 (.CI(n29290), .I0(n2793), .I1(n2819), .CO(n29291));
    SB_CARRY mod_5_add_1272_8 (.CI(n29094), .I0(n1804), .I1(n1829), .CO(n29095));
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n17296), .I2(VCC_net), 
            .I3(n28242), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_4 (.CI(n28242), .I0(n17296), .I1(VCC_net), 
            .CO(n28243));
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n14450), .I2(GND_net), 
            .I3(n28241), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_3 (.CI(n28241), .I0(n14450), .I1(GND_net), 
            .CO(n28242));
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n28241));
    SB_LUT4 mod_5_add_736_8_lut (.I0(n4_adj_4564), .I1(n4_adj_4564), .I2(n1037), 
            .I3(n28240), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_7_lut (.I0(n1005), .I1(n1005), .I2(n1037), .I3(n28239), 
            .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_14 (.CI(n27852), .I0(bit_ctr[12]), .I1(GND_net), .CO(n27853));
    SB_CARRY mod_5_add_736_7 (.CI(n28239), .I0(n1005), .I1(n1037), .CO(n28240));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(n2794), .I1(n2794), .I2(n2819), 
            .I3(n29289), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_7_lut (.I0(n1805), .I1(n1805), .I2(n1829), 
            .I3(n29093), .O(n1904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_18 (.CI(n29289), .I0(n2794), .I1(n2819), .CO(n29290));
    SB_CARRY mod_5_add_1272_7 (.CI(n29093), .I0(n1805), .I1(n1829), .CO(n29094));
    SB_LUT4 mod_5_add_736_6_lut (.I0(n1006), .I1(n1006), .I2(n1037), .I3(n28238), 
            .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_6 (.CI(n28238), .I0(n1006), .I1(n1037), .CO(n28239));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(n2795), .I1(n2795), .I2(n2819), 
            .I3(n29288), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_6_lut (.I0(n1806), .I1(n1806), .I2(n1829), 
            .I3(n29092), .O(n1905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_6 (.CI(n29092), .I0(n1806), .I1(n1829), .CO(n29093));
    SB_LUT4 mod_5_add_736_5_lut (.I0(n1007), .I1(n1007), .I2(n1037), .I3(n28237), 
            .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_5 (.CI(n28237), .I0(n1007), .I1(n1037), .CO(n28238));
    SB_CARRY mod_5_add_1942_17 (.CI(n29288), .I0(n2795), .I1(n2819), .CO(n29289));
    SB_LUT4 mod_5_add_1272_5_lut (.I0(n1807), .I1(n1807), .I2(n1829), 
            .I3(n29091), .O(n1906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n28236), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1272_5 (.CI(n29091), .I0(n1807), .I1(n1829), .CO(n29092));
    SB_CARRY mod_5_add_736_4 (.CI(n28236), .I0(n1008), .I1(n1037), .CO(n28237));
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n43645), 
            .I3(n28235), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_3 (.CI(n28235), .I0(n1009), .I1(n43645), .CO(n28236));
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n43645), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1942_16_lut (.I0(n2796), .I1(n2796), .I2(n2819), 
            .I3(n29287), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_4_lut (.I0(n1808), .I1(n1808), .I2(n1829), 
            .I3(n29090), .O(n1907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_16 (.CI(n29287), .I0(n2796), .I1(n2819), .CO(n29288));
    SB_CARRY mod_5_add_1272_4 (.CI(n29090), .I0(n1808), .I1(n1829), .CO(n29091));
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n43645), 
            .CO(n28235));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(n2797), .I1(n2797), .I2(n2819), 
            .I3(n29286), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1272_3_lut (.I0(n1809), .I1(n1809), .I2(n43644), 
            .I3(n29089), .O(n1908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_3 (.CI(n29089), .I0(n1809), .I1(n43644), .CO(n29090));
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n28234), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n28233), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_8 (.CI(n28233), .I0(n1104), .I1(n1136), .CO(n28234));
    SB_CARRY mod_5_add_1942_15 (.CI(n29286), .I0(n2797), .I1(n2819), .CO(n29287));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(bit_ctr[17]), .I1(bit_ctr[17]), .I2(n43644), 
            .I3(VCC_net), .O(n1909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(n43644), 
            .CO(n29089));
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n28232), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_7 (.CI(n28232), .I0(n1105), .I1(n1136), .CO(n28233));
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n28231), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_6 (.CI(n28231), .I0(n1106), .I1(n1136), .CO(n28232));
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n28230), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_5 (.CI(n28230), .I0(n1107), .I1(n1136), .CO(n28231));
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n28229), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_14_lut (.I0(n2798), .I1(n2798), .I2(n2819), 
            .I3(n29285), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n29088), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_4 (.CI(n28229), .I0(n1108), .I1(n1136), .CO(n28230));
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n43646), 
            .I3(n28228), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1942_14 (.CI(n29285), .I0(n2798), .I1(n2819), .CO(n29286));
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n29087), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_3 (.CI(n28228), .I0(n1109), .I1(n43646), .CO(n28229));
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n43646), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n43646), 
            .CO(n28228));
    SB_LUT4 mod_5_add_1942_13_lut (.I0(n2799), .I1(n2799), .I2(n2819), 
            .I3(n29284), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_14 (.CI(n29087), .I0(n1698), .I1(n1730), .CO(n29088));
    SB_DFF timer_1223__i1 (.Q(timer[1]), .C(clk32MHz), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY mod_5_add_1942_13 (.CI(n29284), .I0(n2799), .I1(n2819), .CO(n29285));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n29086), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_13_lut (.I0(n25779), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(n27851), .O(n40700)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_13 (.CI(n27851), .I0(bit_ctr[11]), .I1(GND_net), .CO(n27852));
    SB_DFF timer_1223__i2 (.Q(timer[2]), .C(clk32MHz), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i3 (.Q(timer[3]), .C(clk32MHz), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i4 (.Q(timer[4]), .C(clk32MHz), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i5 (.Q(timer[5]), .C(clk32MHz), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i6 (.Q(timer[6]), .C(clk32MHz), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i7 (.Q(timer[7]), .C(clk32MHz), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i8 (.Q(timer[8]), .C(clk32MHz), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i9 (.Q(timer[9]), .C(clk32MHz), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i10 (.Q(timer[10]), .C(clk32MHz), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i11 (.Q(timer[11]), .C(clk32MHz), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i12 (.Q(timer[12]), .C(clk32MHz), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i13 (.Q(timer[13]), .C(clk32MHz), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i14 (.Q(timer[14]), .C(clk32MHz), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i15 (.Q(timer[15]), .C(clk32MHz), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i16 (.Q(timer[16]), .C(clk32MHz), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i17 (.Q(timer[17]), .C(clk32MHz), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i18 (.Q(timer[18]), .C(clk32MHz), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i19 (.Q(timer[19]), .C(clk32MHz), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i20 (.Q(timer[20]), .C(clk32MHz), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i21 (.Q(timer[21]), .C(clk32MHz), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i22 (.Q(timer[22]), .C(clk32MHz), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i23 (.Q(timer[23]), .C(clk32MHz), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i24 (.Q(timer[24]), .C(clk32MHz), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i25 (.Q(timer[25]), .C(clk32MHz), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i26 (.Q(timer[26]), .C(clk32MHz), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i27 (.Q(timer[27]), .C(clk32MHz), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i28 (.Q(timer[28]), .C(clk32MHz), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i29 (.Q(timer[29]), .C(clk32MHz), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i30 (.Q(timer[30]), .C(clk32MHz), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1223__i31 (.Q(timer[31]), .C(clk32MHz), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_DFF start_103 (.Q(start), .C(clk32MHz), .D(n33675));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(clk32MHz), .D(n17444));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n28221), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n28220), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n28220), .I0(n1203), .I1(n1235), .CO(n28221));
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n28219), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_8 (.CI(n28219), .I0(n1204), .I1(n1235), .CO(n28220));
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n28218), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_7 (.CI(n28218), .I0(n1205), .I1(n1235), .CO(n28219));
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n28217), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_6 (.CI(n28217), .I0(n1206), .I1(n1235), .CO(n28218));
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n28216), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_5 (.CI(n28216), .I0(n1207), .I1(n1235), .CO(n28217));
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n28215), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_4 (.CI(n28215), .I0(n1208), .I1(n1235), .CO(n28216));
    SB_LUT4 mod_5_add_1942_12_lut (.I0(n2800), .I1(n2800), .I2(n2819), 
            .I3(n29283), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n43648), 
            .I3(n28214), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_12_lut (.I0(n25779), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(n27850), .O(n40699)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_870_3 (.CI(n28214), .I0(n1209), .I1(n43648), .CO(n28215));
    SB_CARRY mod_5_add_1205_13 (.CI(n29086), .I0(n1699), .I1(n1730), .CO(n29087));
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n43648), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n43648), 
            .CO(n28214));
    SB_CARRY mod_5_add_1942_12 (.CI(n29283), .I0(n2800), .I1(n2819), .CO(n29284));
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n29085), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_12 (.CI(n29085), .I0(n1700), .I1(n1730), .CO(n29086));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(n2801), .I1(n2801), .I2(n2819), 
            .I3(n29282), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n29084), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_11 (.CI(n29084), .I0(n1701), .I1(n1730), .CO(n29085));
    SB_CARRY mod_5_add_1942_11 (.CI(n29282), .I0(n2801), .I1(n2819), .CO(n29283));
    SB_LUT4 mod_5_add_1942_10_lut (.I0(n2802), .I1(n2802), .I2(n2819), 
            .I3(n29281), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n29083), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_10 (.CI(n29083), .I0(n1702), .I1(n1730), .CO(n29084));
    SB_CARRY add_21_12 (.CI(n27850), .I0(bit_ctr[10]), .I1(GND_net), .CO(n27851));
    SB_CARRY mod_5_add_1942_10 (.CI(n29281), .I0(n2802), .I1(n2819), .CO(n29282));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n29082), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_9_lut (.I0(n2803), .I1(n2803), .I2(n2819), 
            .I3(n29280), .O(n2902)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_9 (.CI(n29082), .I0(n1703), .I1(n1730), .CO(n29083));
    SB_CARRY mod_5_add_1942_9 (.CI(n29280), .I0(n2803), .I1(n2819), .CO(n29281));
    SB_LUT4 mod_5_add_1942_8_lut (.I0(n2804), .I1(n2804), .I2(n2819), 
            .I3(n29279), .O(n2903)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_8 (.CI(n29279), .I0(n2804), .I1(n2819), .CO(n29280));
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n29081), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_8 (.CI(n29081), .I0(n1704), .I1(n1730), .CO(n29082));
    SB_LUT4 mod_5_add_1942_7_lut (.I0(n2805), .I1(n2805), .I2(n2819), 
            .I3(n29278), .O(n2904)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n29080), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_11_lut (.I0(n25779), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(n27849), .O(n40698)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1942_7 (.CI(n29278), .I0(n2805), .I1(n2819), .CO(n29279));
    SB_CARRY mod_5_add_1205_7 (.CI(n29080), .I0(n1705), .I1(n1730), .CO(n29081));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(n2806), .I1(n2806), .I2(n2819), 
            .I3(n29277), .O(n2905)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_11 (.CI(n27849), .I0(bit_ctr[9]), .I1(GND_net), .CO(n27850));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n29079), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1942_6 (.CI(n29277), .I0(n2806), .I1(n2819), .CO(n29278));
    SB_CARRY mod_5_add_1205_6 (.CI(n29079), .I0(n1706), .I1(n1730), .CO(n29080));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n29078), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1942_5_lut (.I0(n2807), .I1(n2807), .I2(n2819), 
            .I3(n29276), .O(n2906)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_10_lut (.I0(n25779), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(n27848), .O(n40707)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1205_5 (.CI(n29078), .I0(n1707), .I1(n1730), .CO(n29079));
    SB_CARRY mod_5_add_1942_5 (.CI(n29276), .I0(n2807), .I1(n2819), .CO(n29277));
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n29077), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_4 (.CI(n29077), .I0(n1708), .I1(n1730), .CO(n29078));
    SB_CARRY add_21_10 (.CI(n27848), .I0(bit_ctr[8]), .I1(GND_net), .CO(n27849));
    SB_LUT4 add_21_9_lut (.I0(n25779), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(n27847), .O(n40706)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1942_4_lut (.I0(n2808), .I1(n2808), .I2(n2819), 
            .I3(n29275), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n43647), 
            .I3(n29076), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 i1_2_lut_adj_1644 (.I0(n2103), .I1(n2097), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4565));
    defparam i1_2_lut_adj_1644.LUT_INIT = 16'heeee;
    SB_CARRY add_21_9 (.CI(n27847), .I0(bit_ctr[7]), .I1(GND_net), .CO(n27848));
    SB_CARRY mod_5_add_1942_4 (.CI(n29275), .I0(n2808), .I1(n2819), .CO(n29276));
    SB_LUT4 i20155_2_lut (.I0(bit_ctr[14]), .I1(n2109), .I2(GND_net), 
            .I3(GND_net), .O(n24876));
    defparam i20155_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mod_5_add_1205_3 (.CI(n29076), .I0(n1709), .I1(n43647), .CO(n29077));
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1301), .I1(n1301), .I2(n1334), 
            .I3(n28204), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n43647), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1942_3_lut (.I0(n2809), .I1(n2809), .I2(n43643), 
            .I3(n29274), .O(n2908)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n43647), 
            .CO(n29076));
    SB_LUT4 add_21_8_lut (.I0(n25779), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(n27846), .O(n40701)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1942_3 (.CI(n29274), .I0(n2809), .I1(n43643), .CO(n29275));
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1598), .I1(n1598), .I2(n1631), 
            .I3(n29075), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_937_10_lut (.I0(n1302), .I1(n1302), .I2(n1334), 
            .I3(n28203), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_10 (.CI(n28203), .I0(n1302), .I1(n1334), .CO(n28204));
    SB_LUT4 mod_5_add_937_9_lut (.I0(n1303), .I1(n1303), .I2(n1334), .I3(n28202), 
            .O(n1402)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_8 (.CI(n27846), .I0(bit_ctr[6]), .I1(GND_net), .CO(n27847));
    SB_LUT4 mod_5_add_1942_2_lut (.I0(bit_ctr[7]), .I1(bit_ctr[7]), .I2(n43643), 
            .I3(VCC_net), .O(n2909)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(n1599), .I1(n1599), .I2(n1631), 
            .I3(n29074), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i13_4_lut_adj_1645 (.I0(n2102), .I1(n2099), .I2(n2100), .I3(n18_adj_4565), 
            .O(n30_adj_4566));
    defparam i13_4_lut_adj_1645.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_7_lut (.I0(n25779), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(n27845), .O(n40711)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_21_7 (.CI(n27845), .I0(bit_ctr[5]), .I1(GND_net), .CO(n27846));
    SB_CARRY mod_5_add_1138_13 (.CI(n29074), .I0(n1599), .I1(n1631), .CO(n29075));
    SB_LUT4 add_21_6_lut (.I0(n25779), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(n27844), .O(n40710)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_937_9 (.CI(n28202), .I0(n1303), .I1(n1334), .CO(n28203));
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(n43643), 
            .CO(n29274));
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2687), .I1(n2687), .I2(n2720), 
            .I3(n29273), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_12_lut (.I0(n1600), .I1(n1600), .I2(n1631), 
            .I3(n29073), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_12 (.CI(n29073), .I0(n1600), .I1(n1631), .CO(n29074));
    SB_LUT4 mod_5_add_937_8_lut (.I0(n1304), .I1(n1304), .I2(n1334), .I3(n28201), 
            .O(n1403)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i11_4_lut_adj_1646 (.I0(n2098), .I1(n2106), .I2(n2093), .I3(n24876), 
            .O(n28_adj_4567));
    defparam i11_4_lut_adj_1646.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1875_24_lut (.I0(n2688), .I1(n2688), .I2(n2720), 
            .I3(n29272), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_8 (.CI(n28201), .I0(n1304), .I1(n1334), .CO(n28202));
    SB_LUT4 mod_5_add_1138_11_lut (.I0(n1601), .I1(n1601), .I2(n1631), 
            .I3(n29072), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_6 (.CI(n27844), .I0(bit_ctr[4]), .I1(GND_net), .CO(n27845));
    SB_CARRY mod_5_add_1875_24 (.CI(n29272), .I0(n2688), .I1(n2720), .CO(n29273));
    SB_LUT4 add_21_5_lut (.I0(n25779), .I1(bit_ctr[3]), .I2(GND_net), 
            .I3(n27843), .O(n40705)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_937_7_lut (.I0(n1305), .I1(n1305), .I2(n1334), .I3(n28200), 
            .O(n1404)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_23_lut (.I0(n2689), .I1(n2689), .I2(n2720), 
            .I3(n29271), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_11 (.CI(n29072), .I0(n1601), .I1(n1631), .CO(n29073));
    SB_CARRY mod_5_add_937_7 (.CI(n28200), .I0(n1305), .I1(n1334), .CO(n28201));
    SB_CARRY add_21_5 (.CI(n27843), .I0(bit_ctr[3]), .I1(GND_net), .CO(n27844));
    SB_LUT4 mod_5_add_937_6_lut (.I0(n1306), .I1(n1306), .I2(n1334), .I3(n28199), 
            .O(n1405)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_10_lut (.I0(n1602), .I1(n1602), .I2(n1631), 
            .I3(n29071), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_23 (.CI(n29271), .I0(n2689), .I1(n2720), .CO(n29272));
    SB_CARRY mod_5_add_1138_10 (.CI(n29071), .I0(n1602), .I1(n1631), .CO(n29072));
    SB_LUT4 mod_5_add_1875_22_lut (.I0(n2690), .I1(n2690), .I2(n2720), 
            .I3(n29270), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_937_6 (.CI(n28199), .I0(n1306), .I1(n1334), .CO(n28200));
    SB_LUT4 mod_5_add_937_5_lut (.I0(n1307), .I1(n1307), .I2(n1334), .I3(n28198), 
            .O(n1406)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_9_lut (.I0(n1603), .I1(n1603), .I2(n1631), 
            .I3(n29070), .O(n1702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_9 (.CI(n29070), .I0(n1603), .I1(n1631), .CO(n29071));
    SB_CARRY mod_5_add_937_5 (.CI(n28198), .I0(n1307), .I1(n1334), .CO(n28199));
    SB_CARRY mod_5_add_1875_22 (.CI(n29270), .I0(n2690), .I1(n2720), .CO(n29271));
    SB_LUT4 mod_5_add_1138_8_lut (.I0(n1604), .I1(n1604), .I2(n1631), 
            .I3(n29069), .O(n1703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_4_lut (.I0(n25779), .I1(bit_ctr[2]), .I2(GND_net), 
            .I3(n27842), .O(n40619)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1875_21_lut (.I0(n2691), .I1(n2691), .I2(n2720), 
            .I3(n29269), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_21 (.CI(n29269), .I0(n2691), .I1(n2720), .CO(n29270));
    SB_CARRY mod_5_add_1138_8 (.CI(n29069), .I0(n1604), .I1(n1631), .CO(n29070));
    SB_LUT4 mod_5_add_1875_20_lut (.I0(n2692), .I1(n2692), .I2(n2720), 
            .I3(n29268), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_7_lut (.I0(n1605), .I1(n1605), .I2(n1631), 
            .I3(n29068), .O(n1704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_4 (.CI(n27842), .I0(bit_ctr[2]), .I1(GND_net), .CO(n27843));
    SB_LUT4 mod_5_add_937_4_lut (.I0(n1308), .I1(n1308), .I2(n1334), .I3(n28197), 
            .O(n1407)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_3_lut (.I0(n25779), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(n27841), .O(n40620)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_937_4 (.CI(n28197), .I0(n1308), .I1(n1334), .CO(n28198));
    SB_CARRY mod_5_add_1875_20 (.CI(n29268), .I0(n2692), .I1(n2720), .CO(n29269));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(n2693), .I1(n2693), .I2(n2720), 
            .I3(n29267), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_7 (.CI(n29068), .I0(n1605), .I1(n1631), .CO(n29069));
    SB_LUT4 i12_4_lut_adj_1647 (.I0(n2108), .I1(n2095), .I2(n2096), .I3(n2105), 
            .O(n29_adj_4568));
    defparam i12_4_lut_adj_1647.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_937_3_lut (.I0(n1309), .I1(n1309), .I2(n43649), 
            .I3(n28196), .O(n1408)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_3 (.CI(n28196), .I0(n1309), .I1(n43649), .CO(n28197));
    SB_LUT4 mod_5_add_937_2_lut (.I0(bit_ctr[22]), .I1(bit_ctr[22]), .I2(n43649), 
            .I3(VCC_net), .O(n1409)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(n43649), 
            .CO(n28196));
    SB_CARRY add_21_3 (.CI(n27841), .I0(bit_ctr[1]), .I1(GND_net), .CO(n27842));
    SB_LUT4 mod_5_add_1138_6_lut (.I0(n1606), .I1(n1606), .I2(n1631), 
            .I3(n29067), .O(n1705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_19 (.CI(n29267), .I0(n2693), .I1(n2720), .CO(n29268));
    SB_CARRY mod_5_add_1138_6 (.CI(n29067), .I0(n1606), .I1(n1631), .CO(n29068));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(n1607), .I1(n1607), .I2(n1631), 
            .I3(n29066), .O(n1706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_18_lut (.I0(n2694), .I1(n2694), .I2(n2720), 
            .I3(n29266), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_5 (.CI(n29066), .I0(n1607), .I1(n1631), .CO(n29067));
    SB_CARRY mod_5_add_1875_18 (.CI(n29266), .I0(n2694), .I1(n2720), .CO(n29267));
    SB_LUT4 mod_5_add_1138_4_lut (.I0(n1608), .I1(n1608), .I2(n1631), 
            .I3(n29065), .O(n1707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_17_lut (.I0(n2695), .I1(n2695), .I2(n2720), 
            .I3(n29265), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1138_4 (.CI(n29065), .I0(n1608), .I1(n1631), .CO(n29066));
    SB_CARRY mod_5_add_1875_17 (.CI(n29265), .I0(n2695), .I1(n2720), .CO(n29266));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(n1609), .I1(n1609), .I2(n43650), 
            .I3(n29064), .O(n1708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1138_3 (.CI(n29064), .I0(n1609), .I1(n43650), .CO(n29065));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(n2696), .I1(n2696), .I2(n2720), 
            .I3(n29264), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1138_2_lut (.I0(bit_ctr[19]), .I1(bit_ctr[19]), .I2(n43650), 
            .I3(VCC_net), .O(n1709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 add_21_2_lut (.I0(n25779), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n40616)) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(n43650), 
            .CO(n29064));
    SB_LUT4 i10_4_lut_adj_1648 (.I0(n2101), .I1(n2104), .I2(n2107), .I3(n2094), 
            .O(n27_adj_4569));
    defparam i10_4_lut_adj_1648.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1875_16 (.CI(n29264), .I0(n2696), .I1(n2720), .CO(n29265));
    SB_LUT4 mod_5_add_1875_15_lut (.I0(n2697), .I1(n2697), .I2(n2720), 
            .I3(n29263), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_15 (.CI(n29263), .I0(n2697), .I1(n2720), .CO(n29264));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(n2698), .I1(n2698), .I2(n2720), 
            .I3(n29262), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_14 (.CI(n29262), .I0(n2698), .I1(n2720), .CO(n29263));
    SB_LUT4 mod_5_add_1875_13_lut (.I0(n2699), .I1(n2699), .I2(n2720), 
            .I3(n29261), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_13 (.CI(n29261), .I0(n2699), .I1(n2720), .CO(n29262));
    SB_LUT4 mod_5_add_1875_12_lut (.I0(n2700), .I1(n2700), .I2(n2720), 
            .I3(n29260), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_12 (.CI(n29260), .I0(n2700), .I1(n2720), .CO(n29261));
    SB_LUT4 mod_5_add_1875_11_lut (.I0(n2701), .I1(n2701), .I2(n2720), 
            .I3(n29259), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_11 (.CI(n29259), .I0(n2701), .I1(n2720), .CO(n29260));
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n27841));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(n2702), .I1(n2702), .I2(n2720), 
            .I3(n29258), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_10 (.CI(n29258), .I0(n2702), .I1(n2720), .CO(n29259));
    SB_LUT4 mod_5_add_1875_9_lut (.I0(n2703), .I1(n2703), .I2(n2720), 
            .I3(n29257), .O(n2802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_9 (.CI(n29257), .I0(n2703), .I1(n2720), .CO(n29258));
    SB_LUT4 i16_4_lut_adj_1649 (.I0(n27_adj_4569), .I1(n29_adj_4568), .I2(n28_adj_4567), 
            .I3(n30_adj_4566), .O(n2126));
    defparam i16_4_lut_adj_1649.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1875_8_lut (.I0(n2704), .I1(n2704), .I2(n2720), 
            .I3(n29256), .O(n2803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_8 (.CI(n29256), .I0(n2704), .I1(n2720), .CO(n29257));
    SB_LUT4 mod_5_add_1875_7_lut (.I0(n2705), .I1(n2705), .I2(n2720), 
            .I3(n29255), .O(n2804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_7 (.CI(n29255), .I0(n2705), .I1(n2720), .CO(n29256));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(n2706), .I1(n2706), .I2(n2720), 
            .I3(n29254), .O(n2805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1400), .I1(n1400), .I2(n1433), 
            .I3(n28132), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1875_6 (.CI(n29254), .I0(n2706), .I1(n2720), .CO(n29255));
    SB_LUT4 mod_5_add_1004_11_lut (.I0(n1401), .I1(n1401), .I2(n1433), 
            .I3(n28131), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_11 (.CI(n28131), .I0(n1401), .I1(n1433), .CO(n28132));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(n1402), .I1(n1402), .I2(n1433), 
            .I3(n28130), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_10 (.CI(n28130), .I0(n1402), .I1(n1433), .CO(n28131));
    SB_LUT4 mod_5_add_1004_9_lut (.I0(n1403), .I1(n1403), .I2(n1433), 
            .I3(n28129), .O(n1502)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_5_lut (.I0(n2707), .I1(n2707), .I2(n2720), 
            .I3(n29253), .O(n2806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_9 (.CI(n28129), .I0(n1403), .I1(n1433), .CO(n28130));
    SB_CARRY mod_5_add_1875_5 (.CI(n29253), .I0(n2707), .I1(n2720), .CO(n29254));
    SB_LUT4 mod_5_add_1004_8_lut (.I0(n1404), .I1(n1404), .I2(n1433), 
            .I3(n28128), .O(n1503)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_8 (.CI(n28128), .I0(n1404), .I1(n1433), .CO(n28129));
    SB_LUT4 mod_5_add_1004_7_lut (.I0(n1405), .I1(n1405), .I2(n1433), 
            .I3(n28127), .O(n1504)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_7 (.CI(n28127), .I0(n1405), .I1(n1433), .CO(n28128));
    SB_LUT4 mod_5_add_1004_6_lut (.I0(n1406), .I1(n1406), .I2(n1433), 
            .I3(n28126), .O(n1505)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_6 (.CI(n28126), .I0(n1406), .I1(n1433), .CO(n28127));
    SB_LUT4 mod_5_add_1004_5_lut (.I0(n1407), .I1(n1407), .I2(n1433), 
            .I3(n28125), .O(n1506)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1875_4_lut (.I0(n2708), .I1(n2708), .I2(n2720), 
            .I3(n29252), .O(n2807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_5 (.CI(n28125), .I0(n1407), .I1(n1433), .CO(n28126));
    SB_CARRY mod_5_add_1875_4 (.CI(n29252), .I0(n2708), .I1(n2720), .CO(n29253));
    SB_LUT4 mod_5_add_1004_4_lut (.I0(n1408), .I1(n1408), .I2(n1433), 
            .I3(n28124), .O(n1507)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1004_4 (.CI(n28124), .I0(n1408), .I1(n1433), .CO(n28125));
    SB_LUT4 mod_5_add_1004_3_lut (.I0(n1409), .I1(n1409), .I2(n43652), 
            .I3(n28123), .O(n1508)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1004_3 (.CI(n28123), .I0(n1409), .I1(n43652), .CO(n28124));
    SB_LUT4 mod_5_add_1004_2_lut (.I0(bit_ctr[21]), .I1(bit_ctr[21]), .I2(n43652), 
            .I3(VCC_net), .O(n1509)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(n43652), 
            .CO(n28123));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(n2709), .I1(n2709), .I2(n43651), 
            .I3(n29251), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_3 (.CI(n29251), .I0(n2709), .I1(n43651), .CO(n29252));
    SB_LUT4 mod_5_add_1875_2_lut (.I0(bit_ctr[8]), .I1(bit_ctr[8]), .I2(n43651), 
            .I3(VCC_net), .O(n2809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(n43651), 
            .CO(n29251));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n29250), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n29249), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_23 (.CI(n29249), .I0(n2589), .I1(n2621), .CO(n29250));
    SB_LUT4 sub_14_add_2_33_lut (.I0(one_wire_N_513[25]), .I1(timer[31]), 
            .I2(n1[31]), .I3(n28100), .O(n22_adj_4542)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 sub_14_add_2_32_lut (.I0(one_wire_N_513[24]), .I1(timer[30]), 
            .I2(n1[30]), .I3(n28099), .O(n23)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_32 (.CI(n28099), .I0(timer[30]), .I1(n1[30]), 
            .CO(n28100));
    SB_LUT4 sub_14_add_2_31_lut (.I0(one_wire_N_513[19]), .I1(timer[29]), 
            .I2(n1[29]), .I3(n28098), .O(n28_adj_4548)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_31 (.CI(n28098), .I0(timer[29]), .I1(n1[29]), 
            .CO(n28099));
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n29248), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_30_lut (.I0(one_wire_N_513[26]), .I1(timer[28]), 
            .I2(n1[28]), .I3(n28097), .O(n26_adj_4547)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1808_22 (.CI(n29248), .I0(n2590), .I1(n2621), .CO(n29249));
    SB_CARRY sub_14_add_2_30 (.CI(n28097), .I0(timer[28]), .I1(n1[28]), 
            .CO(n28098));
    SB_LUT4 sub_14_add_2_29_lut (.I0(one_wire_N_513[18]), .I1(timer[27]), 
            .I2(n1[27]), .I3(n28096), .O(n21)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_29 (.CI(n28096), .I0(timer[27]), .I1(n1[27]), 
            .CO(n28097));
    SB_LUT4 sub_14_add_2_28_lut (.I0(GND_net), .I1(timer[26]), .I2(n1[26]), 
            .I3(n28095), .O(one_wire_N_513[26])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_28 (.CI(n28095), .I0(timer[26]), .I1(n1[26]), 
            .CO(n28096));
    SB_LUT4 sub_14_add_2_27_lut (.I0(GND_net), .I1(timer[25]), .I2(n1[25]), 
            .I3(n28094), .O(one_wire_N_513[25])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n29247), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_21 (.CI(n29247), .I0(n2591), .I1(n2621), .CO(n29248));
    SB_CARRY sub_14_add_2_27 (.CI(n28094), .I0(timer[25]), .I1(n1[25]), 
            .CO(n28095));
    SB_LUT4 sub_14_add_2_26_lut (.I0(GND_net), .I1(timer[24]), .I2(n1[24]), 
            .I3(n28093), .O(one_wire_N_513[24])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_26 (.CI(n28093), .I0(timer[24]), .I1(n1[24]), 
            .CO(n28094));
    SB_LUT4 sub_14_add_2_25_lut (.I0(one_wire_N_513[16]), .I1(timer[23]), 
            .I2(n1[23]), .I3(n28092), .O(n30_adj_4550)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_25 (.CI(n28092), .I0(timer[23]), .I1(n1[23]), 
            .CO(n28093));
    SB_LUT4 sub_14_add_2_24_lut (.I0(one_wire_N_513[13]), .I1(timer[22]), 
            .I2(n1[22]), .I3(n28091), .O(n24_adj_4543)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_24 (.CI(n28091), .I0(timer[22]), .I1(n1[22]), 
            .CO(n28092));
    SB_LUT4 sub_14_add_2_23_lut (.I0(one_wire_N_513[14]), .I1(timer[21]), 
            .I2(n1[21]), .I3(n28090), .O(n25_adj_4545)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_23 (.CI(n28090), .I0(timer[21]), .I1(n1[21]), 
            .CO(n28091));
    SB_LUT4 sub_14_add_2_22_lut (.I0(one_wire_N_513[15]), .I1(timer[20]), 
            .I2(n1[20]), .I3(n28089), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_22 (.CI(n28089), .I0(timer[20]), .I1(n1[20]), 
            .CO(n28090));
    SB_LUT4 sub_14_add_2_21_lut (.I0(GND_net), .I1(timer[19]), .I2(n1[19]), 
            .I3(n28088), .O(one_wire_N_513[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_21 (.CI(n28088), .I0(timer[19]), .I1(n1[19]), 
            .CO(n28089));
    SB_LUT4 sub_14_add_2_20_lut (.I0(GND_net), .I1(timer[18]), .I2(n1[18]), 
            .I3(n28087), .O(one_wire_N_513[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_20 (.CI(n28087), .I0(timer[18]), .I1(n1[18]), 
            .CO(n28088));
    SB_LUT4 sub_14_add_2_19_lut (.I0(one_wire_N_513[12]), .I1(timer[17]), 
            .I2(n1[17]), .I3(n28086), .O(n27_adj_4546)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_19 (.CI(n28086), .I0(timer[17]), .I1(n1[17]), 
            .CO(n28087));
    SB_LUT4 sub_14_add_2_18_lut (.I0(GND_net), .I1(timer[16]), .I2(n1[16]), 
            .I3(n28085), .O(one_wire_N_513[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_18 (.CI(n28085), .I0(timer[16]), .I1(n1[16]), 
            .CO(n28086));
    SB_LUT4 sub_14_add_2_17_lut (.I0(GND_net), .I1(timer[15]), .I2(n1[15]), 
            .I3(n28084), .O(one_wire_N_513[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n29246), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_17 (.CI(n28084), .I0(timer[15]), .I1(n1[15]), 
            .CO(n28085));
    SB_LUT4 sub_14_add_2_16_lut (.I0(GND_net), .I1(timer[14]), .I2(n1[14]), 
            .I3(n28083), .O(one_wire_N_513[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_16 (.CI(n28083), .I0(timer[14]), .I1(n1[14]), 
            .CO(n28084));
    SB_LUT4 sub_14_add_2_15_lut (.I0(GND_net), .I1(timer[13]), .I2(n1[13]), 
            .I3(n28082), .O(one_wire_N_513[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_20 (.CI(n29246), .I0(n2592), .I1(n2621), .CO(n29247));
    SB_CARRY sub_14_add_2_15 (.CI(n28082), .I0(timer[13]), .I1(n1[13]), 
            .CO(n28083));
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n29245), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_14_lut (.I0(GND_net), .I1(timer[12]), .I2(n1[12]), 
            .I3(n28081), .O(one_wire_N_513[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_14 (.CI(n28081), .I0(timer[12]), .I1(n1[12]), 
            .CO(n28082));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n28080), .O(\one_wire_N_513[11] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_13 (.CI(n28080), .I0(timer[11]), .I1(n1[11]), 
            .CO(n28081));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n28079), .O(\one_wire_N_513[10] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_12 (.CI(n28079), .I0(timer[10]), .I1(n1[10]), 
            .CO(n28080));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n28078), .O(\one_wire_N_513[9] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_11 (.CI(n28078), .I0(timer[9]), .I1(n1[9]), 
            .CO(n28079));
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n28077), .O(\one_wire_N_513[8] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_10 (.CI(n28077), .I0(timer[8]), .I1(n1[8]), 
            .CO(n28078));
    SB_CARRY mod_5_add_1808_19 (.CI(n29245), .I0(n2593), .I1(n2621), .CO(n29246));
    SB_LUT4 sub_14_add_2_9_lut (.I0(one_wire_N_513[5]), .I1(timer[7]), .I2(n1[7]), 
            .I3(n28076), .O(n11)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_9 (.CI(n28076), .I0(timer[7]), .I1(n1[7]), .CO(n28077));
    SB_LUT4 sub_14_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n28075), .O(\one_wire_N_513[6] )) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_8 (.CI(n28075), .I0(timer[6]), .I1(n1[6]), .CO(n28076));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n29244), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_18 (.CI(n29244), .I0(n2594), .I1(n2621), .CO(n29245));
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n28074), .O(one_wire_N_513[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_7 (.CI(n28074), .I0(timer[5]), .I1(n1[5]), .CO(n28075));
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n28073), .O(one_wire_N_513[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_6 (.CI(n28073), .I0(timer[4]), .I1(n1[4]), .CO(n28074));
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n29243), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n28072), .O(one_wire_N_513[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_5 (.CI(n28072), .I0(timer[3]), .I1(n1[3]), .CO(n28073));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n28071), .O(one_wire_N_513[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_4 (.CI(n28071), .I0(timer[2]), .I1(n1[2]), .CO(n28072));
    SB_CARRY mod_5_add_1808_17 (.CI(n29243), .I0(n2595), .I1(n2621), .CO(n29244));
    SB_LUT4 sub_14_add_2_3_lut (.I0(n4_adj_4592), .I1(timer[1]), .I2(n1[1]), 
            .I3(n28070), .O(n30206)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_3 (.CI(n28070), .I0(timer[1]), .I1(n1[1]), .CO(n28071));
    SB_LUT4 sub_14_add_2_2_lut (.I0(one_wire_N_513[2]), .I1(timer[0]), .I2(n1[0]), 
            .I3(VCC_net), .O(n4_adj_4592)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_2_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n29242), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n28070));
    SB_CARRY mod_5_add_1808_16 (.CI(n29242), .I0(n2596), .I1(n2621), .CO(n29243));
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n29241), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_15 (.CI(n29241), .I0(n2597), .I1(n2621), .CO(n29242));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n29240), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_14 (.CI(n29240), .I0(n2598), .I1(n2621), .CO(n29241));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n29239), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_13 (.CI(n29239), .I0(n2599), .I1(n2621), .CO(n29240));
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n29238), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_12 (.CI(n29238), .I0(n2600), .I1(n2621), .CO(n29239));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n29237), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_11 (.CI(n29237), .I0(n2601), .I1(n2621), .CO(n29238));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n29236), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_10 (.CI(n29236), .I0(n2602), .I1(n2621), .CO(n29237));
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n29235), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i36792_1_lut (.I0(n2225), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43637));
    defparam i36792_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i10_4_lut_adj_1650 (.I0(n2193), .I1(n2194), .I2(n2206), .I3(n2204), 
            .O(n28_adj_4594));
    defparam i10_4_lut_adj_1650.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1651 (.I0(n2203), .I1(n28_adj_4594), .I2(bit_ctr[13]), 
            .I3(n2209), .O(n32_adj_4595));
    defparam i14_4_lut_adj_1651.LUT_INIT = 16'hfeee;
    SB_LUT4 i12_4_lut_adj_1652 (.I0(n2208), .I1(n2201), .I2(n2192), .I3(n2196), 
            .O(n30_adj_4596));
    defparam i12_4_lut_adj_1652.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1653 (.I0(n2195), .I1(n2207), .I2(n2205), .I3(n2199), 
            .O(n31_adj_4597));
    defparam i13_4_lut_adj_1653.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i11_4_lut_adj_1654 (.I0(n2202), .I1(n2197), .I2(n2198), .I3(n2200), 
            .O(n29_adj_4598));
    defparam i11_4_lut_adj_1654.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1655 (.I0(n29_adj_4598), .I1(n31_adj_4597), .I2(n30_adj_4596), 
            .I3(n32_adj_4595), .O(n2225));
    defparam i17_4_lut_adj_1655.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36789_1_lut (.I0(n2324), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43634));
    defparam i36789_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut (.I0(n24984), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[1] ), .O(n36198));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 i23_3_lut_4_lut (.I0(n24922), .I1(one_wire_N_513[4]), .I2(n30047), 
            .I3(\state[0] ), .O(n35720));
    defparam i23_3_lut_4_lut.LUT_INIT = 16'hf0ee;
    SB_LUT4 i9_2_lut (.I0(n3084), .I1(n3092), .I2(GND_net), .I3(GND_net), 
            .O(n36_adj_4599));
    defparam i9_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i19_4_lut_adj_1656 (.I0(n3085), .I1(n3094), .I2(n3093), .I3(n3108), 
            .O(n46_adj_4600));
    defparam i19_4_lut_adj_1656.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1657 (.I0(n3087), .I1(n3107), .I2(n3088), .I3(n3086), 
            .O(n42_adj_4601));
    defparam i15_4_lut_adj_1657.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1658 (.I0(bit_ctr[4]), .I1(n3103), .I2(n3109), 
            .I3(GND_net), .O(n34_adj_4602));
    defparam i7_3_lut_adj_1658.LUT_INIT = 16'hecec;
    SB_LUT4 i16_4_lut_adj_1659 (.I0(n3100), .I1(n3083), .I2(n3089), .I3(n3101), 
            .O(n43_adj_4603));
    defparam i16_4_lut_adj_1659.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(n3104), .I1(n46_adj_4600), .I2(n36_adj_4599), 
            .I3(n3091), .O(n50_adj_4604));
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1660 (.I0(n3105), .I1(n42_adj_4601), .I2(n3098), 
            .I3(n3096), .O(n48));
    defparam i21_4_lut_adj_1660.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1661 (.I0(n43_adj_4603), .I1(n3099), .I2(n34_adj_4602), 
            .I3(n3090), .O(n49));
    defparam i22_4_lut_adj_1661.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1662 (.I0(n3102), .I1(n3095), .I2(n3106), .I3(n3097), 
            .O(n47_adj_4605));
    defparam i20_4_lut_adj_1662.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut (.I0(n47_adj_4605), .I1(n49), .I2(n48), .I3(n50_adj_4604), 
            .O(n3116));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36806_1_lut (.I0(n2720), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43651));
    defparam i36806_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36807_1_lut (.I0(n1433), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43652));
    defparam i36807_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19848_2_lut (.I0(bit_ctr[21]), .I1(n1409), .I2(GND_net), 
            .I3(GND_net), .O(n24567));
    defparam i19848_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i6_4_lut_adj_1663 (.I0(n1405), .I1(n24567), .I2(n1403), .I3(n1406), 
            .O(n16_adj_4606));
    defparam i6_4_lut_adj_1663.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1664 (.I0(n1402), .I1(n1404), .I2(n1400), .I3(n1407), 
            .O(n17_adj_4607));
    defparam i7_4_lut_adj_1664.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1665 (.I0(n17_adj_4607), .I1(n1408), .I2(n16_adj_4606), 
            .I3(n1401), .O(n1433));
    defparam i9_4_lut_adj_1665.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i471_3_lut_3_lut_4_lut_4_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), 
            .I2(n24488), .I3(bit_ctr[29]), .O(n708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i471_3_lut_3_lut_4_lut_4_lut.LUT_INIT = 16'hd622;
    SB_LUT4 i36805_1_lut (.I0(n1631), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43650));
    defparam i36805_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36804_1_lut (.I0(n1334), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43649));
    defparam i36804_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_2_lut (.I0(n2693), .I1(n2704), .I2(GND_net), .I3(GND_net), 
            .O(n28_adj_4608));
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i15_4_lut_adj_1666 (.I0(n2699), .I1(n2706), .I2(n2694), .I3(n2691), 
            .O(n38_adj_4609));
    defparam i15_4_lut_adj_1666.LUT_INIT = 16'hfffe;
    SB_LUT4 i20183_2_lut (.I0(bit_ctr[8]), .I1(n2709), .I2(GND_net), .I3(GND_net), 
            .O(n24904));
    defparam i20183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13_4_lut_adj_1667 (.I0(n2701), .I1(n2696), .I2(n2697), .I3(n24904), 
            .O(n36_adj_4610));
    defparam i13_4_lut_adj_1667.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1668 (.I0(n2700), .I1(n38_adj_4609), .I2(n28_adj_4608), 
            .I3(n2705), .O(n42_adj_4611));
    defparam i19_4_lut_adj_1668.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1669 (.I0(n2702), .I1(n2690), .I2(n2689), .I3(n2708), 
            .O(n40_adj_4612));
    defparam i17_4_lut_adj_1669.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1670 (.I0(n2687), .I1(n36_adj_4610), .I2(n2703), 
            .I3(n2695), .O(n41_adj_4613));
    defparam i18_4_lut_adj_1670.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1671 (.I0(n2688), .I1(n2698), .I2(n2692), .I3(n2707), 
            .O(n39_adj_4614));
    defparam i16_4_lut_adj_1671.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1672 (.I0(n39_adj_4614), .I1(n41_adj_4613), .I2(n40_adj_4612), 
            .I3(n42_adj_4611), .O(n2720));
    defparam i22_4_lut_adj_1672.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1673 (.I0(n1608), .I1(n1606), .I2(n1604), .I3(n1603), 
            .O(n20_adj_4615));
    defparam i8_4_lut_adj_1673.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1674 (.I0(bit_ctr[19]), .I1(n1602), .I2(n1609), 
            .I3(GND_net), .O(n13_adj_4616));
    defparam i1_3_lut_adj_1674.LUT_INIT = 16'hecec;
    SB_LUT4 i6_2_lut (.I0(n1598), .I1(n1600), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4617));
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1675 (.I0(n13_adj_4616), .I1(n20_adj_4615), .I2(n1605), 
            .I3(n1599), .O(n22_adj_4618));
    defparam i10_4_lut_adj_1675.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1676 (.I0(n1601), .I1(n22_adj_4618), .I2(n18_adj_4617), 
            .I3(n1607), .O(n1631));
    defparam i11_4_lut_adj_1676.LUT_INIT = 16'hfffe;
    SB_LUT4 i36798_1_lut (.I0(n2819), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43643));
    defparam i36798_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_2_lut_adj_1677 (.I0(n1304), .I1(n1305), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_4619));
    defparam i1_2_lut_adj_1677.LUT_INIT = 16'heeee;
    SB_LUT4 i3_3_lut_adj_1678 (.I0(bit_ctr[22]), .I1(n1303), .I2(n1309), 
            .I3(GND_net), .O(n12_adj_4620));
    defparam i3_3_lut_adj_1678.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1679 (.I0(n1306), .I1(n1308), .I2(n1302), .I3(n10_adj_4619), 
            .O(n16_adj_4621));
    defparam i7_4_lut_adj_1679.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1680 (.I0(n1307), .I1(n16_adj_4621), .I2(n12_adj_4620), 
            .I3(n1301), .O(n1334));
    defparam i8_4_lut_adj_1680.LUT_INIT = 16'hfffe;
    SB_LUT4 i36802_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43647));
    defparam i36802_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36803_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43648));
    defparam i36803_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6_4_lut_adj_1681 (.I0(n1205), .I1(n1204), .I2(n1203), .I3(n1207), 
            .O(n14_adj_4622));
    defparam i6_4_lut_adj_1681.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1682 (.I0(bit_ctr[23]), .I1(n1206), .I2(n1209), 
            .I3(GND_net), .O(n9_adj_4623));
    defparam i1_3_lut_adj_1682.LUT_INIT = 16'hecec;
    SB_LUT4 i7_4_lut_adj_1683 (.I0(n9_adj_4623), .I1(n14_adj_4622), .I2(n1202), 
            .I3(n1208), .O(n1235));
    defparam i7_4_lut_adj_1683.LUT_INIT = 16'hfffe;
    SB_LUT4 i36801_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43646));
    defparam i36801_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_3_lut (.I0(bit_ctr[18]), .I1(n1699), .I2(n1709), .I3(GND_net), 
            .O(n17_adj_4624));
    defparam i4_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i8_4_lut_adj_1684 (.I0(n1698), .I1(n1707), .I2(n1703), .I3(n1705), 
            .O(n21_adj_4625));
    defparam i8_4_lut_adj_1684.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_3_lut_adj_1685 (.I0(n1704), .I1(n1701), .I2(n1708), .I3(GND_net), 
            .O(n20_adj_4626));
    defparam i7_3_lut_adj_1685.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1686 (.I0(n21_adj_4625), .I1(n17_adj_4624), .I2(n1702), 
            .I3(n1697), .O(n24_adj_4627));
    defparam i11_4_lut_adj_1686.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1687 (.I0(n1700), .I1(n24_adj_4627), .I2(n20_adj_4626), 
            .I3(n1706), .O(n1730));
    defparam i12_4_lut_adj_1687.LUT_INIT = 16'hfffe;
    SB_LUT4 i20079_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n24800));
    defparam i20079_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1688 (.I0(n1105), .I1(n1103), .I2(n24800), .I3(n1108), 
            .O(n12_adj_4628));
    defparam i5_4_lut_adj_1688.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1689 (.I0(n1107), .I1(n12_adj_4628), .I2(n1106), 
            .I3(n1104), .O(n1136));
    defparam i6_4_lut_adj_1689.LUT_INIT = 16'hfffe;
    SB_LUT4 i36799_1_lut (.I0(n1829), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43644));
    defparam i36799_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36800_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43645));
    defparam i36800_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36768_2_lut (.I0(n31409), .I1(n971[28]), .I2(GND_net), .I3(GND_net), 
            .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam i36768_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i36770_2_lut (.I0(n31409), .I1(n971[29]), .I2(GND_net), .I3(GND_net), 
            .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam i36770_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n31409), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i675_3_lut (.I0(n14450), .I1(n971[27]), .I2(n31409), 
            .I3(GND_net), .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i672_3_lut (.I0(n906), .I1(n971[30]), .I2(n31409), .I3(GND_net), 
            .O(n1005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i672_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31760_3_lut (.I0(n905), .I1(n906), .I2(n35829), .I3(GND_net), 
            .O(n38528));
    defparam i31760_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(bit_ctr[26]), .I1(n38528), .I2(n17296), .I3(n14450), 
            .O(n31409));
    defparam i4_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 i31801_3_lut (.I0(n971[28]), .I1(n971[31]), .I2(n971[29]), 
            .I3(GND_net), .O(n38573));
    defparam i31801_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_adj_1690 (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), 
            .I3(GND_net), .O(n6_adj_4629));
    defparam i2_3_lut_adj_1690.LUT_INIT = 16'heaea;
    SB_LUT4 i3_4_lut (.I0(n31409), .I1(n6_adj_4629), .I2(n1005), .I3(n38573), 
            .O(n1037));
    defparam i3_4_lut.LUT_INIT = 16'hfdfc;
    SB_LUT4 i36764_2_lut (.I0(n31409), .I1(n971[31]), .I2(GND_net), .I3(GND_net), 
            .O(n4_adj_4564));   // verilog/neopixel.v(22[26:36])
    defparam i36764_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1691 (.I0(bit_ctr[27]), .I1(n838), .I2(GND_net), 
            .I3(GND_net), .O(n14450));
    defparam i1_2_lut_adj_1691.LUT_INIT = 16'h9999;
    SB_LUT4 mod_5_i605_3_lut (.I0(n807), .I1(n60), .I2(n838), .I3(GND_net), 
            .O(n906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i605_3_lut.LUT_INIT = 16'ha9a9;
    SB_LUT4 i19999_2_lut (.I0(bit_ctr[30]), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(GND_net), .O(n608));   // verilog/neopixel.v(22[26:36])
    defparam i19999_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_4_lut_adj_1692 (.I0(n708), .I1(n24488), .I2(n35702), .I3(n608), 
            .O(n35706));
    defparam i2_4_lut_adj_1692.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_2_lut_adj_1693 (.I0(bit_ctr[28]), .I1(n35706), .I2(GND_net), 
            .I3(GND_net), .O(n14452));
    defparam i1_2_lut_adj_1693.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut (.I0(n24984), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(GND_net), .O(n13425));   // verilog/neopixel.v(36[4] 116[11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i20061_2_lut_4_lut (.I0(\one_wire_N_513[9] ), .I1(\one_wire_N_513[11] ), 
            .I2(\one_wire_N_513[10] ), .I3(n15961), .O(n24782));
    defparam i20061_2_lut_4_lut.LUT_INIT = 16'hffc8;
    SB_LUT4 i31689_3_lut (.I0(n35706), .I1(n708), .I2(n35702), .I3(GND_net), 
            .O(n807));   // verilog/neopixel.v(22[26:36])
    defparam i31689_3_lut.LUT_INIT = 16'h8282;
    SB_LUT4 mod_5_i604_4_lut (.I0(n807), .I1(n838), .I2(n60), .I3(GND_net), 
            .O(n905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i604_4_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i20119_2_lut (.I0(bit_ctr[17]), .I1(n1809), .I2(GND_net), 
            .I3(GND_net), .O(n24840));
    defparam i20119_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_2_lut (.I0(n1807), .I1(n1801), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4630));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1694 (.I0(n1802), .I1(n1798), .I2(n1808), .I3(n1797), 
            .O(n24_adj_4631));
    defparam i10_4_lut_adj_1694.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1695 (.I0(n1803), .I1(n1799), .I2(n24840), .I3(n1805), 
            .O(n22_adj_4632));
    defparam i8_4_lut_adj_1695.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1696 (.I0(n1804), .I1(n24_adj_4631), .I2(n18_adj_4630), 
            .I3(n1806), .O(n26_adj_4633));
    defparam i12_4_lut_adj_1696.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1697 (.I0(n1796), .I1(n26_adj_4633), .I2(n22_adj_4632), 
            .I3(n1800), .O(n1829));
    defparam i13_4_lut_adj_1697.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1698 (.I0(n2798), .I1(n2804), .I2(n2791), .I3(n2795), 
            .O(n40_adj_4634));
    defparam i16_4_lut_adj_1698.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1699 (.I0(n2796), .I1(n2793), .I2(n2788), .I3(n2808), 
            .O(n38_adj_4635));
    defparam i14_4_lut_adj_1699.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1700 (.I0(n2789), .I1(n2800), .I2(n2803), .I3(n2805), 
            .O(n39_adj_4636));
    defparam i15_4_lut_adj_1700.LUT_INIT = 16'hfffe;
    SB_LUT4 i29117_2_lut_3_lut (.I0(n35873), .I1(one_wire_N_513[4]), .I2(n35738), 
            .I3(GND_net), .O(n35879));
    defparam i29117_2_lut_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i13_4_lut_adj_1701 (.I0(n2792), .I1(n2787), .I2(n2801), .I3(n2799), 
            .O(n37_adj_4637));
    defparam i13_4_lut_adj_1701.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_2_lut (.I0(n2786), .I1(n2797), .I2(GND_net), .I3(GND_net), 
            .O(n34_adj_4638));
    defparam i10_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i18_4_lut_adj_1702 (.I0(n2794), .I1(n2806), .I2(n2807), .I3(n2790), 
            .O(n42_adj_4639));
    defparam i18_4_lut_adj_1702.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1703 (.I0(n37_adj_4637), .I1(n39_adj_4636), .I2(n38_adj_4635), 
            .I3(n40_adj_4634), .O(n46_adj_4640));
    defparam i22_4_lut_adj_1703.LUT_INIT = 16'hfffe;
    SB_LUT4 i20261_2_lut_3_lut (.I0(n24488), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(GND_net), .O(n24982));   // verilog/neopixel.v(22[26:36])
    defparam i20261_2_lut_3_lut.LUT_INIT = 16'hbaba;
    SB_LUT4 i9_3_lut (.I0(bit_ctr[7]), .I1(n2802), .I2(n2809), .I3(GND_net), 
            .O(n33_adj_4641));
    defparam i9_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i23_4_lut_adj_1704 (.I0(n33_adj_4641), .I1(n46_adj_4640), .I2(n42_adj_4639), 
            .I3(n34_adj_4638), .O(n2819));
    defparam i23_4_lut_adj_1704.LUT_INIT = 16'hfffe;
    SB_LUT4 i34518_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n35706), .I2(bit_ctr[27]), 
            .I3(n838), .O(n17296));
    defparam i34518_3_lut_4_lut.LUT_INIT = 16'h6696;
    SB_LUT4 i36797_1_lut (.I0(n1928), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43642));
    defparam i36797_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i29087_2_lut (.I0(one_wire_N_513[4]), .I1(n35738), .I2(GND_net), 
            .I3(GND_net), .O(n35847));
    defparam i29087_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i130_4_lut (.I0(n24747), .I1(n35879), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[1] ), .O(n103));
    defparam i130_4_lut.LUT_INIT = 16'h3530;
    SB_LUT4 i1_4_lut_adj_1705 (.I0(n35873), .I1(n35847), .I2(n4), .I3(n34976), 
            .O(n34897));
    defparam i1_4_lut_adj_1705.LUT_INIT = 16'h1505;
    SB_LUT4 i1_4_lut_adj_1706 (.I0(n15961), .I1(\state[0] ), .I2(n34897), 
            .I3(n103), .O(n17155));
    defparam i1_4_lut_adj_1706.LUT_INIT = 16'h5150;
    SB_LUT4 i89_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_576 ));   // verilog/neopixel.v(35[12] 117[6])
    defparam i89_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36796_1_lut (.I0(n2918), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43641));
    defparam i36796_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i20049_2_lut (.I0(bit_ctr[3]), .I1(n3209), .I2(GND_net), .I3(GND_net), 
            .O(n24770));
    defparam i20049_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i12_4_lut_adj_1707 (.I0(n3192), .I1(n3182), .I2(n3201), .I3(n3200), 
            .O(n28_adj_4642));
    defparam i12_4_lut_adj_1707.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1708 (.I0(n3206), .I1(n3197), .I2(n3183), .I3(n3188), 
            .O(n26_adj_4643));
    defparam i10_4_lut_adj_1708.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1709 (.I0(n3208), .I1(n3199), .I2(n3196), .I3(n3185), 
            .O(n27_adj_4644));
    defparam i11_4_lut_adj_1709.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1710 (.I0(n3189), .I1(n3184), .I2(n3193), .I3(n3190), 
            .O(n25_adj_4645));
    defparam i9_4_lut_adj_1710.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut_adj_1711 (.I0(n3194), .I1(n3195), .I2(n3202), .I3(n3191), 
            .O(n20_adj_4646));
    defparam i8_4_lut_adj_1711.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1712 (.I0(n3198), .I1(n3186), .I2(n24770), .I3(n3205), 
            .O(n19_adj_4647));
    defparam i7_4_lut_adj_1712.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1713 (.I0(n25_adj_4645), .I1(n27_adj_4644), .I2(n26_adj_4643), 
            .I3(n28_adj_4642), .O(n37402));
    defparam i15_4_lut_adj_1713.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1714 (.I0(n3204), .I1(n3207), .I2(n3187), .I3(n3203), 
            .O(n21_adj_4648));
    defparam i9_4_lut_adj_1714.LUT_INIT = 16'hfffe;
    SB_LUT4 i27_4_lut (.I0(n21_adj_4648), .I1(n37402), .I2(n19_adj_4647), 
            .I3(n20_adj_4646), .O(n24824));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i20026_3_lut (.I0(\one_wire_N_513[9] ), .I1(\one_wire_N_513[11] ), 
            .I2(\one_wire_N_513[10] ), .I3(GND_net), .O(n24747));
    defparam i20026_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i234_2_lut (.I0(n24782), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n1167));   // verilog/neopixel.v(103[9] 111[12])
    defparam i234_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i1_4_lut_adj_1715 (.I0(\state[0] ), .I1(n13425), .I2(n1167), 
            .I3(\state[1] ), .O(n17203));
    defparam i1_4_lut_adj_1715.LUT_INIT = 16'haf33;
    SB_LUT4 i15_4_lut_adj_1716 (.I0(n13425), .I1(n1167), .I2(\state[1] ), 
            .I3(\state[0] ), .O(n35833));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15_4_lut_adj_1716.LUT_INIT = 16'h0535;
    SB_LUT4 i28950_2_lut_3_lut_4_lut (.I0(bit_ctr[29]), .I1(n24488), .I2(n608), 
            .I3(bit_ctr[28]), .O(n35702));
    defparam i28950_2_lut_3_lut_4_lut.LUT_INIT = 16'h5600;
    SB_LUT4 i2843_2_lut_3_lut_4_lut (.I0(bit_ctr[28]), .I1(n35706), .I2(bit_ctr[27]), 
            .I3(n35682), .O(n60));   // verilog/neopixel.v(22[26:36])
    defparam i2843_2_lut_3_lut_4_lut.LUT_INIT = 16'hff60;
    SB_LUT4 mux_665_Mux_0_i3_3_lut_3_lut (.I0(\neo_pixel_transmitter.done ), 
            .I1(start), .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_570 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_665_Mux_0_i3_3_lut_3_lut.LUT_INIT = 16'ha1a1;
    SB_LUT4 i1_3_lut_2_lut (.I0(\state[0] ), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n35021));
    defparam i1_3_lut_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut (.I0(n30047), .I1(start), .I2(\neo_pixel_transmitter.done ), 
            .I3(n15776), .O(n1164));   // verilog/neopixel.v(79[18] 99[12])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hcfdf;
    SB_LUT4 i2_2_lut_3_lut (.I0(n15776), .I1(n24922), .I2(one_wire_N_513[4]), 
            .I3(GND_net), .O(n24962));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i11_4_lut_adj_1717 (.I0(n1895), .I1(n1902), .I2(n1899), .I3(n1897), 
            .O(n26_adj_4649));
    defparam i11_4_lut_adj_1717.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1718 (.I0(n1907), .I1(bit_ctr[16]), .I2(n1909), 
            .I3(GND_net), .O(n19_adj_4650));
    defparam i4_3_lut_adj_1718.LUT_INIT = 16'heaea;
    SB_LUT4 i1_2_lut_adj_1719 (.I0(n1908), .I1(n1900), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4651));
    defparam i1_2_lut_adj_1719.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1720 (.I0(n1904), .I1(n1901), .I2(n1906), .I3(n1898), 
            .O(n24_adj_4652));
    defparam i9_4_lut_adj_1720.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1721 (.I0(n19_adj_4650), .I1(n26_adj_4649), .I2(n1905), 
            .I3(n1903), .O(n28_adj_4653));
    defparam i13_4_lut_adj_1721.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1722 (.I0(n1896), .I1(n28_adj_4653), .I2(n24_adj_4652), 
            .I3(n16_adj_4651), .O(n1928));
    defparam i14_4_lut_adj_1722.LUT_INIT = 16'hfffe;
    SB_LUT4 i36795_1_lut (.I0(n2027), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43640));
    defparam i36795_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i28949_4_lut (.I0(n15776), .I1(n30047), .I2(n4), .I3(\state[0] ), 
            .O(n24984));   // verilog/neopixel.v(36[4] 116[11])
    defparam i28949_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i3_4_lut_adj_1723 (.I0(n24698), .I1(\state[1] ), .I2(n15776), 
            .I3(n35720), .O(n36438));
    defparam i3_4_lut_adj_1723.LUT_INIT = 16'heeef;
    SB_LUT4 i2_4_lut_adj_1724 (.I0(\state[1] ), .I1(n36438), .I2(start), 
            .I3(n36198), .O(n36533));
    defparam i2_4_lut_adj_1724.LUT_INIT = 16'h8c00;
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis lattice_noprune=1, syn_instantiated=1, LSE_LINE_FILE_ID=49, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=35, LSE_RLINE=38, syn_preserve=0 */ ;   // verilog/TinyFPGA_B.v(35[10] 38[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module coms
//

module coms (clk32MHz, GND_net, rx_data, \data_in_frame[20] , \data_in_frame[8] , 
            n18251, setpoint, n36556, n18252, n18231, n18232, n18233, 
            n18234, n18235, n18236, n18237, n34167, \byte_transmit_counter[7] , 
            n34267, \byte_transmit_counter[4] , n34225, \byte_transmit_counter[5] , 
            n34421, \byte_transmit_counter[2] , n34315, \byte_transmit_counter[3] , 
            n34419, \byte_transmit_counter[1] , n43830, n18249, n18250, 
            n18247, n18248, n18245, n18246, n18243, n18244, n18241, 
            n18242, n18238, n18239, n18240, n18230, n18145, PWMLimit, 
            n18146, n18147, n18148, n18149, n18150, n18151, n34409, 
            \byte_transmit_counter[0] , n18137, n18138, n18139, n18140, 
            n18141, n18142, \data_in_frame[21] , n18155, n18156, \data_in_frame[5] , 
            n18152, n18153, n18154, n18143, n18144, n18133, \data_in_frame[24] , 
            n18134, n18135, n18136, n18126, n18127, n18128, n18129, 
            n18130, n18131, n18132, \data_in_frame[22] , \data_in_frame[4] , 
            \data_in_frame[13] , \data_in_frame[12] , \data_in_frame[3] , 
            \data_in_frame[2] , \data_in_frame[11] , \data_in_frame[1] , 
            \FRAME_MATCHER.state[3] , \FRAME_MATCHER.state[1] , n15963, 
            n13302, \data_out_frame[20] , \data_out_frame[5] , \data_out_frame[6] , 
            \data_out_frame[7] , n17934, control_mode, rx_data_ready, 
            n17933, n17932, n17931, n17930, n17929, n17928, n17927, 
            n17926, n17925, n17924, n17923, n17922, n17921, n17920, 
            n17919, \data_out_frame[19] , n17918, n17917, n17916, 
            n17915, \data_in_frame[9] , n17914, n17913, n17912, n17911, 
            \data_out_frame[18] , n17910, \data_in_frame[14][1] , n17909, 
            n35644, n17908, \data_in_frame[10] , n17907, n17906, n17905, 
            n40740, n34978, n17904, n40742, n40743, n17903, \data_out_frame[17] , 
            n17902, n40744, n37132, n16086, n17011, n35463, n35626, 
            n17901, n17900, n40747, n17899, n17898, n17897, n17896, 
            n17895, \data_out_frame[16] , n17894, n17893, n17892, 
            n17891, PIN_11_c, n17890, n17889, n17888, n17887, \data_out_frame[15] , 
            n17886, n17885, n17884, n17883, n17882, n17881, n17880, 
            n17879, \data_out_frame[14] , n17878, n17877, n17876, 
            n17875, n17874, n17873, n40746, n17872, n17871, \data_out_frame[13] , 
            n17870, n17869, n17868, n17867, n17866, n17865, n17864, 
            n17863, \data_out_frame[12] , n17862, n17861, n17860, 
            n17859, n17858, n17857, n17856, n17855, \data_out_frame[11] , 
            n17854, n17853, n17852, n17851, n17850, n17849, n17848, 
            n17847, \data_out_frame[10] , n17846, n17845, n40745, 
            n17844, n17843, n17842, n17841, n17840, n17839, \data_out_frame[9] , 
            n17838, n17837, n17836, n17835, n17834, n17833, n17832, 
            n17831, \data_out_frame[8] , n17830, n17829, n17828, n17827, 
            n17826, n17825, n17824, n17823, n17822, n17821, n17820, 
            n17819, n17818, n17817, n17816, n17815, n17814, n17813, 
            n17812, n17811, n17810, n17809, n17808, n17807, n37622, 
            n4408, n17806, n17805, n17804, n17803, n17802, n17801, 
            n17800, n17799, \data_in[3] , n17798, n17797, n17796, 
            n17795, n17794, n17793, n17792, n17791, \data_in[2] , 
            n17790, n17789, n17788, n17787, n17786, n17785, n17784, 
            n17783, \data_in[1] , n17782, n17781, n17780, n17779, 
            n17778, n17777, n17776, n17775, \data_in[0] , n17774, 
            n17773, n17772, n17771, n17770, n17769, n17768, \Ki[15] , 
            n17767, \Ki[14] , n17766, \Ki[13] , n17765, \Ki[12] , 
            n17764, \Ki[11] , n17763, \Ki[10] , n17762, \Ki[9] , 
            n17761, \Ki[8] , n17760, \Ki[7] , n17759, \Ki[6] , n17758, 
            \Ki[5] , n17757, \Ki[4] , n17756, \Ki[3] , n17755, \Ki[2] , 
            n17754, \Ki[1] , n17753, \Kp[15] , n17752, \Kp[14] , 
            n17751, \Kp[13] , n17750, \Kp[12] , n17749, \Kp[11] , 
            n17748, \Kp[10] , n17747, \Kp[9] , n17746, \Kp[8] , 
            n17745, \Kp[7] , n17744, \Kp[6] , n17743, \Kp[5] , n17742, 
            \Kp[4] , n17741, \Kp[3] , n17740, \Kp[2] , n17739, \Kp[1] , 
            n17738, gearBoxRatio, n17737, n17736, n17735, n17734, 
            n17733, n17732, n17731, n17730, n17729, n17728, n17727, 
            n17726, n17725, n17724, n17723, n17722, n17721, n17720, 
            n4593, n17719, n17718, n17717, n17716, n4387, n4397, 
            n4396, n17714, IntegralLimit, n4395, n17713, n17712, 
            n17711, n17710, n17709, n17708, n17707, n17706, n17705, 
            n17704, n17703, n17702, n17701, n17700, n17699, n4399, 
            n17698, n17697, n17696, n17695, n17694, n17693, n17692, 
            n63, n4398, n4401, n4400, n4403, n4402, n18021, n18020, 
            n18019, n18018, n18017, n18016, n18015, LED_c, n4405, 
            n4404, n4407, n4406, n18014, n17616, n3894, n788, 
            n34343, n17593, n17591, n17590, n17589, \Ki[0] , n17588, 
            \Kp[0] , n17587, n17445, \data_in_frame[6][7] , n2774, 
            n122, n15957, n2957, n5, n44342, n24190, n36526, tx_active, 
            n24918, n3, n4394, n4393, n4392, n4391, n4390, n4389, 
            \FRAME_MATCHER.state_31__N_2661[0] , n34989, n4388, n15960, 
            n63_adj_3, n35562, n15994, n4386, n4409, n5_adj_4, n17500, 
            \r_Clock_Count[3] , n17497, \r_Clock_Count[4] , n17494, 
            \r_Clock_Count[5] , n17491, \r_Clock_Count[6] , n17488, 
            \r_Clock_Count[7] , n17485, \r_Clock_Count[8] , n17513, 
            r_Bit_Index, n17510, n17506, \r_Clock_Count[1] , n17503, 
            \r_Clock_Count[2] , r_SM_Main, n17637, n313, n314, n315, 
            n316, n317, n318, n319, n320, VCC_net, n17505, tx_o, 
            tx_enable, n17607, n17606, n17605, n19670, n4, n4720, 
            n17256, n17385, n3_adj_5, n8950, n29, n17537, r_Bit_Index_adj_14, 
            n17540, n24794, \r_SM_Main[1]_adj_9 , r_Rx_Data, PIN_13_N_105, 
            \r_SM_Main[2]_adj_10 , n15851, n15740, n17250, n40690, 
            n40689, n17656, n17623, n17622, n17621, n17620, n17619, 
            n17618, n17598, n17541, n43694, n17376, n4698, n23989, 
            n4_adj_11, n4_adj_12, n4_adj_13) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input clk32MHz;
    input GND_net;
    output [7:0]rx_data;
    output [7:0]\data_in_frame[20] ;
    output [7:0]\data_in_frame[8] ;
    input n18251;
    output [23:0]setpoint;
    output n36556;
    input n18252;
    input n18231;
    input n18232;
    input n18233;
    input n18234;
    input n18235;
    input n18236;
    input n18237;
    input n34167;
    output \byte_transmit_counter[7] ;
    input n34267;
    output \byte_transmit_counter[4] ;
    input n34225;
    output \byte_transmit_counter[5] ;
    input n34421;
    output \byte_transmit_counter[2] ;
    input n34315;
    output \byte_transmit_counter[3] ;
    input n34419;
    output \byte_transmit_counter[1] ;
    input n43830;
    input n18249;
    input n18250;
    input n18247;
    input n18248;
    input n18245;
    input n18246;
    input n18243;
    input n18244;
    input n18241;
    input n18242;
    input n18238;
    input n18239;
    input n18240;
    input n18230;
    input n18145;
    output [23:0]PWMLimit;
    input n18146;
    input n18147;
    input n18148;
    input n18149;
    input n18150;
    input n18151;
    input n34409;
    output \byte_transmit_counter[0] ;
    input n18137;
    input n18138;
    input n18139;
    input n18140;
    input n18141;
    input n18142;
    output [7:0]\data_in_frame[21] ;
    input n18155;
    input n18156;
    output [7:0]\data_in_frame[5] ;
    input n18152;
    input n18153;
    input n18154;
    input n18143;
    input n18144;
    input n18133;
    output [7:0]\data_in_frame[24] ;
    input n18134;
    input n18135;
    input n18136;
    input n18126;
    input n18127;
    input n18128;
    input n18129;
    input n18130;
    input n18131;
    input n18132;
    output [7:0]\data_in_frame[22] ;
    output [7:0]\data_in_frame[4] ;
    output [7:0]\data_in_frame[13] ;
    output [7:0]\data_in_frame[12] ;
    output [7:0]\data_in_frame[3] ;
    output [7:0]\data_in_frame[2] ;
    output [7:0]\data_in_frame[11] ;
    output [7:0]\data_in_frame[1] ;
    output \FRAME_MATCHER.state[3] ;
    output \FRAME_MATCHER.state[1] ;
    output n15963;
    output n13302;
    output [7:0]\data_out_frame[20] ;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[6] ;
    output [7:0]\data_out_frame[7] ;
    input n17934;
    output [7:0]control_mode;
    output rx_data_ready;
    input n17933;
    input n17932;
    input n17931;
    input n17930;
    input n17929;
    input n17928;
    input n17927;
    input n17926;
    input n17925;
    input n17924;
    input n17923;
    input n17922;
    input n17921;
    input n17920;
    input n17919;
    output [7:0]\data_out_frame[19] ;
    input n17918;
    input n17917;
    input n17916;
    input n17915;
    output [7:0]\data_in_frame[9] ;
    input n17914;
    input n17913;
    input n17912;
    input n17911;
    output [7:0]\data_out_frame[18] ;
    input n17910;
    output \data_in_frame[14][1] ;
    input n17909;
    output n35644;
    input n17908;
    output [7:0]\data_in_frame[10] ;
    input n17907;
    input n17906;
    input n17905;
    output n40740;
    input n34978;
    input n17904;
    output n40742;
    output n40743;
    input n17903;
    output [7:0]\data_out_frame[17] ;
    input n17902;
    output n40744;
    input n37132;
    output n16086;
    output n17011;
    output n35463;
    output n35626;
    input n17901;
    input n17900;
    output n40747;
    input n17899;
    input n17898;
    input n17897;
    input n17896;
    input n17895;
    output [7:0]\data_out_frame[16] ;
    input n17894;
    input n17893;
    input n17892;
    input n17891;
    output PIN_11_c;
    input n17890;
    input n17889;
    input n17888;
    input n17887;
    output [7:0]\data_out_frame[15] ;
    input n17886;
    input n17885;
    input n17884;
    input n17883;
    input n17882;
    input n17881;
    input n17880;
    input n17879;
    output [7:0]\data_out_frame[14] ;
    input n17878;
    input n17877;
    input n17876;
    input n17875;
    input n17874;
    input n17873;
    output n40746;
    input n17872;
    input n17871;
    output [7:0]\data_out_frame[13] ;
    input n17870;
    input n17869;
    input n17868;
    input n17867;
    input n17866;
    input n17865;
    input n17864;
    input n17863;
    output [7:0]\data_out_frame[12] ;
    input n17862;
    input n17861;
    input n17860;
    input n17859;
    input n17858;
    input n17857;
    input n17856;
    input n17855;
    output [7:0]\data_out_frame[11] ;
    input n17854;
    input n17853;
    input n17852;
    input n17851;
    input n17850;
    input n17849;
    input n17848;
    input n17847;
    output [7:0]\data_out_frame[10] ;
    input n17846;
    input n17845;
    output n40745;
    input n17844;
    input n17843;
    input n17842;
    input n17841;
    input n17840;
    input n17839;
    output [7:0]\data_out_frame[9] ;
    input n17838;
    input n17837;
    input n17836;
    input n17835;
    input n17834;
    input n17833;
    input n17832;
    input n17831;
    output [7:0]\data_out_frame[8] ;
    input n17830;
    input n17829;
    input n17828;
    input n17827;
    input n17826;
    input n17825;
    input n17824;
    input n17823;
    input n17822;
    input n17821;
    input n17820;
    input n17819;
    input n17818;
    input n17817;
    input n17816;
    input n17815;
    input n17814;
    input n17813;
    input n17812;
    input n17811;
    input n17810;
    input n17809;
    input n17808;
    input n17807;
    output n37622;
    output n4408;
    input n17806;
    input n17805;
    input n17804;
    input n17803;
    input n17802;
    input n17801;
    input n17800;
    input n17799;
    output [7:0]\data_in[3] ;
    input n17798;
    input n17797;
    input n17796;
    input n17795;
    input n17794;
    input n17793;
    input n17792;
    input n17791;
    output [7:0]\data_in[2] ;
    input n17790;
    input n17789;
    input n17788;
    input n17787;
    input n17786;
    input n17785;
    input n17784;
    input n17783;
    output [7:0]\data_in[1] ;
    input n17782;
    input n17781;
    input n17780;
    input n17779;
    input n17778;
    input n17777;
    input n17776;
    input n17775;
    output [7:0]\data_in[0] ;
    input n17774;
    input n17773;
    input n17772;
    input n17771;
    input n17770;
    input n17769;
    input n17768;
    output \Ki[15] ;
    input n17767;
    output \Ki[14] ;
    input n17766;
    output \Ki[13] ;
    input n17765;
    output \Ki[12] ;
    input n17764;
    output \Ki[11] ;
    input n17763;
    output \Ki[10] ;
    input n17762;
    output \Ki[9] ;
    input n17761;
    output \Ki[8] ;
    input n17760;
    output \Ki[7] ;
    input n17759;
    output \Ki[6] ;
    input n17758;
    output \Ki[5] ;
    input n17757;
    output \Ki[4] ;
    input n17756;
    output \Ki[3] ;
    input n17755;
    output \Ki[2] ;
    input n17754;
    output \Ki[1] ;
    input n17753;
    output \Kp[15] ;
    input n17752;
    output \Kp[14] ;
    input n17751;
    output \Kp[13] ;
    input n17750;
    output \Kp[12] ;
    input n17749;
    output \Kp[11] ;
    input n17748;
    output \Kp[10] ;
    input n17747;
    output \Kp[9] ;
    input n17746;
    output \Kp[8] ;
    input n17745;
    output \Kp[7] ;
    input n17744;
    output \Kp[6] ;
    input n17743;
    output \Kp[5] ;
    input n17742;
    output \Kp[4] ;
    input n17741;
    output \Kp[3] ;
    input n17740;
    output \Kp[2] ;
    input n17739;
    output \Kp[1] ;
    input n17738;
    output [23:0]gearBoxRatio;
    input n17737;
    input n17736;
    input n17735;
    input n17734;
    input n17733;
    input n17732;
    input n17731;
    input n17730;
    input n17729;
    input n17728;
    input n17727;
    input n17726;
    input n17725;
    input n17724;
    input n17723;
    input n17722;
    input n17721;
    input n17720;
    output n4593;
    input n17719;
    input n17718;
    input n17717;
    input n17716;
    output n4387;
    output n4397;
    output n4396;
    input n17714;
    output [23:0]IntegralLimit;
    output n4395;
    input n17713;
    input n17712;
    input n17711;
    input n17710;
    input n17709;
    input n17708;
    input n17707;
    input n17706;
    input n17705;
    input n17704;
    input n17703;
    input n17702;
    input n17701;
    input n17700;
    input n17699;
    output n4399;
    input n17698;
    input n17697;
    input n17696;
    input n17695;
    input n17694;
    input n17693;
    input n17692;
    output n63;
    output n4398;
    output n4401;
    output n4400;
    output n4403;
    output n4402;
    input n18021;
    input n18020;
    input n18019;
    input n18018;
    input n18017;
    input n18016;
    input n18015;
    output LED_c;
    output n4405;
    output n4404;
    output n4407;
    output n4406;
    input n18014;
    input n17616;
    output n3894;
    output n788;
    input n34343;
    input n17593;
    input n17591;
    input n17590;
    input n17589;
    output \Ki[0] ;
    input n17588;
    output \Kp[0] ;
    input n17587;
    input n17445;
    output \data_in_frame[6][7] ;
    output n2774;
    output n122;
    output n15957;
    output n2957;
    output n5;
    output n44342;
    output n24190;
    output n36526;
    output tx_active;
    output n24918;
    output n3;
    output n4394;
    output n4393;
    output n4392;
    output n4391;
    output n4390;
    output n4389;
    output \FRAME_MATCHER.state_31__N_2661[0] ;
    output n34989;
    output n4388;
    output n15960;
    output n63_adj_3;
    output n35562;
    output n15994;
    output n4386;
    output n4409;
    output n5_adj_4;
    input n17500;
    output \r_Clock_Count[3] ;
    input n17497;
    output \r_Clock_Count[4] ;
    input n17494;
    output \r_Clock_Count[5] ;
    input n17491;
    output \r_Clock_Count[6] ;
    input n17488;
    output \r_Clock_Count[7] ;
    input n17485;
    output \r_Clock_Count[8] ;
    input n17513;
    output [2:0]r_Bit_Index;
    input n17510;
    input n17506;
    output \r_Clock_Count[1] ;
    input n17503;
    output \r_Clock_Count[2] ;
    output [2:0]r_SM_Main;
    input n17637;
    output n313;
    output n314;
    output n315;
    output n316;
    output n317;
    output n318;
    output n319;
    output n320;
    input VCC_net;
    output n17505;
    output tx_o;
    output tx_enable;
    input n17607;
    input n17606;
    input n17605;
    output n19670;
    output n4;
    output n4720;
    output n17256;
    output n17385;
    output n3_adj_5;
    output n8950;
    output n29;
    input n17537;
    output [2:0]r_Bit_Index_adj_14;
    input n17540;
    input n24794;
    output \r_SM_Main[1]_adj_9 ;
    output r_Rx_Data;
    input PIN_13_N_105;
    output \r_SM_Main[2]_adj_10 ;
    output n15851;
    output n15740;
    output n17250;
    output n40690;
    output n40689;
    input n17656;
    input n17623;
    input n17622;
    input n17621;
    input n17620;
    input n17619;
    input n17618;
    input n17598;
    input n17541;
    output n43694;
    output n17376;
    output n4698;
    output n23989;
    output n4_adj_11;
    output n4_adj_12;
    output n4_adj_13;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire LED_c /* synthesis SET_AS_NETWORK=LED_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(4[10:13])
    
    wire n30588;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(95[12:25])
    
    wire n35173, n6, n30586, n17988;
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(95[12:25])
    
    wire n18092, n18091, n18090, n18089, n18088, n18087, n18086, 
        n18085;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(95[12:25])
    
    wire n18084, n18083, n18082;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(114[11:12])
    
    wire n161, n27884, n18081, n18080, n35357, n35487, n6_adj_4259, 
        n17987, n17986, n2, n3_c, n8, n35006, n18094, n18079, 
        n18078, n18077;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(95[12:25])
    
    wire n17985, n17984, n18076, n18075, n18101, n17998, n17997;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(95[12:25])
    
    wire n17996, n17995, n17994, n18100, n18099, n17993, n17992, 
        n18098, n13414, n31, n15950, n17991, n18288;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(101[12:33])
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(111[11:16])
    
    wire n8_adj_4260, n18122;
    wire [7:0]\data_in_frame[23] ;   // verilog/coms.v(95[12:25])
    
    wire n18123, n18102, n18103, n18104, n17983, n17982, n18093, 
        n18095, n17981, n17990, n18124, n18125, n17980, n18118, 
        n18119, n18120, n18121, n18116, n18117, n18114, n18115, 
        n18112, n18113, n18110, n18111, n18108, n18109, n17979, 
        n18105, n18106, n18107, n18096, n18097, n17978, n17977, 
        n17976, n17975, n17974, n17973, n17972, n17971, n17970, 
        n17969, n17968, n18039, n18038, n18037, n18036, n17967, 
        n17966, n17965, n18035, n18034, n18033, n18032, n18031, 
        n17964, n17963, n17962, n18048;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(95[12:25])
    
    wire n17961, n17960, n17959, n17958, n17957, n18030, n18029, 
        n18028, n18027, n17956, n17955, n17954, n17953, n17952, 
        n17951, n17950, n17949, n17948, n17947, n17946, n17945, 
        n17944, n17943, n17942, n17941;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(95[12:25])
    
    wire n17940, n17939, n17938, n18026, n38543, n30, n34891, 
        n28, n29_c, n38681, n38680;
    wire [7:0]tx_data;   // verilog/coms.v(104[13:20])
    
    wire n27, n18025;
    wire [31:0]\FRAME_MATCHER.state_31__N_2725 ;
    
    wire n15886, n34898, n38526, n13013, n18074;
    wire [7:0]\data_out_frame[21] ;   // verilog/coms.v(96[12:26])
    
    wire n19, n6_adj_4261, n5_c;
    wire [7:0]\data_out_frame[22] ;   // verilog/coms.v(96[12:26])
    
    wire n38653, n43712, n38654, n18073, n40522, n38661, n18072, 
        n38663, n43772, n43766, n38662, n17937, n17936, n17935;
    wire [0:0]n3332;
    wire [2:0]r_SM_Main_2__N_3585;
    
    wire n35671, \FRAME_MATCHER.rx_data_ready_prev , n18071, n18070, 
        n35300, n30523, n15609, n6_adj_4262, n18024, n36755, n37377, 
        Kp_23__N_805, n38678, n38677, n35558, n35590, n16777, n35438, 
        n35360, n16386, n35543, n18040, n18023, n18047, n18069;
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(95[12:25])
    
    wire n18068, n18046, n35182, n16156, n35499, n20, n35413, 
        n35110, n30671, n35581, n19_adj_4263, n35391, n35154, n16044, 
        n21, n15568, n35578, n35327, n35454, n16, n30578, n35629, 
        n35224, n17, n18067, n24966, n24738, n101, n5_adj_4264, 
        n36982, n4498, n16034, n37006, n37597, n16883, n12, n16272, 
        n35354, n31482, n7, n35227, Kp_23__N_1186, n35518, n35294, 
        n16642, n35533, n35385, n16142, n35122, n16552, n16645, 
        n16464, n16782, n16231, n35167, n35617, n30529, n35135, 
        n14, n35555;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(95[12:25])
    
    wire n15, n37527, n16835, n11, n36431, n31528, n30677, n35347, 
        n10, n35276, n35508, n8_adj_4265, n37028, n27926, n40622, 
        n27925, \FRAME_MATCHER.i_31__N_2624 , n18045, n18044, n14_adj_4266, 
        n18043, n27924, n27923, n18042, n38675, n38674, n27922, 
        n10_adj_4267, n36306, n31558, n30683, n30689, n35147, n35394, 
        n35370, n35144, n31571, n12_adj_4268, n35552, n30592, n35367, 
        n30807, n35341, n16202, n35493, Kp_23__N_1802, n35602, n10_adj_4269, 
        n35546, n35364, n15_adj_4270, n35273, n35218, n21_adj_4271, 
        n30812, n35599, n20_adj_4272, n18, n35157, n24, n35176, 
        n37548, n31470, n12_adj_4273, n18_adj_4274, n35511, n35037, 
        n30721, n14_adj_4275, n35515, n35259, n17_adj_4276, n35410, 
        n13, n9, n17023, n11_adj_4277, n31460, n35407, n8_adj_4278, 
        n16838, n36572, n35344, n24_adj_4279, n22, n36394, n38515, 
        n35466, n21_adj_4280, n35279, n31474, n36878, n37403, n14_adj_4281, 
        n36317, n37411, n27921, n37080, n37572, n18041, n20_adj_4282, 
        n19_adj_4283, n30_adj_4284, n25, n31_adj_4285, n26, n35101, 
        n35051, n16494, n15531, n35170, n16399, n4462, n35783, 
        n37191, n34998, n35416, n27920, n36436, tx_transmit_N_3482, 
        n35104, n16953, n16555, n6_adj_4286, n6_adj_4287, n17042, 
        n16038, n5_adj_4288, n35048, n35044, n6_adj_4289, Kp_23__N_1003, 
        n35138, n8_adj_4290, n18_adj_4291, n24_adj_4292, n22_adj_4293, 
        n35268, n26_adj_4294, n37530, n35441, n35098, n35245, n30669, 
        n6_adj_4295, Kp_23__N_949, n6_adj_4296, n14_adj_4297, n9_adj_4298, 
        n16360, n16115, n37247, n16876, n16_adj_4299, n22_adj_4300, 
        n20_adj_4301, n24_adj_4302, n4385, n24968, n24910, n12_adj_4303, 
        n24686, n35536, n6_adj_4304, n14_adj_4305, n30584, n31464, 
        n16345, n4_c, n36548, n16029, n35426, n35256, n28_adj_4306, 
        n32, n16006, n35221, n38569, n9_adj_4307, n6_adj_4308, n4_adj_4309, 
        n16445, n16716, n16239, n10_adj_4310, n35151, n35584, n37560, 
        n36894, n31480, n35566, n35587, n16714, n16772, n30582, 
        n10_adj_4311, n35638, n86, n8_adj_4312, n16184, n35318, 
        n36368, n35521, n35297, n31017, n35230, n35376, n8_adj_4313, 
        n6_adj_4314, n18022, n63_c, n63_adj_4315, n10389;
    wire [31:0]n23;
    
    wire n70, n67, n34465, n7_adj_4317, n7_adj_4318, n34451, n34463, 
        n34461, n38672, n38671, n7_adj_4319, n34459, n8_adj_4320, 
        n34457, n34469, n7_adj_4321, n34449, n7_adj_4322, n43805, 
        n43808, n43799, n43802, n43793, n43796, n23914, n23912, 
        n2_adj_4323, n3_adj_4324, n18000, n34447, n34445, n34455, 
        n34443, n34467, n34441, n2_adj_4325, n3_adj_4326, n34429, 
        n2_adj_4327, n3_adj_4328, n2_adj_4329, n3_adj_4330, n2_adj_4331, 
        n3_adj_4332, n2_adj_4333, n3_adj_4334, n2_adj_4335, n3_adj_4336, 
        n2_adj_4337, n3_adj_4338, n2_adj_4339, n3_adj_4340, n2_adj_4341, 
        n3_adj_4342, n2_adj_4343, n3_adj_4344, n2_adj_4345, n3_adj_4346, 
        n2_adj_4347, n3_adj_4348, n2_adj_4349, n3_adj_4350, n2_adj_4351, 
        n3_adj_4352, n2_adj_4353, n3_adj_4354, n2_adj_4355, n3_adj_4356, 
        n2_adj_4357, n3_adj_4358, n2_adj_4359, n3_adj_4360, n2_adj_4361, 
        n3_adj_4362, n2_adj_4363, n3_adj_4364, n2_adj_4365, n3_adj_4366, 
        n2_adj_4367, n3_adj_4368, n2_adj_4369, n3_adj_4370, n2_adj_4371, 
        n3_adj_4372, n2_adj_4373, n3_adj_4374, n2_adj_4375, n3_adj_4376, 
        n2_adj_4377, n3_adj_4378, n2_adj_4379, n3_adj_4380, n2_adj_4381, 
        n3_adj_4382, n2_adj_4383, n3_adj_4384, n34453, n36265, n17205, 
        n36416, n37044, n36758, n36181, n36199, n37556, n36904, 
        n35353, n35271, n36143, n36260, n35383, n36345, n36347, 
        n37510, n34439, n17348, n34927, n37152, n34329, n44032, 
        n34437, n34333, n10_adj_4385, n34431, n34331, n34433, n34397, 
        n34435, n34395, n34393, n34391, n34335, n34401, n34389, 
        n34339, n34387, n34351, n34385, n34383, n24679, n24681, 
        n8_adj_4386, n34381, n8_adj_4387, n34349, n34347, n34345, 
        n34273, n34337, n34341, n34379, n8_adj_4388, n8_adj_4389, 
        n34323, n15_adj_4390, n46, n1, n43787, n8_adj_4391, n34984, 
        n18006, n18007, n18008, n18009, n18010, n18011, n18012, 
        n18013, n6_adj_4392, n37642, n2058, n9_adj_4393, n36539, 
        n15939, n37335, n18066, n15759, n15848, n16_adj_4394, n17_adj_4395, 
        n24712, n18054, n18055, n18065, n15858, n16_adj_4396, n17_adj_4397, 
        n18056, n18057, n18058, n18059, n18060, n18061, n15460, 
        n37314, n31476, n18064, n18063, n18062, n35082, n31530, 
        n4_adj_4398, n8_adj_4399, n15845, n35575, n43790, n27914, 
        n27913, n27912, n17999, n4_adj_4400, n15722, n9_adj_4401, 
        n12_adj_4402, n19_adj_4403, n40680, n43781, n9015, n44, 
        n35388, n42, n43, n41, n7_adj_4404, n40, n17_adj_4405, 
        n16_adj_4406, n43784, n39, n50, n45, n15765, n15992, n18005, 
        n18004, n18003, n17592, n27911, n27910, n17989, n27909, 
        n27908, n27907, n27906, n27905, n8_adj_4407, n27904, n6_adj_4408, 
        n27903, n27902, n27901, n27900, n27899, n27898, n27897, 
        n27896, n27895, n27894, n31118, n35249, n27893, n27892, 
        n10_adj_4409, n27891, n14_adj_4410, n27890, n10_adj_4411, 
        n31457, n35067, n38564, n9_adj_4412, n27889, n18002, n18001, 
        n18053, n18052, n18051, n18050, n27888, n38538, n27887, 
        n27886, n18049, n21_adj_4413, n27885, n20_adj_4414, n24_adj_4415, 
        n43775, n23947, n43_adj_4416, n24684, n43778, n43769, n43763, 
        n43757, n43760, n35641, n16812, n35185, n30512, n6_adj_4418, 
        n43751, n43754, n43745, n43748, n43739, n43742, n30704, 
        n14_adj_4419, n43733, n43736, n43727, n43730, n43721, n43724, 
        n18_adj_4420, n43715, n43718, n24_adj_4421, n43709, n22_adj_4422, 
        n16870, n35125, n16587, n6_adj_4423, n35057, n35651, n35188, 
        n10_adj_4424, n34995, n38499, n10_adj_4425, n35429, n1286, 
        n16937, n30598, n35422, n43703, n35490, n35141, n14107, 
        n35654, n16214, n35565, n35635, n35212, n43706, n35475, 
        n35596, n8_adj_4426, n30558, n26_adj_4427, n43697, n6_adj_4428, 
        n35530, n16_adj_4429, n7_adj_4430, n8_adj_4431, n43700, n25_adj_4433, 
        n35432, n38666, n38665, n30545, n31254, n35107, n31610, 
        n30653, n31455, n35081, n16566, n35285, n35079, n30516, 
        n30667, n6_adj_4434, n35524, n35525, n31518, n5_adj_4435, 
        n15861, n7_adj_4436, n14_adj_4437, n6_adj_4438, n10_adj_4439, 
        n35091, n6_adj_4440, n38669, n38668, n12_adj_4442, n15958, 
        n41108, n5_adj_4443, n38649, n38651, n43670, n43664, n38650, 
        n19_adj_4444, n41104, n5_adj_4445, n38695, n38696, n38679, 
        n43682, n43676, n16246, n14_adj_4446, n19_adj_4447, n41099, 
        n5_adj_4448, n38692, n38693, n38676, n43688, n19_adj_4449, 
        n6_adj_4450, n5_adj_4451, n38689, n38690, n38673, n35164, 
        n31068, n35472, n19_adj_4452, n6_adj_4453, Kp_23__N_1768, 
        n5_adj_4454, n38686, n38687, n38670, n15_adj_4455, n10_adj_4456, 
        n16659, n43685, n19_adj_4457, n6_adj_4458, n5_adj_4459, n38683, 
        n38684, n38667, n14_adj_4460, n37297, n19_adj_4461, n6_adj_4462, 
        n5_adj_4463, n38656, n38657, n43679, n38664, n8_adj_4464, 
        n12_adj_4465, n8_adj_4466, n16486, n98, n30730, n96, n97, 
        n95, n35309, n90, n88, n89, n87, n94, n35303, n35315, 
        n92, n93, n91, n99, n110, n108, n109, n107, n13144, 
        n13181, n65, n35746, n30622, n6_adj_4467;
    wire [31:0]\FRAME_MATCHER.state_31__N_2661 ;
    
    wire n5_adj_4468, n5_adj_4469, n35129, n35336, n12_adj_4470, n35382, 
        n35351, n14129, n16020, n10_adj_4471, n7_adj_4472, n35549, 
        n22_adj_4473, n20_adj_4474, n24_adj_4475, n43673, n6_adj_4476, 
        n35502, n6_adj_4477, n31552, n30681, n35614, n6_adj_4478, 
        n31504, n6_adj_4479, n35070, n31140, n31595, n16163, n35033, 
        n18_adj_4480, n17033, n30_adj_4481, n35505, n28_adj_4482, 
        n35288, n17080, n29_adj_4483, n35397, n35262, n27_adj_4484, 
        n12_adj_4485, n6_adj_4486, n43667, n43661, n31510, n12_adj_4487, 
        n35478, n35196, n16_adj_4488, n35379, n35265, n16949, n35060, 
        n35404, n35647, n52, n35484, n59, n35608, n40_adj_4489, 
        n35448, n35527, n38, n35236, n31478, n39_adj_4490, n37, 
        n35400, n35306, n35064, n56, n54, n35054, n35460, n55, 
        n53, n58, n64, n16729, n57, n65_adj_4491, n37570, n42_adj_4492, 
        n46_adj_4493, n41_adj_4494, n35321, n35322, n10_adj_4495, 
        n31178, n35611, n35330, n11_adj_4496, n13_adj_4497, n35041, 
        n35113, n6_adj_4498, n37407, n16982, n30618, n35119, n7_adj_4499, 
        n16530, n1608, n35161, n16806, n35481, n35593, n35076, 
        n1205, n26_adj_4500, n35572, n30_adj_4501, n34, n35657, 
        n29_adj_4502, n35469, n10_adj_4503, n17071, n35209, n14_adj_4504, 
        n35206, n14123, n10_adj_4505, n14180, n35291, n35457, n10_adj_4506, 
        n35324, n14_adj_4507, n30630, n6_adj_4509, n35451, n35132, 
        n10_adj_4510, n16482, n35242, n35496, n35605, n10_adj_4511, 
        n16821, n16252, n12_adj_4512, n10_adj_4513, n35032, n15_adj_4514;
    
    SB_LUT4 i4_4_lut (.I0(n30588), .I1(\data_in_frame[19] [7]), .I2(n35173), 
            .I3(n6), .O(n30586));
    defparam i4_4_lut.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(clk32MHz), 
           .D(n17988));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(clk32MHz), 
           .D(n18092));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(clk32MHz), 
           .D(n18091));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(clk32MHz), 
           .D(n18090));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(clk32MHz), 
           .D(n18089));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(clk32MHz), 
           .D(n18088));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(clk32MHz), 
           .D(n18087));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(clk32MHz), 
           .D(n18086));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(clk32MHz), 
           .D(n18085));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(clk32MHz), 
           .D(n18084));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(clk32MHz), 
           .D(n18083));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(clk32MHz), 
           .D(n18082));   // verilog/coms.v(127[12] 295[6])
    SB_CARRY add_44_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n27884));
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(clk32MHz), 
           .D(n18081));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(clk32MHz), 
           .D(n18080));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut (.I0(n35357), .I1(n35487), .I2(GND_net), .I3(GND_net), 
            .O(n6_adj_4259));
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(clk32MHz), 
           .D(n17987));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(clk32MHz), 
           .D(n17986));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(clk32MHz), 
            .D(n2), .S(n3_c));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13355_3_lut_4_lut (.I0(n8), .I1(n35006), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n18094));
    defparam i13355_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(clk32MHz), 
           .D(n18079));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(clk32MHz), 
           .D(n18078));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(clk32MHz), 
           .D(n18077));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(clk32MHz), 
           .D(n17985));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(clk32MHz), 
           .D(n17984));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(clk32MHz), 
           .D(n18076));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(clk32MHz), 
           .D(n18075));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13362_3_lut_4_lut (.I0(n8), .I1(n35006), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n18101));
    defparam i13362_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(clk32MHz), 
           .D(n17998));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(clk32MHz), 
           .D(n17997));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(clk32MHz), 
           .D(n17996));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(clk32MHz), 
           .D(n17995));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(clk32MHz), 
           .D(n17994));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13361_3_lut_4_lut (.I0(n8), .I1(n35006), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n18100));
    defparam i13361_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13360_3_lut_4_lut (.I0(n8), .I1(n35006), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n18099));
    defparam i13360_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(clk32MHz), 
           .D(n17993));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(clk32MHz), 
           .D(n17992));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13359_3_lut_4_lut (.I0(n8), .I1(n35006), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n18098));
    defparam i13359_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF setpoint__i22 (.Q(setpoint[22]), .C(clk32MHz), .D(n18251));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i2_3_lut (.I0(n13414), .I1(n31), .I2(n15950), .I3(GND_net), 
            .O(n36556));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_DFF setpoint__i23 (.Q(setpoint[23]), .C(clk32MHz), .D(n18252));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(clk32MHz), 
           .D(n17991));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i2 (.Q(setpoint[2]), .C(clk32MHz), .D(n18231));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i3 (.Q(setpoint[3]), .C(clk32MHz), .D(n18232));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i4 (.Q(setpoint[4]), .C(clk32MHz), .D(n18233));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i5 (.Q(setpoint[5]), .C(clk32MHz), .D(n18234));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i6 (.Q(setpoint[6]), .C(clk32MHz), .D(n18235));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i7 (.Q(setpoint[7]), .C(clk32MHz), .D(n18236));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i8 (.Q(setpoint[8]), .C(clk32MHz), .D(n18237));   // verilog/coms.v(127[12] 295[6])
    SB_DFF byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(clk32MHz), 
           .D(n18288));   // verilog/coms.v(127[12] 295[6])
    SB_DFF byte_transmit_counter_i0_i7 (.Q(\byte_transmit_counter[7] ), .C(clk32MHz), 
           .D(n34167));   // verilog/coms.v(127[12] 295[6])
    SB_DFF byte_transmit_counter_i0_i4 (.Q(\byte_transmit_counter[4] ), .C(clk32MHz), 
           .D(n34267));   // verilog/coms.v(127[12] 295[6])
    SB_DFF byte_transmit_counter_i0_i5 (.Q(\byte_transmit_counter[5] ), .C(clk32MHz), 
           .D(n34225));   // verilog/coms.v(127[12] 295[6])
    SB_DFF byte_transmit_counter_i0_i2 (.Q(\byte_transmit_counter[2] ), .C(clk32MHz), 
           .D(n34421));   // verilog/coms.v(127[12] 295[6])
    SB_DFF byte_transmit_counter_i0_i3 (.Q(\byte_transmit_counter[3] ), .C(clk32MHz), 
           .D(n34315));   // verilog/coms.v(127[12] 295[6])
    SB_DFF byte_transmit_counter_i0_i1 (.Q(\byte_transmit_counter[1] ), .C(clk32MHz), 
           .D(n34419));   // verilog/coms.v(127[12] 295[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state [2]), .C(clk32MHz), 
           .D(n43830));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i20 (.Q(setpoint[20]), .C(clk32MHz), .D(n18249));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 equal_116_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4260));   // verilog/coms.v(154[7:23])
    defparam equal_116_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_DFF setpoint__i21 (.Q(setpoint[21]), .C(clk32MHz), .D(n18250));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i18 (.Q(setpoint[18]), .C(clk32MHz), .D(n18247));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i19 (.Q(setpoint[19]), .C(clk32MHz), .D(n18248));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i16 (.Q(setpoint[16]), .C(clk32MHz), .D(n18245));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i17 (.Q(setpoint[17]), .C(clk32MHz), .D(n18246));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i14 (.Q(setpoint[14]), .C(clk32MHz), .D(n18243));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i15 (.Q(setpoint[15]), .C(clk32MHz), .D(n18244));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i12 (.Q(setpoint[12]), .C(clk32MHz), .D(n18241));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i13 (.Q(setpoint[13]), .C(clk32MHz), .D(n18242));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i9 (.Q(setpoint[9]), .C(clk32MHz), .D(n18238));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i10 (.Q(setpoint[10]), .C(clk32MHz), .D(n18239));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i11 (.Q(setpoint[11]), .C(clk32MHz), .D(n18240));   // verilog/coms.v(127[12] 295[6])
    SB_DFF setpoint__i1 (.Q(setpoint[1]), .C(clk32MHz), .D(n18230));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 equal_101_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8));   // verilog/coms.v(154[7:23])
    defparam equal_101_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(clk32MHz), .D(n18145));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(clk32MHz), .D(n18146));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(clk32MHz), .D(n18147));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(clk32MHz), .D(n18148));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(clk32MHz), .D(n18149));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(clk32MHz), .D(n18150));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(clk32MHz), .D(n18151));   // verilog/coms.v(127[12] 295[6])
    SB_DFF byte_transmit_counter_i0_i0 (.Q(\byte_transmit_counter[0] ), .C(clk32MHz), 
           .D(n34409));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(clk32MHz), .D(n18137));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(clk32MHz), .D(n18138));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(clk32MHz), .D(n18139));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(clk32MHz), .D(n18140));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(clk32MHz), .D(n18141));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(clk32MHz), .D(n18142));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i189 (.Q(\data_in_frame[23] [4]), .C(clk32MHz), 
           .D(n18122));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i190 (.Q(\data_in_frame[23] [5]), .C(clk32MHz), 
           .D(n18123));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(clk32MHz), 
           .D(n18098));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(clk32MHz), 
           .D(n18099));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(clk32MHz), 
           .D(n18100));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(clk32MHz), 
           .D(n18101));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(clk32MHz), 
           .D(n18102));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(clk32MHz), 
           .D(n18103));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(clk32MHz), 
           .D(n18104));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(clk32MHz), 
           .D(n17983));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(clk32MHz), 
           .D(n17982));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(clk32MHz), 
           .D(n18093));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(clk32MHz), 
           .D(n18094));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(clk32MHz), 
           .D(n18095));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(clk32MHz), .D(n18155));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(clk32MHz), .D(n18156));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(clk32MHz), 
           .D(n17981));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(clk32MHz), .D(n18152));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(clk32MHz), .D(n18153));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(clk32MHz), .D(n18154));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(clk32MHz), .D(n18143));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(clk32MHz), .D(n18144));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i200 (.Q(\data_in_frame[24] [7]), .C(clk32MHz), 
           .D(n18133));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(clk32MHz), .D(n18134));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(clk32MHz), .D(n18135));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(clk32MHz), .D(n18136));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(clk32MHz), 
           .D(n17990));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i191 (.Q(\data_in_frame[23] [6]), .C(clk32MHz), 
           .D(n18124));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i192 (.Q(\data_in_frame[23] [7]), .C(clk32MHz), 
           .D(n18125));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i193 (.Q(\data_in_frame[24] [0]), .C(clk32MHz), 
           .D(n18126));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i194 (.Q(\data_in_frame[24] [1]), .C(clk32MHz), 
           .D(n18127));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i195 (.Q(\data_in_frame[24] [2]), .C(clk32MHz), 
           .D(n18128));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i196 (.Q(\data_in_frame[24] [3]), .C(clk32MHz), 
           .D(n18129));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i197 (.Q(\data_in_frame[24] [4]), .C(clk32MHz), 
           .D(n18130));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i198 (.Q(\data_in_frame[24] [5]), .C(clk32MHz), 
           .D(n18131));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i199 (.Q(\data_in_frame[24] [6]), .C(clk32MHz), 
           .D(n18132));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(clk32MHz), 
           .D(n17980));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i185 (.Q(\data_in_frame[23] [0]), .C(clk32MHz), 
           .D(n18118));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i186 (.Q(\data_in_frame[23] [1]), .C(clk32MHz), 
           .D(n18119));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i187 (.Q(\data_in_frame[23] [2]), .C(clk32MHz), 
           .D(n18120));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i188 (.Q(\data_in_frame[23] [3]), .C(clk32MHz), 
           .D(n18121));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i183 (.Q(\data_in_frame[22] [6]), .C(clk32MHz), 
           .D(n18116));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i184 (.Q(\data_in_frame[22] [7]), .C(clk32MHz), 
           .D(n18117));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i181 (.Q(\data_in_frame[22] [4]), .C(clk32MHz), 
           .D(n18114));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i182 (.Q(\data_in_frame[22] [5]), .C(clk32MHz), 
           .D(n18115));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i179 (.Q(\data_in_frame[22] [2]), .C(clk32MHz), 
           .D(n18112));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i180 (.Q(\data_in_frame[22] [3]), .C(clk32MHz), 
           .D(n18113));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i177 (.Q(\data_in_frame[22] [0]), .C(clk32MHz), 
           .D(n18110));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i178 (.Q(\data_in_frame[22] [1]), .C(clk32MHz), 
           .D(n18111));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(clk32MHz), 
           .D(n18108));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(clk32MHz), 
           .D(n18109));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(clk32MHz), 
           .D(n17979));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(clk32MHz), 
           .D(n18105));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(clk32MHz), 
           .D(n18106));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(clk32MHz), 
           .D(n18107));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(clk32MHz), 
           .D(n18096));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(clk32MHz), 
           .D(n18097));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(clk32MHz), 
           .D(n17978));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(clk32MHz), 
           .D(n17977));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(clk32MHz), 
           .D(n17976));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(clk32MHz), 
           .D(n17975));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(clk32MHz), 
           .D(n17974));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(clk32MHz), 
           .D(n17973));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(clk32MHz), 
           .D(n17972));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(clk32MHz), 
           .D(n17971));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(clk32MHz), 
           .D(n17970));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(clk32MHz), 
           .D(n17969));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(clk32MHz), 
           .D(n17968));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(clk32MHz), 
           .D(n18039));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(clk32MHz), 
           .D(n18038));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(clk32MHz), 
           .D(n18037));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(clk32MHz), 
           .D(n18036));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(clk32MHz), 
           .D(n17967));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(clk32MHz), 
           .D(n17966));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(clk32MHz), 
           .D(n17965));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(clk32MHz), 
           .D(n18035));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(clk32MHz), 
           .D(n18034));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(clk32MHz), 
           .D(n18033));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(clk32MHz), 
           .D(n18032));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(clk32MHz), 
           .D(n18031));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(clk32MHz), 
           .D(n17964));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(clk32MHz), 
           .D(n17963));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(clk32MHz), 
           .D(n17962));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(clk32MHz), 
           .D(n18048));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(clk32MHz), 
           .D(n17961));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(clk32MHz), 
           .D(n17960));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(clk32MHz), 
           .D(n17959));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(clk32MHz), 
           .D(n17958));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(clk32MHz), 
           .D(n17957));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(clk32MHz), 
           .D(n18030));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(clk32MHz), 
           .D(n18029));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(clk32MHz), 
           .D(n18028));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(clk32MHz), 
           .D(n18027));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(clk32MHz), 
           .D(n17956));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(clk32MHz), 
           .D(n17955));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(clk32MHz), 
           .D(n17954));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(clk32MHz), 
           .D(n17953));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(clk32MHz), 
           .D(n17952));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(clk32MHz), 
           .D(n17951));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(clk32MHz), 
           .D(n17950));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(clk32MHz), 
           .D(n17949));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(clk32MHz), 
           .D(n17948));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(clk32MHz), 
           .D(n17947));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(clk32MHz), 
           .D(n17946));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(clk32MHz), 
           .D(n17945));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(clk32MHz), 
           .D(n17944));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(clk32MHz), 
           .D(n17943));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(clk32MHz), 
           .D(n17942));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(clk32MHz), 
           .D(n17941));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(clk32MHz), 
           .D(n17940));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(clk32MHz), 
           .D(n17939));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(clk32MHz), 
           .D(n17938));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(clk32MHz), 
           .D(n18026));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i31774_2_lut (.I0(\data_in_frame[1] [7]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n38543));
    defparam i31774_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut (.I0(n38543), .I1(\data_in_frame[2] [3]), .I2(\data_in_frame[2] [0]), 
            .I3(\data_in_frame[2] [6]), .O(n30));
    defparam i13_4_lut.LUT_INIT = 16'h0010;
    SB_LUT4 i11_4_lut (.I0(n34891), .I1(\data_in_frame[2] [4]), .I2(\data_in_frame[2] [1]), 
            .I3(\data_in_frame[1] [5]), .O(n28));
    defparam i11_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i12_4_lut (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(\data_in_frame[2] [5]), .I3(\data_in_frame[2] [7]), .O(n29_c));
    defparam i12_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut (.I0(\byte_transmit_counter[4] ), 
            .I1(\byte_transmit_counter[3] ), .I2(n38681), .I3(n38680), 
            .O(tx_data[6]));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i10_4_lut (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[1] [3]), .O(n27));
    defparam i10_4_lut.LUT_INIT = 16'h8000;
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(clk32MHz), 
           .D(n18025));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i16_4_lut (.I0(n27), .I1(n29_c), .I2(n28), .I3(n30), .O(\FRAME_MATCHER.state_31__N_2725 [3]));
    defparam i16_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_997 (.I0(\FRAME_MATCHER.state[3] ), .I1(n15886), 
            .I2(GND_net), .I3(GND_net), .O(n34898));
    defparam i1_2_lut_adj_997.LUT_INIT = 16'h2222;
    SB_LUT4 i31758_2_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n38526));
    defparam i31758_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut (.I0(\FRAME_MATCHER.state[1] ), .I1(n34898), .I2(n38526), 
            .I3(\FRAME_MATCHER.state [0]), .O(n13013));
    defparam i1_4_lut.LUT_INIT = 16'hccce;
    SB_LUT4 i3_4_lut (.I0(\FRAME_MATCHER.state_31__N_2725 [3]), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(n15963), .I3(n13013), .O(n13302));   // verilog/coms.v(127[12] 295[6])
    defparam i3_4_lut.LUT_INIT = 16'h0800;
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(clk32MHz), 
           .D(n18074));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i19_3_lut (.I0(\data_out_frame[20] [0]), 
            .I1(\data_out_frame[21] [0]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i6_4_lut (.I0(\data_out_frame[5] [0]), 
            .I1(\byte_transmit_counter[0] ), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[1] ), .O(n6_adj_4261));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i6_4_lut.LUT_INIT = 16'hb0bc;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i5_3_lut (.I0(\data_out_frame[6] [0]), 
            .I1(\data_out_frame[7] [0]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_c));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31807_4_lut (.I0(n19), .I1(\data_out_frame[22] [0]), .I2(\byte_transmit_counter[1] ), 
            .I3(\byte_transmit_counter[0] ), .O(n38653));
    defparam i31807_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31808_3_lut (.I0(n43712), .I1(n38653), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n38654));
    defparam i31808_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(clk32MHz), 
           .D(n18073));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i31815_3_lut (.I0(n5_c), .I1(n6_adj_4261), .I2(n40522), .I3(GND_net), 
            .O(n38661));
    defparam i31815_3_lut.LUT_INIT = 16'hacac;
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(clk32MHz), 
           .D(n18072));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i31817_4_lut (.I0(n38661), .I1(n38654), .I2(\byte_transmit_counter[4] ), 
            .I3(\byte_transmit_counter[3] ), .O(n38663));
    defparam i31817_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31816_3_lut (.I0(n43772), .I1(n43766), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n38662));
    defparam i31816_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(clk32MHz), 
           .D(n17937));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(clk32MHz), 
           .D(n17936));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(clk32MHz), 
           .D(n17935));   // verilog/coms.v(127[12] 295[6])
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(clk32MHz), .D(n17934));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSR tx_transmit_3494 (.Q(r_SM_Main_2__N_3585[0]), .C(clk32MHz), 
            .D(n3332[0]), .R(n35671));   // verilog/coms.v(127[12] 295[6])
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3495  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(clk32MHz), .D(rx_data_ready));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(clk32MHz), 
           .D(n18071));   // verilog/coms.v(127[12] 295[6])
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(clk32MHz), .D(n17933));   // verilog/coms.v(127[12] 295[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(clk32MHz), .D(n17932));   // verilog/coms.v(127[12] 295[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(clk32MHz), .D(n17931));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(clk32MHz), 
           .D(n18070));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i3_4_lut_adj_998 (.I0(n30586), .I1(n35300), .I2(n30523), .I3(\data_in_frame[18] [0]), 
            .O(n15609));
    defparam i3_4_lut_adj_998.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_999 (.I0(\data_in_frame[20] [2]), .I1(\data_in_frame[22] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4262));
    defparam i1_2_lut_adj_999.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(clk32MHz), 
           .D(n18024));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i4_4_lut_adj_1000 (.I0(n36755), .I1(\data_in_frame[18] [1]), 
            .I2(n35300), .I3(n6_adj_4262), .O(n37377));
    defparam i4_4_lut_adj_1000.LUT_INIT = 16'h9669;
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(clk32MHz), .D(n17930));   // verilog/coms.v(127[12] 295[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(clk32MHz), .D(n17929));   // verilog/coms.v(127[12] 295[6])
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(clk32MHz), .D(n17928));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(clk32MHz), 
           .D(n17927));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(clk32MHz), 
           .D(n17926));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(clk32MHz), 
           .D(n17925));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(clk32MHz), 
           .D(n17924));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(clk32MHz), 
           .D(n17923));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(clk32MHz), 
           .D(n17922));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(clk32MHz), 
           .D(n17921));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(clk32MHz), 
           .D(n17920));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(clk32MHz), 
           .D(n17919));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(clk32MHz), 
           .D(n17918));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(clk32MHz), 
           .D(n17917));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(clk32MHz), 
           .D(n17916));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(clk32MHz), 
           .D(n17915));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 data_in_frame_9__7__I_0_3513_2_lut (.I0(\data_in_frame[9] [7]), 
            .I1(\data_in_frame[9] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_805));   // verilog/coms.v(70[16:27])
    defparam data_in_frame_9__7__I_0_3513_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(clk32MHz), 
           .D(n17914));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(clk32MHz), 
           .D(n17913));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut (.I0(\byte_transmit_counter[4] ), 
            .I1(\byte_transmit_counter[3] ), .I2(n38678), .I3(n38677), 
            .O(tx_data[5]));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(clk32MHz), 
           .D(n17912));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_adj_1001 (.I0(\data_in_frame[7] [2]), .I1(\data_in_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n35558));
    defparam i1_2_lut_adj_1001.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1002 (.I0(\data_in_frame[6] [5]), .I1(n35590), 
            .I2(n16777), .I3(GND_net), .O(n35438));   // verilog/coms.v(84[17:63])
    defparam i2_3_lut_adj_1002.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(clk32MHz), 
           .D(n17911));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(clk32MHz), 
           .D(n17910));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i3_4_lut_adj_1003 (.I0(\data_in_frame[9] [5]), .I1(n35360), 
            .I2(n16386), .I3(\data_in_frame[11] [6]), .O(n35543));
    defparam i3_4_lut_adj_1003.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(clk32MHz), 
           .D(n18040));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(clk32MHz), 
           .D(n18023));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14][1] ), .C(clk32MHz), 
           .D(n18047));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(clk32MHz), 
           .D(n18069));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(clk32MHz), 
           .D(n17909));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(clk32MHz), 
           .D(n18068));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(clk32MHz), 
           .D(n18046));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i28923_3_lut (.I0(n15886), .I1(n15963), .I2(\FRAME_MATCHER.state[3] ), 
            .I3(GND_net), .O(n35671));
    defparam i28923_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i8_4_lut (.I0(n35182), .I1(n35644), .I2(n16156), .I3(n35499), 
            .O(n20));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(n35413), .I1(n35110), .I2(n30671), .I3(n35581), 
            .O(n19_adj_4263));
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n35391), .I1(\data_in_frame[1] [1]), .I2(n35154), 
            .I3(n16044), .O(n21));
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut (.I0(n21), .I1(n19_adj_4263), .I2(n20), .I3(GND_net), 
            .O(n15568));
    defparam i11_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1004 (.I0(\data_in_frame[6] [0]), .I1(n35578), 
            .I2(\data_in_frame[8] [7]), .I3(GND_net), .O(n35327));
    defparam i2_3_lut_adj_1004.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1005 (.I0(\data_in_frame[7] [6]), .I1(\data_in_frame[8] [0]), 
            .I2(\data_in_frame[7] [7]), .I3(GND_net), .O(n35454));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1005.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut (.I0(\data_in_frame[7] [3]), .I1(\data_in_frame[7] [0]), 
            .I2(n35454), .I3(n35327), .O(n16));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1006 (.I0(n30578), .I1(n35438), .I2(n35629), 
            .I3(n35224), .O(n17));
    defparam i7_4_lut_adj_1006.LUT_INIT = 16'h6996;
    SB_LUT4 i13368_3_lut_4_lut (.I0(n8_adj_4260), .I1(n35006), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n18107));
    defparam i13368_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(clk32MHz), 
           .D(n18067));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(clk32MHz), 
           .D(n17908));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i3_4_lut_adj_1007 (.I0(n24966), .I1(n24738), .I2(n101), .I3(n5_adj_4264), 
            .O(n36982));
    defparam i3_4_lut_adj_1007.LUT_INIT = 16'hfffb;
    SB_LUT4 mux_788_i1_3_lut (.I0(n36982), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n4498), .I3(GND_net), .O(n3332[0]));   // verilog/coms.v(145[4] 294[11])
    defparam mux_788_i1_3_lut.LUT_INIT = 16'h5c5c;
    SB_LUT4 i9_4_lut_adj_1008 (.I0(n17), .I1(n16034), .I2(n16), .I3(\data_in_frame[8] [4]), 
            .O(n37006));
    defparam i9_4_lut_adj_1008.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1009 (.I0(n37597), .I1(\data_in_frame[13] [2]), 
            .I2(\data_in_frame[10] [7]), .I3(GND_net), .O(n35487));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1009.LUT_INIT = 16'h6969;
    SB_LUT4 i6_4_lut_adj_1010 (.I0(n16883), .I1(n12), .I2(n35487), .I3(\data_in_frame[13] [1]), 
            .O(n16272));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_1010.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1011 (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[17] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n35354));
    defparam i1_2_lut_adj_1011.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut (.I0(n31482), .I1(\data_in_frame[20] [1]), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13367_3_lut_4_lut (.I0(n8_adj_4260), .I1(n35006), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n18106));
    defparam i13367_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(153[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_adj_1012 (.I0(n16156), .I1(\data_in_frame[6] [4]), 
            .I2(\data_in_frame[6] [5]), .I3(GND_net), .O(n35227));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1012.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1013 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[8] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16034));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_adj_1013.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1014 (.I0(n16034), .I1(Kp_23__N_1186), .I2(n35227), 
            .I3(n37006), .O(n35518));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1014.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1015 (.I0(\data_in_frame[10] [7]), .I1(n37006), 
            .I2(GND_net), .I3(GND_net), .O(n35294));
    defparam i1_2_lut_adj_1015.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1016 (.I0(\data_in_frame[8] [2]), .I1(n35154), 
            .I2(\data_in_frame[6] [0]), .I3(\data_in_frame[6] [1]), .O(n16642));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_1016.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1017 (.I0(\data_in_frame[10] [4]), .I1(n16642), 
            .I2(GND_net), .I3(GND_net), .O(n35533));
    defparam i1_2_lut_adj_1017.LUT_INIT = 16'h6666;
    SB_LUT4 i13366_3_lut_4_lut (.I0(n8_adj_4260), .I1(n35006), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n18105));
    defparam i13366_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(clk32MHz), 
           .D(n17907));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18] [2]), .C(clk32MHz), 
           .D(n17906));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_adj_1018 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35385));
    defparam i1_2_lut_adj_1018.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1019 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16142));   // verilog/coms.v(71[16:41])
    defparam i1_2_lut_adj_1019.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1020 (.I0(\data_in_frame[6] [2]), .I1(n35122), 
            .I2(n16552), .I3(GND_net), .O(n16645));   // verilog/coms.v(72[16:42])
    defparam i2_3_lut_adj_1020.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1021 (.I0(n16464), .I1(n35224), .I2(n16782), 
            .I3(GND_net), .O(n16231));   // verilog/coms.v(71[16:41])
    defparam i2_3_lut_adj_1021.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1022 (.I0(n16231), .I1(n16645), .I2(GND_net), 
            .I3(GND_net), .O(n35167));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1022.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1023 (.I0(\data_in_frame[8] [5]), .I1(Kp_23__N_1186), 
            .I2(GND_net), .I3(GND_net), .O(n35617));
    defparam i1_2_lut_adj_1023.LUT_INIT = 16'h6666;
    SB_LUT4 i5_3_lut (.I0(n30529), .I1(n35617), .I2(n35135), .I3(GND_net), 
            .O(n14));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1024 (.I0(n35385), .I1(n35555), .I2(\data_in_frame[15] [2]), 
            .I3(n16645), .O(n15));
    defparam i6_4_lut_adj_1024.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1025 (.I0(n15), .I1(\data_in_frame[12] [6]), .I2(n14), 
            .I3(\data_in_frame[11] [0]), .O(n37527));
    defparam i8_4_lut_adj_1025.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1026 (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[17] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16835));
    defparam i1_2_lut_adj_1026.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1027 (.I0(\data_in_frame[21] [5]), .I1(\data_in_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n11));
    defparam i1_2_lut_adj_1027.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1028 (.I0(\data_in_frame[24] [4]), .I1(n37377), 
            .I2(n15609), .I3(\data_in_frame[22] [2]), .O(n36431));
    defparam i3_4_lut_adj_1028.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1029 (.I0(n31528), .I1(n30677), .I2(\data_in_frame[22] [6]), 
            .I3(n35347), .O(n10));
    defparam i4_4_lut_adj_1029.LUT_INIT = 16'h9669;
    SB_LUT4 i3_3_lut (.I0(\data_in_frame[23] [1]), .I1(n35276), .I2(n35508), 
            .I3(GND_net), .O(n8_adj_4265));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_adj_1030 (.I0(\data_in_frame[20] [4]), .I1(n10), .I2(\data_in_frame[24] [7]), 
            .I3(GND_net), .O(n37028));
    defparam i5_3_lut_adj_1030.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18] [1]), .C(clk32MHz), 
           .D(n17905));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 add_3597_9_lut (.I0(n34978), .I1(\byte_transmit_counter[7] ), 
            .I2(GND_net), .I3(n27926), .O(n40740)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3597_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3597_8_lut (.I0(\FRAME_MATCHER.i_31__N_2624 ), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n27925), .O(n40622)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3597_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3597_8 (.CI(n27925), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n27926));
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(clk32MHz), 
           .D(n18045));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(clk32MHz), 
           .D(n18044));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18] [0]), .C(clk32MHz), 
           .D(n17904));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i6_4_lut_adj_1031 (.I0(n35543), .I1(\data_in_frame[9] [4]), 
            .I2(\data_in_frame[12] [0]), .I3(n30671), .O(n14_adj_4266));
    defparam i6_4_lut_adj_1031.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(clk32MHz), 
           .D(n18043));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 add_3597_7_lut (.I0(n34978), .I1(\byte_transmit_counter[5] ), 
            .I2(GND_net), .I3(n27924), .O(n40742)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3597_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3597_7 (.CI(n27924), .I0(\byte_transmit_counter[5] ), .I1(GND_net), 
            .CO(n27925));
    SB_LUT4 add_3597_6_lut (.I0(n34978), .I1(\byte_transmit_counter[4] ), 
            .I2(GND_net), .I3(n27923), .O(n40743)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3597_6_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(clk32MHz), 
           .D(n18042));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(clk32MHz), 
           .D(n17903));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i31_3_lut_4_lut (.I0(\byte_transmit_counter[4] ), 
            .I1(\byte_transmit_counter[3] ), .I2(n38675), .I3(n38674), 
            .O(tx_data[4]));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i13370_3_lut_4_lut (.I0(n8_adj_4260), .I1(n35006), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n18109));
    defparam i13370_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(clk32MHz), 
           .D(n17902));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13369_3_lut_4_lut (.I0(n8_adj_4260), .I1(n35006), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n18108));
    defparam i13369_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_3597_6 (.CI(n27923), .I0(\byte_transmit_counter[4] ), .I1(GND_net), 
            .CO(n27924));
    SB_LUT4 add_3597_5_lut (.I0(\FRAME_MATCHER.i_31__N_2624 ), .I1(\byte_transmit_counter[3] ), 
            .I2(GND_net), .I3(n27922), .O(n40744)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3597_5_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i7_4_lut_adj_1032 (.I0(\data_in_frame[14] [2]), .I1(n14_adj_4266), 
            .I2(n10_adj_4267), .I3(\data_in_frame[12] [1]), .O(n36306));
    defparam i7_4_lut_adj_1032.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1033 (.I0(n37132), .I1(\data_in_frame[16] [3]), 
            .I2(n36306), .I3(GND_net), .O(n31558));
    defparam i2_3_lut_adj_1033.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1034 (.I0(n30683), .I1(\data_in_frame[15] [7]), 
            .I2(n30689), .I3(GND_net), .O(n35147));
    defparam i2_3_lut_adj_1034.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1035 (.I0(\data_in_frame[9] [4]), .I1(\data_in_frame[9] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16086));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1035.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1036 (.I0(\data_in_frame[7] [3]), .I1(\data_in_frame[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35394));
    defparam i1_2_lut_adj_1036.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1037 (.I0(\data_in_frame[9] [5]), .I1(n17011), 
            .I2(n35394), .I3(n30671), .O(n35370));
    defparam i3_4_lut_adj_1037.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut (.I0(n35144), .I1(n35370), .I2(\data_in_frame[14] [0]), 
            .I3(n31571), .O(n12_adj_4268));
    defparam i5_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1038 (.I0(\data_in_frame[11] [6]), .I1(n12_adj_4268), 
            .I2(n35552), .I3(\data_in_frame[13] [7]), .O(n30592));
    defparam i6_4_lut_adj_1038.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1039 (.I0(\data_in_frame[13] [7]), .I1(\data_in_frame[12] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35463));
    defparam i1_2_lut_adj_1039.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1040 (.I0(\data_in_frame[11] [5]), .I1(\data_in_frame[11] [7]), 
            .I2(\data_in_frame[7] [5]), .I3(GND_net), .O(n35626));
    defparam i2_3_lut_adj_1040.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1041 (.I0(n30592), .I1(\data_in_frame[16] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35367));
    defparam i1_2_lut_adj_1041.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1042 (.I0(n30592), .I1(n35147), .I2(\data_in_frame[16] [1]), 
            .I3(GND_net), .O(n30807));   // verilog/coms.v(84[17:70])
    defparam i2_3_lut_adj_1042.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1043 (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[18] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n35341));
    defparam i1_2_lut_adj_1043.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1044 (.I0(\data_in_frame[20] [3]), .I1(\data_in_frame[20] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n16202));
    defparam i1_2_lut_adj_1044.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1045 (.I0(n35493), .I1(Kp_23__N_1802), .I2(\data_in_frame[23] [0]), 
            .I3(n35602), .O(n10_adj_4269));
    defparam i4_4_lut_adj_1045.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1046 (.I0(n35546), .I1(\data_in_frame[18] [7]), 
            .I2(\data_in_frame[23] [2]), .I3(n35364), .O(n15_adj_4270));
    defparam i6_4_lut_adj_1046.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1047 (.I0(n35273), .I1(\data_in_frame[19] [3]), 
            .I2(n35218), .I3(n30586), .O(n21_adj_4271));
    defparam i8_4_lut_adj_1047.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut (.I0(n30812), .I1(\data_in_frame[21] [6]), .I2(n35599), 
            .I3(GND_net), .O(n20_adj_4272));
    defparam i7_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut_adj_1048 (.I0(n21_adj_4271), .I1(n35493), .I2(n18), 
            .I3(n35157), .O(n24));
    defparam i11_4_lut_adj_1048.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut (.I0(\data_in_frame[24] [3]), .I1(n35176), .I2(\data_in_frame[22] [2]), 
            .I3(\data_in_frame[22] [1]), .O(n37548));
    defparam i2_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1049 (.I0(\data_in_frame[16] [7]), .I1(n11), .I2(n31470), 
            .I3(n12_adj_4273), .O(n18_adj_4274));
    defparam i8_4_lut_adj_1049.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1050 (.I0(n35511), .I1(\data_in_frame[23] [4]), 
            .I2(n35037), .I3(n30721), .O(n14_adj_4275));
    defparam i6_4_lut_adj_1050.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1051 (.I0(n35515), .I1(n35364), .I2(n35259), 
            .I3(\data_in_frame[21] [4]), .O(n17_adj_4276));
    defparam i7_4_lut_adj_1051.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1052 (.I0(\data_in_frame[21] [2]), .I1(n35410), 
            .I2(\data_in_frame[19] [2]), .I3(\data_in_frame[21] [3]), .O(n13));
    defparam i5_4_lut_adj_1052.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1053 (.I0(\data_in_frame[21] [1]), .I1(\data_in_frame[19] [1]), 
            .I2(\data_in_frame[21] [2]), .I3(GND_net), .O(n9));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1053.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1054 (.I0(n17023), .I1(\data_in_frame[18] [7]), 
            .I2(n35276), .I3(\data_in_frame[17] [0]), .O(n11_adj_4277));   // verilog/coms.v(75[16:43])
    defparam i4_4_lut_adj_1054.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1055 (.I0(\data_in_frame[21] [4]), .I1(n31460), 
            .I2(\data_in_frame[21] [3]), .I3(n35407), .O(n8_adj_4278));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_1055.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1056 (.I0(n11_adj_4277), .I1(n9), .I2(\data_in_frame[23] [3]), 
            .I3(n16838), .O(n36572));   // verilog/coms.v(75[16:43])
    defparam i6_4_lut_adj_1056.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1057 (.I0(n36431), .I1(n30677), .I2(n35344), 
            .I3(\data_in_frame[24] [6]), .O(n24_adj_4279));
    defparam i8_4_lut_adj_1057.LUT_INIT = 16'hebbe;
    SB_LUT4 i6_4_lut_adj_1058 (.I0(\data_in_frame[22] [7]), .I1(n37028), 
            .I2(n8_adj_4265), .I3(n35347), .O(n22));
    defparam i6_4_lut_adj_1058.LUT_INIT = 16'hdeed;
    SB_LUT4 i31750_4_lut (.I0(\data_in_frame[24] [5]), .I1(n36394), .I2(n35344), 
            .I3(n37377), .O(n38515));
    defparam i31750_4_lut.LUT_INIT = 16'h4884;
    SB_LUT4 i5_4_lut_adj_1059 (.I0(\data_in_frame[24] [2]), .I1(n36572), 
            .I2(n35466), .I3(\data_in_frame[22] [1]), .O(n21_adj_4280));
    defparam i5_4_lut_adj_1059.LUT_INIT = 16'hb77b;
    SB_LUT4 i5_4_lut_adj_1060 (.I0(n35279), .I1(n10_adj_4269), .I2(\data_in_frame[20] [7]), 
            .I3(n31474), .O(n36878));
    defparam i5_4_lut_adj_1060.LUT_INIT = 16'h9669;
    SB_LUT4 i8_4_lut_adj_1061 (.I0(n15_adj_4270), .I1(n37403), .I2(n14_adj_4281), 
            .I3(\data_in_frame[21] [1]), .O(n36317));
    defparam i8_4_lut_adj_1061.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut_adj_1062 (.I0(\data_in_frame[23] [7]), .I1(n24), .I2(n20_adj_4272), 
            .I3(\data_in_frame[20] [5]), .O(n37411));
    defparam i12_4_lut_adj_1062.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(clk32MHz), 
           .D(n17901));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(clk32MHz), 
           .D(n17900));   // verilog/coms.v(127[12] 295[6])
    SB_CARRY add_3597_5 (.CI(n27922), .I0(\byte_transmit_counter[3] ), .I1(GND_net), 
            .CO(n27923));
    SB_LUT4 add_3597_4_lut (.I0(\FRAME_MATCHER.i_31__N_2624 ), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(n27921), .O(n40747)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3597_4_lut.LUT_INIT = 16'h8228;
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(clk32MHz), 
           .D(n17899));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i3_4_lut_adj_1063 (.I0(n37080), .I1(n35466), .I2(n15609), 
            .I3(\data_in_frame[24] [0]), .O(n37572));
    defparam i3_4_lut_adj_1063.LUT_INIT = 16'h9669;
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(clk32MHz), 
           .D(n18041));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(clk32MHz), 
           .D(n17898));   // verilog/coms.v(127[12] 295[6])
    SB_CARRY add_3597_4 (.CI(n27921), .I0(\byte_transmit_counter[2] ), .I1(GND_net), 
            .CO(n27922));
    SB_LUT4 i13365_3_lut_4_lut (.I0(n8_adj_4260), .I1(n35006), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n18104));
    defparam i13365_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(clk32MHz), 
           .D(n17897));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(clk32MHz), 
           .D(n17896));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(clk32MHz), 
           .D(n17895));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(clk32MHz), 
           .D(n17894));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i4_4_lut_adj_1064 (.I0(n37548), .I1(n37080), .I2(n35176), 
            .I3(\data_in_frame[24] [1]), .O(n20_adj_4282));
    defparam i4_4_lut_adj_1064.LUT_INIT = 16'hbeeb;
    SB_LUT4 i3_4_lut_adj_1065 (.I0(n13), .I1(n17_adj_4276), .I2(n14_adj_4275), 
            .I3(n18_adj_4274), .O(n19_adj_4283));
    defparam i3_4_lut_adj_1065.LUT_INIT = 16'hb7ed;
    SB_LUT4 i14_4_lut (.I0(n21_adj_4280), .I1(n38515), .I2(n22), .I3(n24_adj_4279), 
            .O(n30_adj_4284));
    defparam i14_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i9_4_lut_adj_1066 (.I0(n37572), .I1(n37411), .I2(n36317), 
            .I3(n36878), .O(n25));
    defparam i9_4_lut_adj_1066.LUT_INIT = 16'hffef;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n30_adj_4284), .I2(n19_adj_4283), 
            .I3(n20_adj_4282), .O(n31));
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i13364_3_lut_4_lut (.I0(n8_adj_4260), .I1(n35006), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n18103));
    defparam i13364_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13363_3_lut_4_lut (.I0(n8_adj_4260), .I1(n35006), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n18102));
    defparam i13363_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1067 (.I0(n13414), .I1(n31), .I2(n31_adj_4285), 
            .I3(\FRAME_MATCHER.state[1] ), .O(n26));   // verilog/coms.v(111[11:16])
    defparam i1_4_lut_adj_1067.LUT_INIT = 16'hfaee;
    SB_LUT4 i3_4_lut_adj_1068 (.I0(\data_in_frame[0] [6]), .I1(n35101), 
            .I2(n35051), .I3(n16494), .O(n15531));   // verilog/coms.v(77[16:27])
    defparam i3_4_lut_adj_1068.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1069 (.I0(\data_in_frame[4] [0]), .I1(n35170), 
            .I2(\data_in_frame[3] [6]), .I3(\data_in_frame[3] [7]), .O(n16552));   // verilog/coms.v(72[16:42])
    defparam i3_4_lut_adj_1069.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1070 (.I0(\data_in_frame[5] [3]), .I1(n15531), 
            .I2(GND_net), .I3(GND_net), .O(n16399));
    defparam i1_2_lut_adj_1070.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1071 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[2] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35051));   // verilog/coms.v(69[16:69])
    defparam i1_2_lut_adj_1071.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(clk32MHz), 
           .D(n17893));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(clk32MHz), 
           .D(n17892));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(clk32MHz), 
           .D(n17891));   // verilog/coms.v(127[12] 295[6])
    SB_DFFESR driver_enable_3498 (.Q(PIN_11_c), .C(clk32MHz), .E(n35783), 
            .D(n4462), .R(n37191));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(clk32MHz), 
           .D(n17890));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(clk32MHz), 
           .D(n17889));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(clk32MHz), 
           .D(n17888));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(clk32MHz), 
           .D(n17887));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(clk32MHz), 
           .D(n17886));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(clk32MHz), 
           .D(n17885));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(clk32MHz), 
           .D(n17884));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(clk32MHz), 
           .D(n17883));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(clk32MHz), 
           .D(n17882));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(clk32MHz), 
           .D(n17881));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(clk32MHz), 
           .D(n17880));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13235_3_lut_4_lut (.I0(n8_adj_4260), .I1(n34998), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n17974));
    defparam i13235_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(clk32MHz), 
           .D(n17879));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(clk32MHz), 
           .D(n17878));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(clk32MHz), 
           .D(n17877));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(clk32MHz), 
           .D(n17876));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(clk32MHz), 
           .D(n17875));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(clk32MHz), 
           .D(n17874));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(clk32MHz), 
           .D(n17873));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i3_4_lut_adj_1072 (.I0(\data_in_frame[5] [1]), .I1(\data_in_frame[1] [0]), 
            .I2(n35416), .I3(n35051), .O(n30671));   // verilog/coms.v(69[16:69])
    defparam i3_4_lut_adj_1072.LUT_INIT = 16'h6996;
    SB_LUT4 add_3597_3_lut (.I0(\FRAME_MATCHER.i_31__N_2624 ), .I1(\byte_transmit_counter[1] ), 
            .I2(GND_net), .I3(n27920), .O(n40746)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3597_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3597_3 (.CI(n27920), .I0(\byte_transmit_counter[1] ), .I1(GND_net), 
            .CO(n27921));
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(clk32MHz), 
           .D(n17872));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(clk32MHz), 
           .D(n17871));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(clk32MHz), 
           .D(n17870));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(clk32MHz), 
           .D(n17869));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(clk32MHz), 
           .D(n17868));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(clk32MHz), 
           .D(n17867));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(clk32MHz), 
           .D(n17866));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(clk32MHz), 
           .D(n17865));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(clk32MHz), 
           .D(n17864));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(clk32MHz), 
           .D(n17863));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(clk32MHz), 
           .D(n17862));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(clk32MHz), 
           .D(n17861));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(clk32MHz), 
           .D(n17860));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13236_3_lut_4_lut (.I0(n8_adj_4260), .I1(n34998), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n17975));
    defparam i13236_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(clk32MHz), 
           .D(n17859));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(clk32MHz), 
           .D(n17858));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(clk32MHz), 
           .D(n17857));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(clk32MHz), 
           .D(n17856));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(clk32MHz), 
           .D(n17855));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(clk32MHz), 
           .D(n17854));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(clk32MHz), 
           .D(n17853));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(clk32MHz), 
           .D(n17852));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_adj_1073 (.I0(\data_in_frame[20] [5]), .I1(n36436), 
            .I2(GND_net), .I3(GND_net), .O(n35347));
    defparam i1_2_lut_adj_1073.LUT_INIT = 16'h9999;
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(clk32MHz), 
           .D(n17851));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(clk32MHz), 
           .D(n17850));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(clk32MHz), 
           .D(n17849));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(clk32MHz), 
           .D(n17848));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(clk32MHz), 
           .D(n17847));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(clk32MHz), 
           .D(n17846));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(clk32MHz), 
           .D(n17845));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i36773_3_lut (.I0(\FRAME_MATCHER.state[3] ), .I1(n35671), .I2(n15886), 
            .I3(GND_net), .O(n37191));
    defparam i36773_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i36776_4_lut (.I0(n35671), .I1(\FRAME_MATCHER.state[3] ), .I2(n4462), 
            .I3(n4498), .O(n35783));
    defparam i36776_4_lut.LUT_INIT = 16'h5011;
    SB_LUT4 add_3597_2_lut (.I0(\FRAME_MATCHER.i_31__N_2624 ), .I1(\byte_transmit_counter[0] ), 
            .I2(tx_transmit_N_3482), .I3(GND_net), .O(n40745)) /* synthesis syn_instantiated=1 */ ;
    defparam add_3597_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i36056_2_lut (.I0(\FRAME_MATCHER.state[1] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(GND_net), .I3(GND_net), .O(n4462));   // verilog/coms.v(145[4] 294[11])
    defparam i36056_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i13237_3_lut_4_lut (.I0(n8_adj_4260), .I1(n34998), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n17976));
    defparam i13237_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(clk32MHz), 
           .D(n17844));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i2_3_lut_adj_1074 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[3] [7]), .I3(GND_net), .O(n35182));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_adj_1074.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1075 (.I0(\data_in_frame[4] [4]), .I1(n35104), 
            .I2(GND_net), .I3(GND_net), .O(n16953));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1075.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1076 (.I0(\data_in_frame[1] [7]), .I1(n35182), 
            .I2(\data_in_frame[1] [5]), .I3(GND_net), .O(n16782));   // verilog/coms.v(69[16:27])
    defparam i2_3_lut_adj_1076.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1077 (.I0(\data_in_frame[1] [7]), .I1(n35413), 
            .I2(GND_net), .I3(GND_net), .O(n16555));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1077.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1078 (.I0(\data_in_frame[3] [3]), .I1(\data_in_frame[5] [4]), 
            .I2(\data_in_frame[1] [2]), .I3(n6_adj_4286), .O(n16386));   // verilog/coms.v(72[16:34])
    defparam i4_4_lut_adj_1078.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1079 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[0] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4287));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1079.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1080 (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[2] [1]), 
            .I2(\data_in_frame[1] [6]), .I3(n6_adj_4287), .O(n17042));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1080.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1081 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n16038));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_adj_1081.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1082 (.I0(\data_in_frame[2] [4]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n5_adj_4288));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_adj_1082.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1083 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35048));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1083.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(clk32MHz), 
           .D(n17843));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(clk32MHz), 
           .D(n17842));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(clk32MHz), 
           .D(n17841));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(clk32MHz), 
           .D(n17840));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(clk32MHz), 
           .D(n17839));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_adj_1084 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[2] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35044));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1084.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(clk32MHz), 
           .D(n17838));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_adj_1085 (.I0(\data_in_frame[3] [2]), .I1(\data_in_frame[3] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16494));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_adj_1085.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(clk32MHz), 
           .D(n17837));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_adj_1086 (.I0(n5_adj_4288), .I1(n6_adj_4289), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1003));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1086.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1087 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n35138));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1087.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(clk32MHz), 
           .D(n17836));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_adj_1088 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35170));   // verilog/coms.v(72[16:42])
    defparam i1_2_lut_adj_1088.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(clk32MHz), 
           .D(n17835));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i4_4_lut_adj_1089 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [0]), 
            .I2(n8_adj_4290), .I3(\data_in_frame[1] [1]), .O(n18_adj_4291));   // verilog/coms.v(77[16:27])
    defparam i4_4_lut_adj_1089.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1090 (.I0(\data_in_frame[2] [1]), .I1(n35138), 
            .I2(\data_in_frame[0] [6]), .I3(\data_in_frame[0] [7]), .O(n24_adj_4292));   // verilog/coms.v(77[16:27])
    defparam i10_4_lut_adj_1090.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(clk32MHz), 
           .D(n17834));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i8_4_lut_adj_1091 (.I0(Kp_23__N_1003), .I1(\data_in_frame[2] [0]), 
            .I2(n16494), .I3(n35104), .O(n22_adj_4293));   // verilog/coms.v(77[16:27])
    defparam i8_4_lut_adj_1091.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1092 (.I0(\data_in_frame[2] [7]), .I1(n24_adj_4292), 
            .I2(n18_adj_4291), .I3(n35268), .O(n26_adj_4294));   // verilog/coms.v(77[16:27])
    defparam i12_4_lut_adj_1092.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(clk32MHz), 
           .D(n17833));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13_4_lut_adj_1093 (.I0(n35048), .I1(n26_adj_4294), .I2(n22_adj_4293), 
            .I3(\data_in_frame[0] [5]), .O(n37530));   // verilog/coms.v(77[16:27])
    defparam i13_4_lut_adj_1093.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1094 (.I0(n16038), .I1(n37530), .I2(n35441), 
            .I3(\data_in_frame[3] [7]), .O(n35098));   // verilog/coms.v(69[16:27])
    defparam i3_4_lut_adj_1094.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(clk32MHz), 
           .D(n17832));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_adj_1095 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n16044));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1095.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(clk32MHz), 
           .D(n17831));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_adj_1096 (.I0(\data_in_frame[3] [3]), .I1(\data_in_frame[3] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35441));   // verilog/coms.v(72[16:34])
    defparam i1_2_lut_adj_1096.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(clk32MHz), 
           .D(n17830));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(clk32MHz), 
           .D(n17829));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_adj_1097 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n35101));   // verilog/coms.v(72[16:34])
    defparam i1_2_lut_adj_1097.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(clk32MHz), 
           .D(n17828));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_adj_1098 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[2] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35268));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_1098.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(clk32MHz), 
           .D(n17827));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(clk32MHz), 
           .D(n17826));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i2_3_lut_adj_1099 (.I0(\data_in_frame[5] [2]), .I1(n35245), 
            .I2(\data_in_frame[3] [1]), .I3(GND_net), .O(n35499));
    defparam i2_3_lut_adj_1099.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(clk32MHz), 
           .D(n17825));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(clk32MHz), 
           .D(n17824));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(clk32MHz), 
           .D(n17823));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(clk32MHz), 
           .D(n17822));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i3_4_lut_adj_1100 (.I0(\data_in_frame[5] [0]), .I1(n16044), 
            .I2(n35416), .I3(n35245), .O(n30669));
    defparam i3_4_lut_adj_1100.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(clk32MHz), 
           .D(n17821));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i2_2_lut_adj_1101 (.I0(n35098), .I1(\data_in_frame[3] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4295));   // verilog/coms.v(69[16:27])
    defparam i2_2_lut_adj_1101.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(clk32MHz), 
           .D(n17820));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_4_lut_adj_1102 (.I0(\data_in_frame[4] [7]), .I1(n6_adj_4289), 
            .I2(n6_adj_4295), .I3(\data_in_frame[1] [5]), .O(n17011));
    defparam i1_4_lut_adj_1102.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(clk32MHz), 
           .D(n17819));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i3_4_lut_adj_1103 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[3] [4]), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[3] [5]), .O(Kp_23__N_949));   // verilog/coms.v(75[16:43])
    defparam i3_4_lut_adj_1103.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(clk32MHz), 
           .D(n17818));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_adj_1104 (.I0(\data_in_frame[5] [6]), .I1(Kp_23__N_949), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4296));
    defparam i1_2_lut_adj_1104.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(clk32MHz), 
           .D(n17817));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i2_3_lut_adj_1105 (.I0(\data_in_frame[1] [5]), .I1(n35110), 
            .I2(\data_in_frame[1] [3]), .I3(GND_net), .O(n16464));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_adj_1105.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(clk32MHz), 
           .D(n17816));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i6_4_lut_adj_1106 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[0] [4]), .I3(\data_in_frame[0] [0]), .O(n14_adj_4297));
    defparam i6_4_lut_adj_1106.LUT_INIT = 16'hfbff;
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(clk32MHz), 
           .D(n17815));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_adj_1107 (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4298));
    defparam i1_2_lut_adj_1107.LUT_INIT = 16'heeee;
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(clk32MHz), 
           .D(n17814));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i7_4_lut_adj_1108 (.I0(n9_adj_4298), .I1(n14_adj_4297), .I2(\data_in_frame[0] [5]), 
            .I3(\data_in_frame[0] [2]), .O(n13414));
    defparam i7_4_lut_adj_1108.LUT_INIT = 16'hfeff;
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(clk32MHz), 
           .D(n17813));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i3_4_lut_adj_1109 (.I0(n17011), .I1(n30669), .I2(n16360), 
            .I3(n16115), .O(n37247));   // verilog/coms.v(231[9:81])
    defparam i3_4_lut_adj_1109.LUT_INIT = 16'hefff;
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(clk32MHz), 
           .D(n17812));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i3_2_lut (.I0(n16876), .I1(n17042), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4299));   // verilog/coms.v(231[9:81])
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(clk32MHz), 
           .D(n17811));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i9_4_lut_adj_1110 (.I0(n16386), .I1(n16555), .I2(n16782), 
            .I3(n16953), .O(n22_adj_4300));   // verilog/coms.v(231[9:81])
    defparam i9_4_lut_adj_1110.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(clk32MHz), 
           .D(n17810));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i7_3_lut_adj_1111 (.I0(n30671), .I1(n37247), .I2(n16777), 
            .I3(GND_net), .O(n20_adj_4301));   // verilog/coms.v(231[9:81])
    defparam i7_3_lut_adj_1111.LUT_INIT = 16'hfefe;
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(clk32MHz), 
           .D(n17809));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i11_4_lut_adj_1112 (.I0(n16464), .I1(n22_adj_4300), .I2(n16_adj_4299), 
            .I3(n6_adj_4296), .O(n24_adj_4302));   // verilog/coms.v(231[9:81])
    defparam i11_4_lut_adj_1112.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(clk32MHz), 
           .D(n17808));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i12_4_lut_adj_1113 (.I0(n16399), .I1(n24_adj_4302), .I2(n20_adj_4301), 
            .I3(n16552), .O(n31_adj_4285));   // verilog/coms.v(231[9:81])
    defparam i12_4_lut_adj_1113.LUT_INIT = 16'hfffe;
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(clk32MHz), 
           .D(n17807));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i2_3_lut_adj_1114 (.I0(n31_adj_4285), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(n13414), .I3(GND_net), .O(n4385));
    defparam i2_3_lut_adj_1114.LUT_INIT = 16'h0404;
    SB_LUT4 i5_4_lut_adj_1115 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n24968), .I3(n24910), .O(n12_adj_4303));
    defparam i5_4_lut_adj_1115.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1116 (.I0(\FRAME_MATCHER.state [2]), .I1(n12_adj_4303), 
            .I2(n26), .I3(n24686), .O(n37622));
    defparam i6_4_lut_adj_1116.LUT_INIT = 16'hfffd;
    SB_LUT4 mux_1080_i23_3_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n4385), .I3(GND_net), .O(n4408));
    defparam mux_1080_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(clk32MHz), 
           .D(n17806));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(clk32MHz), 
           .D(n17805));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(clk32MHz), 
           .D(n17804));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i4_4_lut_adj_1117 (.I0(n35341), .I1(n36755), .I2(n35536), 
            .I3(n6_adj_4304), .O(n30677));
    defparam i4_4_lut_adj_1117.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1118 (.I0(\data_in_frame[17] [4]), .I1(n16272), 
            .I2(GND_net), .I3(GND_net), .O(n35173));
    defparam i1_2_lut_adj_1118.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1119 (.I0(n30669), .I1(\data_in_frame[7] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35360));
    defparam i1_2_lut_adj_1119.LUT_INIT = 16'h9999;
    SB_LUT4 i6_4_lut_adj_1120 (.I0(n16360), .I1(\data_in_frame[7] [3]), 
            .I2(n16876), .I3(\data_in_frame[11] [4]), .O(n14_adj_4305));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_1120.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(clk32MHz), 
           .D(n17803));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(clk32MHz), 
           .D(n17802));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(clk32MHz), 
           .D(n17801));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(clk32MHz), 
           .D(n17800));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(clk32MHz), .D(n17799));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(clk32MHz), .D(n17798));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(clk32MHz), .D(n17797));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(clk32MHz), .D(n17796));   // verilog/coms.v(127[12] 295[6])
    SB_CARRY add_3597_2 (.CI(GND_net), .I0(\byte_transmit_counter[0] ), 
            .I1(tx_transmit_N_3482), .CO(n27920));
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(clk32MHz), .D(n17795));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(clk32MHz), .D(n17794));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(clk32MHz), .D(n17793));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(clk32MHz), .D(n17792));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(clk32MHz), .D(n17791));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(clk32MHz), .D(n17790));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(clk32MHz), .D(n17789));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(clk32MHz), .D(n17788));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(clk32MHz), .D(n17787));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(clk32MHz), .D(n17786));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(clk32MHz), .D(n17785));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(clk32MHz), .D(n17784));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(clk32MHz), .D(n17783));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(clk32MHz), .D(n17782));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(clk32MHz), .D(n17781));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(clk32MHz), .D(n17780));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(clk32MHz), .D(n17779));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13238_3_lut_4_lut (.I0(n8_adj_4260), .I1(n34998), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n17977));
    defparam i13238_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13239_3_lut_4_lut (.I0(n8_adj_4260), .I1(n34998), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n17978));
    defparam i13239_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(clk32MHz), .D(n17778));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(clk32MHz), .D(n17777));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(clk32MHz), .D(n17776));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13240_3_lut_4_lut (.I0(n8_adj_4260), .I1(n34998), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n17979));
    defparam i13240_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(clk32MHz), .D(n17775));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(clk32MHz), .D(n17774));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13241_3_lut_4_lut (.I0(n8_adj_4260), .I1(n34998), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n17980));
    defparam i13241_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(clk32MHz), .D(n17773));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13242_3_lut_4_lut (.I0(n8_adj_4260), .I1(n34998), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n17981));
    defparam i13242_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(clk32MHz), .D(n17772));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(clk32MHz), .D(n17771));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(clk32MHz), .D(n17770));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(clk32MHz), .D(n17769));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(clk32MHz), .D(n17768));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(clk32MHz), .D(n17767));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(clk32MHz), .D(n17766));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(clk32MHz), .D(n17765));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(clk32MHz), .D(n17764));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(clk32MHz), .D(n17763));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(clk32MHz), .D(n17762));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_3_lut (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(n30584), .I3(GND_net), .O(n31464));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(clk32MHz), .D(n17761));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(clk32MHz), .D(n17760));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(clk32MHz), .D(n17759));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(clk32MHz), .D(n17758));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(clk32MHz), .D(n17757));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(clk32MHz), .D(n17756));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(clk32MHz), .D(n17755));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(clk32MHz), .D(n17754));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(clk32MHz), .D(n17753));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(clk32MHz), .D(n17752));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(clk32MHz), .D(n17751));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(clk32MHz), .D(n17750));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(clk32MHz), .D(n17749));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(clk32MHz), .D(n17748));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(clk32MHz), .D(n17747));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(clk32MHz), .D(n17746));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(clk32MHz), .D(n17745));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i2_3_lut_4_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[8] [2]), .I3(\data_out_frame[6] [1]), .O(n16345));   // verilog/coms.v(84[17:28])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1121 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[8] [0]), .I3(GND_net), .O(n4_c));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_3_lut_adj_1121.LUT_INIT = 16'h9696;
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(clk32MHz), .D(n17744));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(clk32MHz), .D(n17743));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(clk32MHz), .D(n17742));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(clk32MHz), .D(n17741));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(clk32MHz), .D(n17740));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1122 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[7] [3]), 
            .I2(n36548), .I3(n16029), .O(n35426));
    defparam i2_3_lut_4_lut_adj_1122.LUT_INIT = 16'h6996;
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(clk32MHz), .D(n17739));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i23 (.Q(gearBoxRatio[23]), .C(clk32MHz), .D(n17738));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i22 (.Q(gearBoxRatio[22]), .C(clk32MHz), .D(n17737));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i21 (.Q(gearBoxRatio[21]), .C(clk32MHz), .D(n17736));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i14_3_lut_4_lut (.I0(\data_out_frame[9] [4]), .I1(n35256), .I2(n28_adj_4306), 
            .I3(\data_out_frame[10] [0]), .O(n32));   // verilog/coms.v(84[17:63])
    defparam i14_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF gearBoxRatio_i0_i20 (.Q(gearBoxRatio[20]), .C(clk32MHz), .D(n17735));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i19 (.Q(gearBoxRatio[19]), .C(clk32MHz), .D(n17734));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i18 (.Q(gearBoxRatio[18]), .C(clk32MHz), .D(n17733));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i17 (.Q(gearBoxRatio[17]), .C(clk32MHz), .D(n17732));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i16 (.Q(gearBoxRatio[16]), .C(clk32MHz), .D(n17731));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i15 (.Q(gearBoxRatio[15]), .C(clk32MHz), .D(n17730));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i14 (.Q(gearBoxRatio[14]), .C(clk32MHz), .D(n17729));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i13 (.Q(gearBoxRatio[13]), .C(clk32MHz), .D(n17728));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i12 (.Q(gearBoxRatio[12]), .C(clk32MHz), .D(n17727));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1123 (.I0(\data_out_frame[9] [4]), .I1(n35256), 
            .I2(n16006), .I3(\data_out_frame[9] [5]), .O(n35221));   // verilog/coms.v(84[17:63])
    defparam i2_3_lut_4_lut_adj_1123.LUT_INIT = 16'h6996;
    SB_DFF gearBoxRatio_i0_i11 (.Q(gearBoxRatio[11]), .C(clk32MHz), .D(n17726));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i10 (.Q(gearBoxRatio[10]), .C(clk32MHz), .D(n17725));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i9 (.Q(gearBoxRatio[9]), .C(clk32MHz), .D(n17724));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i8 (.Q(gearBoxRatio[8]), .C(clk32MHz), .D(n17723));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i7 (.Q(gearBoxRatio[7]), .C(clk32MHz), .D(n17722));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i6 (.Q(gearBoxRatio[6]), .C(clk32MHz), .D(n17721));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i5 (.Q(gearBoxRatio[5]), .C(clk32MHz), .D(n17720));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1124 (.I0(\data_in_frame[2] [3]), .I1(n35048), 
            .I2(\data_in_frame[4] [5]), .I3(n5_adj_4288), .O(n16777));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_4_lut_adj_1124.LUT_INIT = 16'h6996;
    SB_LUT4 i31797_4_lut (.I0(\data_in_frame[0] [3]), .I1(\data_in_frame[0] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(\data_in_frame[0] [7]), .O(n38569));
    defparam i31797_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1125 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4307));
    defparam i1_2_lut_adj_1125.LUT_INIT = 16'h8888;
    SB_LUT4 i7_4_lut_adj_1126 (.I0(n9_adj_4307), .I1(n38569), .I2(\data_in_frame[0] [6]), 
            .I3(\data_in_frame[0] [0]), .O(n34891));
    defparam i7_4_lut_adj_1126.LUT_INIT = 16'h0200;
    SB_LUT4 i2_3_lut_adj_1127 (.I0(n31), .I1(n34891), .I2(n15950), .I3(GND_net), 
            .O(n4593));
    defparam i2_3_lut_adj_1127.LUT_INIT = 16'h0404;
    SB_LUT4 i2_3_lut_4_lut_adj_1128 (.I0(\data_in_frame[2] [3]), .I1(n35048), 
            .I2(\data_in_frame[0] [0]), .I3(n35044), .O(n35104));   // verilog/coms.v(166[9:87])
    defparam i2_3_lut_4_lut_adj_1128.LUT_INIT = 16'h6996;
    SB_DFF gearBoxRatio_i0_i4 (.Q(gearBoxRatio[4]), .C(clk32MHz), .D(n17719));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i3 (.Q(gearBoxRatio[3]), .C(clk32MHz), .D(n17718));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1129 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[5] [7]), .I3(GND_net), .O(n6_adj_4308));
    defparam i1_2_lut_3_lut_adj_1129.LUT_INIT = 16'h9696;
    SB_DFF gearBoxRatio_i0_i2 (.Q(gearBoxRatio[2]), .C(clk32MHz), .D(n17717));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i4_4_lut_4_lut (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[8] [1]), 
            .I2(n4_adj_4309), .I3(n16445), .O(n30584));
    defparam i4_4_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF gearBoxRatio_i0_i1 (.Q(gearBoxRatio[1]), .C(clk32MHz), .D(n17716));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i5_3_lut_4_lut (.I0(n16345), .I1(n16716), .I2(n16239), .I3(n10_adj_4310), 
            .O(n35151));
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1080_i2_3_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n4385), .I3(GND_net), .O(n4387));
    defparam mux_1080_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1130 (.I0(n16345), .I1(n16716), .I2(\data_out_frame[10] [5]), 
            .I3(\data_out_frame[10] [4]), .O(n35584));
    defparam i2_3_lut_4_lut_adj_1130.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1080_i12_3_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n4385), .I3(GND_net), .O(n4397));
    defparam mux_1080_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1131 (.I0(\data_out_frame[18] [5]), .I1(n37560), 
            .I2(n36894), .I3(\data_out_frame[18] [4]), .O(n31480));
    defparam i2_3_lut_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1080_i11_3_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n4385), .I3(GND_net), .O(n4396));
    defparam mux_1080_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(clk32MHz), .D(n17714));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 mux_1080_i10_3_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n4385), .I3(GND_net), .O(n4395));
    defparam mux_1080_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(clk32MHz), .D(n17713));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(clk32MHz), .D(n17712));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(clk32MHz), .D(n17711));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(clk32MHz), .D(n17710));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(clk32MHz), .D(n17709));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(clk32MHz), .D(n17708));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(clk32MHz), .D(n17707));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(clk32MHz), .D(n17706));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(clk32MHz), .D(n17705));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(clk32MHz), .D(n17704));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(clk32MHz), .D(n17703));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(clk32MHz), .D(n17702));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(clk32MHz), .D(n17701));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(clk32MHz), .D(n17700));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(clk32MHz), .D(n17699));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1132 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[9] [4]), .I3(n35566), .O(n35587));
    defparam i2_3_lut_4_lut_adj_1132.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1133 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[9] [2]), 
            .I2(n16714), .I3(n16772), .O(n30582));
    defparam i2_3_lut_4_lut_adj_1133.LUT_INIT = 16'h6996;
    SB_LUT4 mux_1080_i14_3_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n4385), .I3(GND_net), .O(n4399));
    defparam mux_1080_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(clk32MHz), .D(n17698));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(clk32MHz), .D(n17697));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(clk32MHz), .D(n17696));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(clk32MHz), .D(n17695));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(clk32MHz), .D(n17694));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(clk32MHz), .D(n17693));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(clk32MHz), .D(n17692));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i2_2_lut_3_lut (.I0(\data_in_frame[18] [3]), .I1(n35536), .I2(\data_in_frame[20] [1]), 
            .I3(GND_net), .O(n10_adj_4311));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1134 (.I0(\data_in_frame[18] [3]), .I1(n35536), 
            .I2(\data_in_frame[21] [0]), .I3(GND_net), .O(n35508));
    defparam i1_2_lut_3_lut_adj_1134.LUT_INIT = 16'h9696;
    SB_LUT4 i29_3_lut_4_lut (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[12] [1]), 
            .I2(\data_in_frame[20] [0]), .I3(n35638), .O(n86));
    defparam i29_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1135 (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[12] [1]), 
            .I2(\data_in_frame[11] [7]), .I3(GND_net), .O(n8_adj_4312));
    defparam i1_2_lut_3_lut_adj_1135.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1136 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[18] [0]), 
            .I2(n16184), .I3(n35318), .O(n36368));
    defparam i2_3_lut_4_lut_adj_1136.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1137 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[18] [0]), 
            .I2(n35521), .I3(n35297), .O(n31017));
    defparam i2_3_lut_4_lut_adj_1137.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_4_lut (.I0(n35426), .I1(n35230), .I2(n35376), .I3(\data_out_frame[15] [7]), 
            .O(n8_adj_4313));
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1138 (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state[1] ), 
            .I2(\FRAME_MATCHER.state_31__N_2725 [3]), .I3(\FRAME_MATCHER.state [2]), 
            .O(n6_adj_4314));   // verilog/coms.v(145[4] 294[11])
    defparam i2_3_lut_4_lut_adj_1138.LUT_INIT = 16'h00bf;
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(clk32MHz), 
           .D(n18022));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1139 (.I0(n63_c), .I1(n63_adj_4315), .I2(n63), 
            .I3(GND_net), .O(n10389));   // verilog/coms.v(139[4] 141[7])
    defparam i1_2_lut_3_lut_adj_1139.LUT_INIT = 16'h8080;
    SB_LUT4 i19380_2_lut_3_lut (.I0(n63_c), .I1(n63_adj_4315), .I2(\FRAME_MATCHER.state[1] ), 
            .I3(GND_net), .O(n23[1]));   // verilog/coms.v(139[4] 141[7])
    defparam i19380_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_3_lut_adj_1140 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [31]), 
            .I3(GND_net), .O(n34465));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1140.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1141 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [30]), 
            .I3(GND_net), .O(n7_adj_4317));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1141.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1142 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [29]), 
            .I3(GND_net), .O(n7_adj_4318));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1142.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1143 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [28]), 
            .I3(GND_net), .O(n34451));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1143.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1144 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [27]), 
            .I3(GND_net), .O(n34463));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1144.LUT_INIT = 16'he0e0;
    SB_LUT4 mux_1080_i13_3_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n4385), .I3(GND_net), .O(n4398));
    defparam mux_1080_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1145 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [26]), 
            .I3(GND_net), .O(n34461));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1145.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut (.I0(\byte_transmit_counter[4] ), 
            .I1(\byte_transmit_counter[3] ), .I2(n38672), .I3(n38671), 
            .O(tx_data[3]));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1_2_lut_3_lut_adj_1146 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [25]), 
            .I3(GND_net), .O(n7_adj_4319));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1146.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1147 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [24]), 
            .I3(GND_net), .O(n34459));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1147.LUT_INIT = 16'he0e0;
    SB_LUT4 mux_1080_i16_3_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n4385), .I3(GND_net), .O(n4401));
    defparam mux_1080_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13372_3_lut_4_lut (.I0(n8_adj_4320), .I1(n35006), .I2(rx_data[1]), 
            .I3(\data_in_frame[22] [1]), .O(n18111));
    defparam i13372_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1148 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [23]), 
            .I3(GND_net), .O(n34457));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1148.LUT_INIT = 16'he0e0;
    SB_LUT4 mux_1080_i15_3_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n4385), .I3(GND_net), .O(n4400));
    defparam mux_1080_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1080_i18_3_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n4385), .I3(GND_net), .O(n4403));
    defparam mux_1080_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1149 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [22]), 
            .I3(GND_net), .O(n34469));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1149.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1150 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [21]), 
            .I3(GND_net), .O(n7_adj_4321));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1150.LUT_INIT = 16'he0e0;
    SB_LUT4 i13371_3_lut_4_lut (.I0(n8_adj_4320), .I1(n35006), .I2(rx_data[0]), 
            .I3(\data_in_frame[22] [0]), .O(n18110));
    defparam i13371_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1151 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [20]), 
            .I3(GND_net), .O(n34449));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1151.LUT_INIT = 16'he0e0;
    SB_LUT4 i13374_3_lut_4_lut (.I0(n8_adj_4320), .I1(n35006), .I2(rx_data[3]), 
            .I3(\data_in_frame[22] [3]), .O(n18113));
    defparam i13374_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1152 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [19]), 
            .I3(GND_net), .O(n7_adj_4322));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1152.LUT_INIT = 16'he0e0;
    SB_LUT4 i13373_3_lut_4_lut (.I0(n8_adj_4320), .I1(n35006), .I2(rx_data[2]), 
            .I3(\data_in_frame[22] [2]), .O(n18112));
    defparam i13373_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [6]), .I2(\data_out_frame[19] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n43805));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n43805_bdd_4_lut (.I0(n43805), .I1(\data_out_frame[17] [6]), 
            .I2(\data_out_frame[16] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n43808));
    defparam n43805_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36934 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [5]), .I2(\data_out_frame[19] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n43799));
    defparam byte_transmit_counter_0__bdd_4_lut_36934.LUT_INIT = 16'he4aa;
    SB_LUT4 n43799_bdd_4_lut (.I0(n43799), .I1(\data_out_frame[17] [5]), 
            .I2(\data_out_frame[16] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n43802));
    defparam n43799_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36929 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [4]), .I2(\data_out_frame[19] [4]), 
            .I3(\byte_transmit_counter[1] ), .O(n43793));
    defparam byte_transmit_counter_0__bdd_4_lut_36929.LUT_INIT = 16'he4aa;
    SB_LUT4 n43793_bdd_4_lut (.I0(n43793), .I1(\data_out_frame[17] [4]), 
            .I2(\data_out_frame[16] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n43796));
    defparam n43793_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mux_1080_i17_3_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n4385), .I3(GND_net), .O(n4402));
    defparam mux_1080_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19198_2_lut_3_lut (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [18]), 
            .I3(GND_net), .O(n23914));   // verilog/coms.v(114[11:12])
    defparam i19198_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i13376_3_lut_4_lut (.I0(n8_adj_4320), .I1(n35006), .I2(rx_data[5]), 
            .I3(\data_in_frame[22] [5]), .O(n18115));
    defparam i13376_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i19197_2_lut_3_lut (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [17]), 
            .I3(GND_net), .O(n23912));   // verilog/coms.v(114[11:12])
    defparam i19197_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(clk32MHz), 
            .D(n2_adj_4323), .S(n3_adj_4324));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(clk32MHz), 
           .D(n18000));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1153 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [16]), 
            .I3(GND_net), .O(n34447));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1153.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1154 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [15]), 
            .I3(GND_net), .O(n34445));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1154.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1155 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [14]), 
            .I3(GND_net), .O(n34455));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1155.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1156 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [13]), 
            .I3(GND_net), .O(n34443));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1156.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1157 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [12]), 
            .I3(GND_net), .O(n34467));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1157.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1158 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [11]), 
            .I3(GND_net), .O(n34441));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1158.LUT_INIT = 16'he0e0;
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(clk32MHz), 
           .D(n18021));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(clk32MHz), 
           .D(n18020));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(clk32MHz), 
           .D(n18019));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(clk32MHz), 
           .D(n18018));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(clk32MHz), 
           .D(n18017));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(clk32MHz), 
            .D(n2_adj_4325), .S(n3_adj_4326));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13375_3_lut_4_lut (.I0(n8_adj_4320), .I1(n35006), .I2(rx_data[4]), 
            .I3(\data_in_frame[22] [4]), .O(n18114));
    defparam i13375_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1159 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [10]), 
            .I3(GND_net), .O(n34429));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1159.LUT_INIT = 16'he0e0;
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(clk32MHz), 
            .D(n2_adj_4327), .S(n3_adj_4328));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(clk32MHz), 
            .D(n2_adj_4329), .S(n3_adj_4330));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(clk32MHz), 
            .D(n2_adj_4331), .S(n3_adj_4332));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(clk32MHz), 
            .D(n2_adj_4333), .S(n3_adj_4334));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(clk32MHz), 
            .D(n2_adj_4335), .S(n3_adj_4336));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(clk32MHz), 
            .D(n2_adj_4337), .S(n3_adj_4338));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(clk32MHz), 
            .D(n2_adj_4339), .S(n3_adj_4340));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(clk32MHz), 
            .D(n2_adj_4341), .S(n3_adj_4342));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(clk32MHz), 
            .D(n2_adj_4343), .S(n3_adj_4344));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(clk32MHz), 
            .D(n2_adj_4345), .S(n3_adj_4346));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(clk32MHz), 
            .D(n2_adj_4347), .S(n3_adj_4348));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(clk32MHz), 
            .D(n2_adj_4349), .S(n3_adj_4350));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(clk32MHz), 
            .D(n2_adj_4351), .S(n3_adj_4352));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(clk32MHz), 
            .D(n2_adj_4353), .S(n3_adj_4354));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(clk32MHz), 
            .D(n2_adj_4355), .S(n3_adj_4356));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(clk32MHz), 
            .D(n2_adj_4357), .S(n3_adj_4358));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(clk32MHz), 
            .D(n2_adj_4359), .S(n3_adj_4360));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(clk32MHz), 
            .D(n2_adj_4361), .S(n3_adj_4362));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(clk32MHz), 
            .D(n2_adj_4363), .S(n3_adj_4364));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(clk32MHz), 
            .D(n2_adj_4365), .S(n3_adj_4366));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(clk32MHz), 
            .D(n2_adj_4367), .S(n3_adj_4368));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(clk32MHz), 
            .D(n2_adj_4369), .S(n3_adj_4370));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(clk32MHz), 
            .D(n2_adj_4371), .S(n3_adj_4372));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(clk32MHz), 
            .D(n2_adj_4373), .S(n3_adj_4374));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(clk32MHz), 
            .D(n2_adj_4375), .S(n3_adj_4376));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(clk32MHz), 
            .D(n2_adj_4377), .S(n3_adj_4378));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(clk32MHz), 
            .D(n2_adj_4379), .S(n3_adj_4380));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(clk32MHz), 
            .D(n2_adj_4381), .S(n3_adj_4382));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i [31]), .C(clk32MHz), 
            .D(n2_adj_4383), .S(n3_adj_4384));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(clk32MHz), 
           .D(n18016));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1160 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [9]), 
            .I3(GND_net), .O(n34453));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1160.LUT_INIT = 16'he0e0;
    SB_DFFE data_out_frame_0___i169 (.Q(\data_out_frame[21] [0]), .C(clk32MHz), 
            .E(n17205), .D(n36265));   // verilog/coms.v(127[12] 295[6])
    SB_DFFE data_out_frame_0___i170 (.Q(\data_out_frame[21] [1]), .C(clk32MHz), 
            .E(n17205), .D(n36416));   // verilog/coms.v(127[12] 295[6])
    SB_DFFE data_out_frame_0___i171 (.Q(\data_out_frame[21] [2]), .C(clk32MHz), 
            .E(n17205), .D(n37044));   // verilog/coms.v(127[12] 295[6])
    SB_DFFE data_out_frame_0___i172 (.Q(\data_out_frame[21] [3]), .C(clk32MHz), 
            .E(n17205), .D(n36758));   // verilog/coms.v(127[12] 295[6])
    SB_DFFE data_out_frame_0___i173 (.Q(\data_out_frame[21] [4]), .C(clk32MHz), 
            .E(n17205), .D(n36181));   // verilog/coms.v(127[12] 295[6])
    SB_DFFE data_out_frame_0___i174 (.Q(\data_out_frame[21] [5]), .C(clk32MHz), 
            .E(n17205), .D(n36199));   // verilog/coms.v(127[12] 295[6])
    SB_DFFE data_out_frame_0___i175 (.Q(\data_out_frame[21] [6]), .C(clk32MHz), 
            .E(n17205), .D(n37556));   // verilog/coms.v(127[12] 295[6])
    SB_DFFE data_out_frame_0___i176 (.Q(\data_out_frame[21] [7]), .C(clk32MHz), 
            .E(n17205), .D(n36904));   // verilog/coms.v(127[12] 295[6])
    SB_DFFE data_out_frame_0___i177 (.Q(\data_out_frame[22] [0]), .C(clk32MHz), 
            .E(n17205), .D(n35353));   // verilog/coms.v(127[12] 295[6])
    SB_DFFE data_out_frame_0___i178 (.Q(\data_out_frame[22] [1]), .C(clk32MHz), 
            .E(n17205), .D(n35271));   // verilog/coms.v(127[12] 295[6])
    SB_DFFE data_out_frame_0___i179 (.Q(\data_out_frame[22] [2]), .C(clk32MHz), 
            .E(n17205), .D(n36143));   // verilog/coms.v(127[12] 295[6])
    SB_DFFE data_out_frame_0___i180 (.Q(\data_out_frame[22] [3]), .C(clk32MHz), 
            .E(n17205), .D(n36260));   // verilog/coms.v(127[12] 295[6])
    SB_DFFE data_out_frame_0___i181 (.Q(\data_out_frame[22] [4]), .C(clk32MHz), 
            .E(n17205), .D(n35383));   // verilog/coms.v(127[12] 295[6])
    SB_DFFE data_out_frame_0___i182 (.Q(\data_out_frame[22] [5]), .C(clk32MHz), 
            .E(n17205), .D(n36345));   // verilog/coms.v(127[12] 295[6])
    SB_DFFE data_out_frame_0___i183 (.Q(\data_out_frame[22] [6]), .C(clk32MHz), 
            .E(n17205), .D(n36347));   // verilog/coms.v(127[12] 295[6])
    SB_DFFE data_out_frame_0___i184 (.Q(\data_out_frame[22] [7]), .C(clk32MHz), 
            .E(n17205), .D(n37510));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(clk32MHz), 
           .D(n18015));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1161 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [8]), 
            .I3(GND_net), .O(n34439));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1161.LUT_INIT = 16'he0e0;
    SB_DFFESR LED_3497 (.Q(LED_c), .C(clk32MHz), .E(n34927), .D(n17348), 
            .R(n37152));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state[1] ), .C(clk32MHz), 
            .D(n34329), .S(n44032));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1162 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [7]), 
            .I3(GND_net), .O(n34437));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1162.LUT_INIT = 16'he0e0;
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state[3] ), .C(clk32MHz), 
            .D(n34333), .S(n10_adj_4385));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state [4]), .C(clk32MHz), 
            .D(n34431), .S(n34331));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state [5]), .C(clk32MHz), 
            .D(n34433), .S(n34397));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state [6]), .C(clk32MHz), 
            .D(n34435), .S(n34395));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state [7]), .C(clk32MHz), 
            .D(n34437), .S(n34393));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state [8]), .C(clk32MHz), 
            .D(n34439), .S(n34391));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state [9]), .C(clk32MHz), 
            .D(n34453), .S(n34335));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state [10]), .C(clk32MHz), 
            .D(n34429), .S(n34401));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state [11]), .C(clk32MHz), 
            .D(n34441), .S(n34389));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state [12]), .C(clk32MHz), 
            .D(n34467), .S(n34339));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state [13]), .C(clk32MHz), 
            .D(n34443), .S(n34387));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state [14]), .C(clk32MHz), 
            .D(n34455), .S(n34351));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state [15]), .C(clk32MHz), 
            .D(n34445), .S(n34385));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state [16]), .C(clk32MHz), 
            .D(n34447), .S(n34383));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state [17]), .C(clk32MHz), 
            .D(n23912), .S(n24679));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state [18]), .C(clk32MHz), 
            .D(n23914), .S(n24681));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state [19]), .C(clk32MHz), 
            .D(n7_adj_4322), .S(n8_adj_4386));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state [20]), .C(clk32MHz), 
            .D(n34449), .S(n34381));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state [21]), .C(clk32MHz), 
            .D(n7_adj_4321), .S(n8_adj_4387));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state [22]), .C(clk32MHz), 
            .D(n34469), .S(n34349));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state [23]), .C(clk32MHz), 
            .D(n34457), .S(n34347));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state [24]), .C(clk32MHz), 
            .D(n34459), .S(n34345));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state [25]), .C(clk32MHz), 
            .D(n7_adj_4319), .S(n34273));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state [26]), .C(clk32MHz), 
            .D(n34461), .S(n34337));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state [27]), .C(clk32MHz), 
            .D(n34463), .S(n34341));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state [28]), .C(clk32MHz), 
            .D(n34451), .S(n34379));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state [29]), .C(clk32MHz), 
            .D(n7_adj_4318), .S(n8_adj_4388));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state [30]), .C(clk32MHz), 
            .D(n7_adj_4317), .S(n8_adj_4389));   // verilog/coms.v(127[12] 295[6])
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state [31]), .C(clk32MHz), 
            .D(n34465), .S(n34323));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13378_3_lut_4_lut (.I0(n8_adj_4320), .I1(n35006), .I2(rx_data[7]), 
            .I3(\data_in_frame[22] [7]), .O(n18117));
    defparam i13378_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1163 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [6]), 
            .I3(GND_net), .O(n34435));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1163.LUT_INIT = 16'he0e0;
    SB_LUT4 mux_1080_i20_3_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n4385), .I3(GND_net), .O(n4405));
    defparam mux_1080_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13377_3_lut_4_lut (.I0(n8_adj_4320), .I1(n35006), .I2(rx_data[6]), 
            .I3(\data_in_frame[22] [6]), .O(n18116));
    defparam i13377_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1164 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [5]), 
            .I3(GND_net), .O(n34433));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1164.LUT_INIT = 16'he0e0;
    SB_LUT4 i13227_3_lut_4_lut (.I0(n8), .I1(n34998), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n17966));
    defparam i13227_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1165 (.I0(n70), .I1(n67), .I2(\FRAME_MATCHER.state [4]), 
            .I3(GND_net), .O(n34431));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1165.LUT_INIT = 16'he0e0;
    SB_LUT4 mux_1080_i19_3_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n4385), .I3(GND_net), .O(n4404));
    defparam mux_1080_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut (.I0(n15_adj_4390), .I1(n46), .I2(n1), .I3(\FRAME_MATCHER.state [30]), 
            .O(n8_adj_4389));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1166 (.I0(n15_adj_4390), .I1(n46), .I2(n1), 
            .I3(\FRAME_MATCHER.state [29]), .O(n8_adj_4388));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_4_lut_adj_1166.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1167 (.I0(n15_adj_4390), .I1(n46), .I2(n1), 
            .I3(\FRAME_MATCHER.state [25]), .O(n34273));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_4_lut_adj_1167.LUT_INIT = 16'hfe00;
    SB_LUT4 mux_1080_i22_3_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n4385), .I3(GND_net), .O(n4407));
    defparam mux_1080_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_4_lut_adj_1168 (.I0(n15_adj_4390), .I1(n46), .I2(n1), 
            .I3(\FRAME_MATCHER.state [21]), .O(n8_adj_4387));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_4_lut_adj_1168.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_4_lut_adj_1169 (.I0(n15_adj_4390), .I1(n46), .I2(n1), 
            .I3(\FRAME_MATCHER.state [19]), .O(n8_adj_4386));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_4_lut_adj_1169.LUT_INIT = 16'hfe00;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36924 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [3]), .I2(\data_out_frame[19] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n43787));
    defparam byte_transmit_counter_0__bdd_4_lut_36924.LUT_INIT = 16'he4aa;
    SB_LUT4 i19960_2_lut_4_lut (.I0(n15_adj_4390), .I1(n46), .I2(n1), 
            .I3(\FRAME_MATCHER.state [18]), .O(n24681));   // verilog/coms.v(114[11:12])
    defparam i19960_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i19959_2_lut_4_lut (.I0(n15_adj_4390), .I1(n46), .I2(n1), 
            .I3(\FRAME_MATCHER.state [17]), .O(n24679));   // verilog/coms.v(114[11:12])
    defparam i19959_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i13228_3_lut_4_lut (.I0(n8), .I1(n34998), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n17967));
    defparam i13228_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1170 (.I0(\data_in_frame[21] [7]), .I1(\data_in_frame[21] [6]), 
            .I2(n35157), .I3(GND_net), .O(n35466));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_3_lut_adj_1170.LUT_INIT = 16'h9696;
    SB_LUT4 i13229_3_lut_4_lut (.I0(n8), .I1(n34998), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n17968));
    defparam i13229_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1171 (.I0(\data_in_frame[21] [7]), .I1(\data_in_frame[21] [6]), 
            .I2(n35218), .I3(\data_in_frame[21] [5]), .O(Kp_23__N_1802));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i13267_3_lut_4_lut (.I0(n8_adj_4391), .I1(n34984), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n18006));
    defparam i13267_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13268_3_lut_4_lut (.I0(n8_adj_4391), .I1(n34984), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n18007));
    defparam i13268_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13269_3_lut_4_lut (.I0(n8_adj_4391), .I1(n34984), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n18008));
    defparam i13269_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13270_3_lut_4_lut (.I0(n8_adj_4391), .I1(n34984), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n18009));
    defparam i13270_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13230_3_lut_4_lut (.I0(n8), .I1(n34998), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n17969));
    defparam i13230_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13271_3_lut_4_lut (.I0(n8_adj_4391), .I1(n34984), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n18010));
    defparam i13271_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13272_3_lut_4_lut (.I0(n8_adj_4391), .I1(n34984), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n18011));
    defparam i13272_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13273_3_lut_4_lut (.I0(n8_adj_4391), .I1(n34984), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n18012));
    defparam i13273_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13274_3_lut_4_lut (.I0(n8_adj_4391), .I1(n34984), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n18013));
    defparam i13274_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut (.I0(\byte_transmit_counter[4] ), 
            .I1(\byte_transmit_counter[3] ), .I2(n38663), .I3(n38662), 
            .O(tx_data[0]));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i13231_3_lut_4_lut (.I0(n8), .I1(n34998), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n17970));
    defparam i13231_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1080_i21_3_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n4385), .I3(GND_net), .O(n4406));
    defparam mux_1080_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1172 (.I0(\data_in[2] [6]), .I1(\data_in[1] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4392));
    defparam i1_2_lut_adj_1172.LUT_INIT = 16'hdddd;
    SB_LUT4 i4_4_lut_adj_1173 (.I0(\data_in[0] [5]), .I1(\data_in[1] [6]), 
            .I2(\data_in[3] [7]), .I3(n6_adj_4392), .O(n37642));
    defparam i4_4_lut_adj_1173.LUT_INIT = 16'hffbf;
    SB_LUT4 add_44_2_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i7_4_lut_adj_1174 (.I0(n9_adj_4393), .I1(n14_adj_4305), .I2(n36539), 
            .I3(n17011), .O(n35144));   // verilog/coms.v(74[16:43])
    defparam i7_4_lut_adj_1174.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1175 (.I0(\data_in_frame[11] [5]), .I1(n35144), 
            .I2(\data_in_frame[9] [4]), .I3(GND_net), .O(n30683));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1175.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(clk32MHz), 
           .D(n18014));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(clk32MHz), 
           .D(n18013));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i3_4_lut_adj_1176 (.I0(\data_in[1] [3]), .I1(\data_in[2] [5]), 
            .I2(n15939), .I3(\data_in[0] [1]), .O(n37335));
    defparam i3_4_lut_adj_1176.LUT_INIT = 16'hfffe;
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(clk32MHz), 
           .D(n18066));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i3_4_lut_adj_1177 (.I0(n37335), .I1(n37642), .I2(\data_in[2] [0]), 
            .I3(\data_in[3] [2]), .O(n15759));
    defparam i3_4_lut_adj_1177.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut_adj_1178 (.I0(n15848), .I1(\data_in[3] [3]), .I2(\data_in[2] [1]), 
            .I3(\data_in[3] [6]), .O(n16_adj_4394));
    defparam i6_4_lut_adj_1178.LUT_INIT = 16'hffbf;
    SB_LUT4 i13232_3_lut_4_lut (.I0(n8), .I1(n34998), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n17971));
    defparam i13232_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1179 (.I0(\data_in[2] [3]), .I1(n15759), .I2(\data_in[3] [5]), 
            .I3(\data_in[0] [7]), .O(n17_adj_4395));
    defparam i7_4_lut_adj_1179.LUT_INIT = 16'hffdf;
    SB_LUT4 i13315_3_lut_4_lut (.I0(n24712), .I1(n34984), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n18054));
    defparam i13315_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i9_4_lut_adj_1180 (.I0(n17_adj_4395), .I1(\data_in[0] [2]), 
            .I2(n16_adj_4394), .I3(\data_in[3] [1]), .O(n63_c));
    defparam i9_4_lut_adj_1180.LUT_INIT = 16'hfbff;
    SB_LUT4 i13316_3_lut_4_lut (.I0(n24712), .I1(n34984), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n18055));
    defparam i13316_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(clk32MHz), 
           .D(n18065));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i6_4_lut_adj_1181 (.I0(\data_in[3] [0]), .I1(n15858), .I2(n15759), 
            .I3(\data_in[2] [2]), .O(n16_adj_4396));
    defparam i6_4_lut_adj_1181.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1182 (.I0(\data_in[2] [4]), .I1(\data_in[1] [0]), 
            .I2(\data_in[1] [5]), .I3(\data_in[0] [3]), .O(n17_adj_4397));
    defparam i7_4_lut_adj_1182.LUT_INIT = 16'hfffd;
    SB_LUT4 i13317_3_lut_4_lut (.I0(n24712), .I1(n34984), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n18056));
    defparam i13317_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13318_3_lut_4_lut (.I0(n24712), .I1(n34984), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n18057));
    defparam i13318_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13319_3_lut_4_lut (.I0(n24712), .I1(n34984), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n18058));
    defparam i13319_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13320_3_lut_4_lut (.I0(n24712), .I1(n34984), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n18059));
    defparam i13320_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13321_3_lut_4_lut (.I0(n24712), .I1(n34984), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n18060));
    defparam i13321_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13322_3_lut_4_lut (.I0(n24712), .I1(n34984), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n18061));
    defparam i13322_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13233_3_lut_4_lut (.I0(n8), .I1(n34998), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n17972));
    defparam i13233_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut (.I0(n15460), .I1(n37527), .I2(\data_in_frame[19] [6]), 
            .I3(GND_net), .O(n6));
    defparam i1_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_1183 (.I0(n7), .I1(n37314), .I2(\data_in_frame[17] [6]), 
            .I3(n31476), .O(n35300));
    defparam i4_4_lut_adj_1183.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1184 (.I0(\data_in_frame[20] [0]), .I1(n15460), 
            .I2(GND_net), .I3(GND_net), .O(n30523));
    defparam i1_2_lut_adj_1184.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(clk32MHz), 
           .D(n18064));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13234_3_lut_4_lut (.I0(n8), .I1(n34998), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n17973));
    defparam i13234_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(clk32MHz), 
           .D(n18012));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(clk32MHz), 
           .D(n18063));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i9_4_lut_adj_1185 (.I0(n17_adj_4397), .I1(\data_in[0] [6]), 
            .I2(n16_adj_4396), .I3(\data_in[1] [4]), .O(n63_adj_4315));
    defparam i9_4_lut_adj_1185.LUT_INIT = 16'hfbff;
    SB_DFF setpoint__i0 (.Q(setpoint[0]), .C(clk32MHz), .D(n17616));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(clk32MHz), 
           .D(n18062));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(clk32MHz), 
           .D(n18061));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(clk32MHz), 
           .D(n18060));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(clk32MHz), 
           .D(n18059));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(clk32MHz), 
           .D(n18058));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(clk32MHz), 
           .D(n18011));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(clk32MHz), 
           .D(n18010));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(clk32MHz), 
           .D(n18009));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(clk32MHz), 
           .D(n18008));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i1_4_lut_adj_1186 (.I0(n30683), .I1(\data_in_frame[16] [0]), 
            .I2(n35082), .I3(\data_in_frame[15] [7]), .O(n31530));
    defparam i1_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_LUT4 i13302_3_lut_4_lut (.I0(n8_adj_4260), .I1(n34984), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n18041));
    defparam i13302_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1187 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [3]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4398));
    defparam i1_2_lut_adj_1187.LUT_INIT = 16'h8888;
    SB_LUT4 i19340_4_lut (.I0(n8_adj_4399), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n15845), .I3(n4_adj_4398), .O(n3894));   // verilog/coms.v(251[9:58])
    defparam i19340_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i33651_2_lut (.I0(\byte_transmit_counter[2] ), .I1(\byte_transmit_counter[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n40522));
    defparam i33651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_adj_1188 (.I0(\byte_transmit_counter[7] ), .I1(byte_transmit_counter[6]), 
            .I2(\byte_transmit_counter[5] ), .I3(GND_net), .O(n5_adj_4264));
    defparam i2_3_lut_adj_1188.LUT_INIT = 16'hfefe;
    SB_LUT4 i13303_3_lut_4_lut (.I0(n8_adj_4260), .I1(n34984), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n18042));
    defparam i13303_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13304_3_lut_4_lut (.I0(n8_adj_4260), .I1(n34984), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n18043));
    defparam i13304_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1189 (.I0(n31476), .I1(\data_in_frame[17] [6]), 
            .I2(n35575), .I3(\data_in_frame[17] [7]), .O(n15460));
    defparam i3_4_lut_adj_1189.LUT_INIT = 16'h6996;
    SB_LUT4 n43787_bdd_4_lut (.I0(n43787), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[16] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n43790));
    defparam n43787_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_44_33_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [31]), .I2(GND_net), 
            .I3(n27914), .O(n2_adj_4383)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_44_32_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n27913), .O(n2_adj_4381)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_32_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_32 (.CI(n27913), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n27914));
    SB_LUT4 add_44_31_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n27912), .O(n2_adj_4379)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_31_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(clk32MHz), 
           .D(n17999));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13305_3_lut_4_lut (.I0(n8_adj_4260), .I1(n34984), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n18044));
    defparam i13305_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13306_3_lut_4_lut (.I0(n8_adj_4260), .I1(n34984), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n18045));
    defparam i13306_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i36753_2_lut (.I0(n24966), .I1(n5_adj_4264), .I2(GND_net), 
            .I3(GND_net), .O(tx_transmit_N_3482));
    defparam i36753_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i19333_4_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [31]), 
            .I2(n4_adj_4400), .I3(\FRAME_MATCHER.i [1]), .O(n788));   // verilog/coms.v(157[9:60])
    defparam i19333_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i13301_3_lut_4_lut (.I0(n8_adj_4260), .I1(n34984), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n18040));
    defparam i13301_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13299_3_lut_4_lut (.I0(n8_adj_4260), .I1(n34984), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n18038));
    defparam i13299_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13300_3_lut_4_lut (.I0(n8_adj_4260), .I1(n34984), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n18039));
    defparam i13300_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13291_3_lut_4_lut (.I0(n8), .I1(n34984), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n18030));
    defparam i13291_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13292_3_lut_4_lut (.I0(n8), .I1(n34984), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n18031));
    defparam i13292_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut (.I0(\FRAME_MATCHER.state[1] ), .I1(n15722), 
            .I2(n9_adj_4401), .I3(n1), .O(n12_adj_4402));   // verilog/coms.v(151[5:27])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hff10;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(\byte_transmit_counter[1] ), 
            .I1(n19_adj_4403), .I2(n40680), .I3(\byte_transmit_counter[2] ), 
            .O(n43781));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 i13293_3_lut_4_lut (.I0(n8), .I1(n34984), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n18032));
    defparam i13293_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4355_2_lut (.I0(n63), .I1(n788), .I2(GND_net), .I3(GND_net), 
            .O(n9015));   // verilog/coms.v(157[6] 159[9])
    defparam i4355_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_44_31 (.CI(n27912), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n27913));
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1190 (.I0(n30671), .I1(n16876), .I2(GND_net), 
            .I3(GND_net), .O(n35388));
    defparam i1_2_lut_adj_1190.LUT_INIT = 16'h6666;
    SB_LUT4 i13294_3_lut_4_lut (.I0(n8), .I1(n34984), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n18033));
    defparam i13294_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i16_4_lut_adj_1191 (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42));
    defparam i16_4_lut_adj_1191.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1192 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41));
    defparam i15_4_lut_adj_1192.LUT_INIT = 16'hfffe;
    SB_LUT4 equal_103_i7_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4404));   // verilog/coms.v(154[7:23])
    defparam equal_103_i7_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i14_4_lut_adj_1193 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40));
    defparam i14_4_lut_adj_1193.LUT_INIT = 16'hfffe;
    SB_LUT4 n43781_bdd_4_lut (.I0(n43781), .I1(n17_adj_4405), .I2(n16_adj_4406), 
            .I3(\byte_transmit_counter[2] ), .O(n43784));
    defparam n43781_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39));
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13295_3_lut_4_lut (.I0(n8), .I1(n34984), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n18034));
    defparam i13295_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43), .I2(n42), .I3(n44), .O(n50));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n45), .I1(n50), .I2(n39), .I3(n40), .O(n15845));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1194 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [3]), 
            .I2(n15845), .I3(GND_net), .O(n15765));
    defparam i2_3_lut_adj_1194.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(n15992), .I1(n10389), .I2(n101), 
            .I3(tx_transmit_N_3482), .O(n70));   // verilog/coms.v(207[5:16])
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h4440;
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(clk32MHz), 
           .D(n18007));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(clk32MHz), 
           .D(n18006));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13296_3_lut_4_lut (.I0(n8), .I1(n34984), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n18035));
    defparam i13296_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(clk32MHz), 
           .D(n18005));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(clk32MHz), 
           .D(n18004));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(clk32MHz), 
           .D(n18003));   // verilog/coms.v(127[12] 295[6])
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state [0]), .C(clk32MHz), 
           .D(n34343));   // verilog/coms.v(127[12] 295[6])
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(clk32MHz), .D(n17593));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(clk32MHz), 
           .D(n17592));   // verilog/coms.v(127[12] 295[6])
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(clk32MHz), .D(n17591));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 add_44_30_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n27911), .O(n2_adj_4377)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_30_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(clk32MHz), .D(n17590));   // verilog/coms.v(127[12] 295[6])
    SB_CARRY add_44_30 (.CI(n27911), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n27912));
    SB_LUT4 add_44_29_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n27910), .O(n2_adj_4375)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_29_lut.LUT_INIT = 16'h8228;
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(clk32MHz), .D(n17589));   // verilog/coms.v(127[12] 295[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(clk32MHz), .D(n17588));   // verilog/coms.v(127[12] 295[6])
    SB_DFF gearBoxRatio_i0_i0 (.Q(gearBoxRatio[0]), .C(clk32MHz), .D(n17587));   // verilog/coms.v(127[12] 295[6])
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(clk32MHz), .D(n17445));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13297_3_lut_4_lut (.I0(n8), .I1(n34984), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n18036));
    defparam i13297_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13298_3_lut_4_lut (.I0(n8), .I1(n34984), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n18037));
    defparam i13298_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6][7] ), .C(clk32MHz), 
           .D(n17989));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(clk32MHz), 
           .D(n18057));   // verilog/coms.v(127[12] 295[6])
    SB_CARRY add_44_29 (.CI(n27910), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n27911));
    SB_LUT4 add_44_28_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n27909), .O(n2_adj_4373)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_28_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_28 (.CI(n27909), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n27910));
    SB_LUT4 add_44_27_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n27908), .O(n2_adj_4371)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_27_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_27 (.CI(n27908), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n27909));
    SB_LUT4 add_44_26_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n27907), .O(n2_adj_4369)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_26 (.CI(n27907), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n27908));
    SB_LUT4 add_44_25_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n27906), .O(n2_adj_4367)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_25_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_25 (.CI(n27906), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n27907));
    SB_LUT4 add_44_24_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n27905), .O(n2_adj_4365)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13354_3_lut_4_lut (.I0(n8_adj_4407), .I1(n35006), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n18093));
    defparam i13354_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_24 (.CI(n27905), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n27906));
    SB_LUT4 i13347_3_lut_4_lut (.I0(n8_adj_4407), .I1(n35006), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n18086));
    defparam i13347_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13219_3_lut_4_lut (.I0(n8_adj_4407), .I1(n34998), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n17958));
    defparam i13219_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_23_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n27904), .O(n2_adj_4363)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_23 (.CI(n27904), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n27905));
    SB_LUT4 i4_4_lut_adj_1195 (.I0(\data_in_frame[6][7] ), .I1(n16777), 
            .I2(n35558), .I3(n6_adj_4408), .O(n31571));
    defparam i4_4_lut_adj_1195.LUT_INIT = 16'h6996;
    SB_LUT4 add_44_22_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n27903), .O(n2_adj_4361)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_22 (.CI(n27903), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n27904));
    SB_LUT4 i13348_3_lut_4_lut (.I0(n8_adj_4407), .I1(n35006), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n18087));
    defparam i13348_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_21_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n27902), .O(n2_adj_4359)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_21_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_21 (.CI(n27902), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n27903));
    SB_LUT4 add_44_20_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n27901), .O(n2_adj_4357)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13349_3_lut_4_lut (.I0(n8_adj_4407), .I1(n35006), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n18088));
    defparam i13349_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_20 (.CI(n27901), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n27902));
    SB_LUT4 add_44_19_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n27900), .O(n2_adj_4355)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13350_3_lut_4_lut (.I0(n8_adj_4407), .I1(n35006), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n18089));
    defparam i13350_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_19 (.CI(n27900), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n27901));
    SB_LUT4 add_44_18_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n27899), .O(n2_adj_4353)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13351_3_lut_4_lut (.I0(n8_adj_4407), .I1(n35006), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n18090));
    defparam i13351_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13352_3_lut_4_lut (.I0(n8_adj_4407), .I1(n35006), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n18091));
    defparam i13352_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_44_18 (.CI(n27899), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n27900));
    SB_LUT4 i13353_3_lut_4_lut (.I0(n8_adj_4407), .I1(n35006), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n18092));
    defparam i13353_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_44_17_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n27898), .O(n2_adj_4351)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_17_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_17 (.CI(n27898), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n27899));
    SB_LUT4 add_44_16_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n27897), .O(n2_adj_4349)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_16_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_16 (.CI(n27897), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n27898));
    SB_LUT4 add_44_15_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n27896), .O(n2_adj_4347)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_15 (.CI(n27896), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n27897));
    SB_LUT4 add_44_14_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n27895), .O(n2_adj_4345)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_14_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_14 (.CI(n27895), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n27896));
    SB_LUT4 add_44_13_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n27894), .O(n2_adj_4343)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i3_4_lut_adj_1196 (.I0(\data_in_frame[11] [4]), .I1(n31571), 
            .I2(\data_in_frame[11] [3]), .I3(n31118), .O(n35249));
    defparam i3_4_lut_adj_1196.LUT_INIT = 16'h6996;
    SB_CARRY add_44_13 (.CI(n27894), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n27895));
    SB_LUT4 add_44_12_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n27893), .O(n2_adj_4341)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_12 (.CI(n27893), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n27894));
    SB_LUT4 add_44_11_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n27892), .O(n2_adj_4339)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i2_2_lut_adj_1197 (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4409));
    defparam i2_2_lut_adj_1197.LUT_INIT = 16'heeee;
    SB_CARRY add_44_11 (.CI(n27892), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n27893));
    SB_LUT4 add_44_10_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n27891), .O(n2_adj_4337)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i6_4_lut_adj_1198 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_4410));
    defparam i6_4_lut_adj_1198.LUT_INIT = 16'hfeff;
    SB_CARRY add_44_10 (.CI(n27891), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n27892));
    SB_LUT4 i13220_3_lut_4_lut (.I0(n8_adj_4407), .I1(n34998), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n17959));
    defparam i13220_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1199 (.I0(\data_in[3] [6]), .I1(n14_adj_4410), 
            .I2(n10_adj_4409), .I3(\data_in[2] [1]), .O(n15858));
    defparam i7_4_lut_adj_1199.LUT_INIT = 16'hfffd;
    SB_LUT4 add_44_9_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n27890), .O(n2_adj_4335)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_4_lut_adj_1200 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_4411));
    defparam i4_4_lut_adj_1200.LUT_INIT = 16'hfdff;
    SB_LUT4 i3_4_lut_adj_1201 (.I0(\data_in_frame[15] [6]), .I1(n31457), 
            .I2(n35067), .I3(\data_in_frame[11] [2]), .O(n35082));
    defparam i3_4_lut_adj_1201.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1202 (.I0(\data_in[3] [4]), .I1(n10_adj_4411), 
            .I2(\data_in[2] [7]), .I3(GND_net), .O(n15939));
    defparam i5_3_lut_adj_1202.LUT_INIT = 16'hdfdf;
    SB_LUT4 i31794_4_lut (.I0(\data_in[1] [5]), .I1(\data_in[1] [0]), .I2(\data_in[2] [2]), 
            .I3(\data_in[0] [3]), .O(n38564));
    defparam i31794_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_adj_1203 (.I0(\data_in[2] [4]), .I1(\data_in[1] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4412));
    defparam i1_2_lut_adj_1203.LUT_INIT = 16'heeee;
    SB_CARRY add_44_9 (.CI(n27890), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n27891));
    SB_LUT4 add_44_8_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n27889), .O(n2_adj_4333)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_8_lut.LUT_INIT = 16'h8228;
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(clk32MHz), 
           .D(n18056));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(clk32MHz), 
           .D(n18055));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(clk32MHz), 
           .D(n18054));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(clk32MHz), 
           .D(n18002));   // verilog/coms.v(127[12] 295[6])
    SB_CARRY add_44_8 (.CI(n27889), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n27890));
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(clk32MHz), 
           .D(n18001));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(clk32MHz), 
           .D(n18053));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(clk32MHz), 
           .D(n18052));   // verilog/coms.v(127[12] 295[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(clk32MHz), 
           .D(n18051));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i13221_3_lut_4_lut (.I0(n8_adj_4407), .I1(n34998), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n17960));
    defparam i13221_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(clk32MHz), 
           .D(n18050));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i7_4_lut_adj_1204 (.I0(n9_adj_4412), .I1(n38564), .I2(\data_in[3] [0]), 
            .I3(\data_in[0] [6]), .O(n15848));
    defparam i7_4_lut_adj_1204.LUT_INIT = 16'hffbf;
    SB_LUT4 add_44_7_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n27888), .O(n2_adj_4331)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_7 (.CI(n27888), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n27889));
    SB_LUT4 i13222_3_lut_4_lut (.I0(n8_adj_4407), .I1(n34998), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n17961));
    defparam i13222_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i31770_2_lut (.I0(\data_in[2] [0]), .I1(\data_in[1] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n38538));
    defparam i31770_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_44_6_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n27887), .O(n2_adj_4329)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_6_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_6 (.CI(n27887), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n27888));
    SB_LUT4 add_44_5_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n27886), .O(n2_adj_4327)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_5 (.CI(n27886), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n27887));
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(clk32MHz), 
           .D(n18049));   // verilog/coms.v(127[12] 295[6])
    SB_LUT4 i8_4_lut_adj_1205 (.I0(n15848), .I1(n15939), .I2(\data_in[3] [7]), 
            .I3(\data_in[2] [6]), .O(n21_adj_4413));
    defparam i8_4_lut_adj_1205.LUT_INIT = 16'hfffe;
    SB_LUT4 add_44_4_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n27885), .O(n2_adj_4325)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i7_3_lut_adj_1206 (.I0(\data_in[0] [1]), .I1(\data_in[2] [5]), 
            .I2(\data_in[1] [6]), .I3(GND_net), .O(n20_adj_4414));
    defparam i7_3_lut_adj_1206.LUT_INIT = 16'hf7f7;
    SB_CARRY add_44_4 (.CI(n27885), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n27886));
    SB_LUT4 add_44_3_lut (.I0(n2058), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n27884), .O(n2_adj_4323)) /* synthesis syn_instantiated=1 */ ;
    defparam add_44_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_44_3 (.CI(n27884), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n27885));
    SB_LUT4 i11_4_lut_adj_1207 (.I0(n21_adj_4413), .I1(n15858), .I2(n38538), 
            .I3(\data_in[0] [5]), .O(n24_adj_4415));
    defparam i11_4_lut_adj_1207.LUT_INIT = 16'hefff;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36919 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [2]), .I2(\data_out_frame[19] [2]), 
            .I3(\byte_transmit_counter[1] ), .O(n43775));
    defparam byte_transmit_counter_0__bdd_4_lut_36919.LUT_INIT = 16'he4aa;
    SB_LUT4 i12_4_lut_adj_1208 (.I0(\data_in[3] [2]), .I1(n24_adj_4415), 
            .I2(n20_adj_4414), .I3(\data_in[1] [2]), .O(n63));
    defparam i12_4_lut_adj_1208.LUT_INIT = 16'hfdff;
    SB_LUT4 i3_4_lut_adj_1209 (.I0(n23947), .I1(n43_adj_4416), .I2(n15950), 
            .I3(n24684), .O(n2774));
    defparam i3_4_lut_adj_1209.LUT_INIT = 16'h8000;
    SB_LUT4 i13223_3_lut_4_lut (.I0(n8_adj_4407), .I1(n34998), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n17962));
    defparam i13223_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i19460_3_lut (.I0(\FRAME_MATCHER.state [2]), .I1(n63_adj_4315), 
            .I2(n63_c), .I3(GND_net), .O(n122));   // verilog/coms.v(139[4] 141[7])
    defparam i19460_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 select_368_Select_2_i5_4_lut (.I0(n122), .I1(n15957), .I2(n2957), 
            .I3(n63), .O(n5));
    defparam select_368_Select_2_i5_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i19463_rep_228_2_lut (.I0(n122), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(n44342));   // verilog/coms.v(142[4] 144[7])
    defparam i19463_rep_228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13224_3_lut_4_lut (.I0(n8_adj_4407), .I1(n34998), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n17963));
    defparam i13224_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13225_3_lut_4_lut (.I0(n8_adj_4407), .I1(n34998), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n17964));
    defparam i13225_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13226_3_lut_4_lut (.I0(n8_adj_4407), .I1(n34998), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n17965));
    defparam i13226_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n43775_bdd_4_lut (.I0(n43775), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(\byte_transmit_counter[1] ), 
            .O(n43778));
    defparam n43775_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36910 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [0]), .I2(\data_out_frame[11] [0]), 
            .I3(\byte_transmit_counter[1] ), .O(n43769));
    defparam byte_transmit_counter_0__bdd_4_lut_36910.LUT_INIT = 16'he4aa;
    SB_LUT4 n43769_bdd_4_lut (.I0(n43769), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[8] [0]), .I3(\byte_transmit_counter[1] ), 
            .O(n43772));
    defparam n43769_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36905 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [0]), .I2(\data_out_frame[15] [0]), 
            .I3(\byte_transmit_counter[1] ), .O(n43763));
    defparam byte_transmit_counter_0__bdd_4_lut_36905.LUT_INIT = 16'he4aa;
    SB_LUT4 n43763_bdd_4_lut (.I0(n43763), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[12] [0]), .I3(\byte_transmit_counter[1] ), 
            .O(n43766));
    defparam n43763_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36900 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [1]), .I2(\data_out_frame[11] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n43757));
    defparam byte_transmit_counter_0__bdd_4_lut_36900.LUT_INIT = 16'he4aa;
    SB_LUT4 i13310_3_lut_4_lut (.I0(n8_adj_4320), .I1(n34984), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n18049));
    defparam i13310_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13311_3_lut_4_lut (.I0(n8_adj_4320), .I1(n34984), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n18050));
    defparam i13311_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13312_3_lut_4_lut (.I0(n8_adj_4320), .I1(n34984), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n18051));
    defparam i13312_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n16386), .I1(\data_in_frame[5] [3]), 
            .I2(n15531), .I3(n30669), .O(n35644));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1210 (.I0(n16386), .I1(\data_in_frame[5] [3]), 
            .I2(n15531), .I3(\data_in_frame[7] [4]), .O(n30578));
    defparam i1_2_lut_3_lut_4_lut_adj_1210.LUT_INIT = 16'h6996;
    SB_LUT4 i13313_3_lut_4_lut (.I0(n8_adj_4320), .I1(n34984), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n18052));
    defparam i13313_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n43757_bdd_4_lut (.I0(n43757), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n43760));
    defparam n43757_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1211 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[6] [2]), 
            .I2(n16115), .I3(\data_in_frame[6] [0]), .O(n35641));   // verilog/coms.v(84[17:63])
    defparam i1_2_lut_4_lut_adj_1211.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(n16812), .I3(n16876), .O(n10_adj_4267));
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1212 (.I0(\data_in_frame[4] [6]), .I1(n5_adj_4288), 
            .I2(n6_adj_4289), .I3(n17011), .O(n35391));
    defparam i1_2_lut_3_lut_4_lut_adj_1212.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1213 (.I0(n16231), .I1(\data_in_frame[10] [4]), 
            .I2(n16642), .I3(n35185), .O(n30512));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1213.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1214 (.I0(\data_out_frame[16] [5]), .I1(n37560), 
            .I2(n36894), .I3(GND_net), .O(n6_adj_4418));
    defparam i2_2_lut_3_lut_adj_1214.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36895 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [1]), .I2(\data_out_frame[15] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n43751));
    defparam byte_transmit_counter_0__bdd_4_lut_36895.LUT_INIT = 16'he4aa;
    SB_LUT4 i13314_3_lut_4_lut (.I0(n8_adj_4320), .I1(n34984), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n18053));
    defparam i13314_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13307_3_lut_4_lut (.I0(n8_adj_4320), .I1(n34984), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n18046));
    defparam i13307_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13308_3_lut_4_lut (.I0(n8_adj_4320), .I1(n34984), .I2(rx_data[1]), 
            .I3(\data_in_frame[14][1] ), .O(n18047));
    defparam i13308_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n43751_bdd_4_lut (.I0(n43751), .I1(\data_out_frame[13] [1]), 
            .I2(\data_out_frame[12] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n43754));
    defparam n43751_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36890 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [2]), .I2(\data_out_frame[11] [2]), 
            .I3(\byte_transmit_counter[1] ), .O(n43745));
    defparam byte_transmit_counter_0__bdd_4_lut_36890.LUT_INIT = 16'he4aa;
    SB_LUT4 n43745_bdd_4_lut (.I0(n43745), .I1(\data_out_frame[9] [2]), 
            .I2(\data_out_frame[8] [2]), .I3(\byte_transmit_counter[1] ), 
            .O(n43748));
    defparam n43745_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36885 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [2]), .I2(\data_out_frame[15] [2]), 
            .I3(\byte_transmit_counter[1] ), .O(n43739));
    defparam byte_transmit_counter_0__bdd_4_lut_36885.LUT_INIT = 16'he4aa;
    SB_LUT4 n43739_bdd_4_lut (.I0(n43739), .I1(\data_out_frame[13] [2]), 
            .I2(\data_out_frame[12] [2]), .I3(\byte_transmit_counter[1] ), 
            .O(n43742));
    defparam n43739_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_3_lut_4_lut_adj_1215 (.I0(\data_out_frame[13] [6]), .I1(n30704), 
            .I2(\data_out_frame[9] [6]), .I3(\data_out_frame[9] [7]), .O(n14_adj_4419));
    defparam i5_3_lut_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36880 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [3]), .I2(\data_out_frame[11] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n43733));
    defparam byte_transmit_counter_0__bdd_4_lut_36880.LUT_INIT = 16'he4aa;
    SB_LUT4 n43733_bdd_4_lut (.I0(n43733), .I1(\data_out_frame[9] [3]), 
            .I2(\data_out_frame[8] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n43736));
    defparam n43733_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13309_3_lut_4_lut (.I0(n8_adj_4320), .I1(n34984), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n18048));
    defparam i13309_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i19472_2_lut (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n24190));
    defparam i19472_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36875 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [3]), .I2(\data_out_frame[15] [3]), 
            .I3(\byte_transmit_counter[1] ), .O(n43727));
    defparam byte_transmit_counter_0__bdd_4_lut_36875.LUT_INIT = 16'he4aa;
    SB_LUT4 n43727_bdd_4_lut (.I0(n43727), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[12] [3]), .I3(\byte_transmit_counter[1] ), 
            .O(n43730));
    defparam n43727_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1216 (.I0(\FRAME_MATCHER.state [6]), .I1(\FRAME_MATCHER.state [5]), 
            .I2(\FRAME_MATCHER.state [4]), .I3(\FRAME_MATCHER.state [7]), 
            .O(n24686));
    defparam i3_4_lut_adj_1216.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36870 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [4]), .I2(\data_out_frame[11] [4]), 
            .I3(\byte_transmit_counter[1] ), .O(n43721));
    defparam byte_transmit_counter_0__bdd_4_lut_36870.LUT_INIT = 16'he4aa;
    SB_LUT4 n43721_bdd_4_lut (.I0(n43721), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[8] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n43724));
    defparam n43721_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i4_2_lut (.I0(\FRAME_MATCHER.state [29]), .I1(\FRAME_MATCHER.state [22]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4420));   // verilog/coms.v(151[5:27])
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36865 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [1]), .I2(\data_out_frame[19] [1]), 
            .I3(\byte_transmit_counter[1] ), .O(n43715));
    defparam byte_transmit_counter_0__bdd_4_lut_36865.LUT_INIT = 16'he4aa;
    SB_LUT4 n43715_bdd_4_lut (.I0(n43715), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(\byte_transmit_counter[1] ), 
            .O(n43718));
    defparam n43715_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i10_4_lut_adj_1217 (.I0(\FRAME_MATCHER.state [16]), .I1(\FRAME_MATCHER.state [19]), 
            .I2(\FRAME_MATCHER.state [23]), .I3(\FRAME_MATCHER.state [26]), 
            .O(n24_adj_4421));   // verilog/coms.v(151[5:27])
    defparam i10_4_lut_adj_1217.LUT_INIT = 16'hfffe;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36860 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [0]), .I2(\data_out_frame[19] [0]), 
            .I3(\byte_transmit_counter[1] ), .O(n43709));
    defparam byte_transmit_counter_0__bdd_4_lut_36860.LUT_INIT = 16'he4aa;
    SB_LUT4 n43709_bdd_4_lut (.I0(n43709), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(\byte_transmit_counter[1] ), 
            .O(n43712));
    defparam n43709_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i8_4_lut_adj_1218 (.I0(\FRAME_MATCHER.state [21]), .I1(\FRAME_MATCHER.state [30]), 
            .I2(\FRAME_MATCHER.state [18]), .I3(\FRAME_MATCHER.state [27]), 
            .O(n22_adj_4422));   // verilog/coms.v(151[5:27])
    defparam i8_4_lut_adj_1218.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1219 (.I0(n37132), .I1(n35367), .I2(\data_in_frame[18] [4]), 
            .I3(n31558), .O(n36436));
    defparam i2_3_lut_4_lut_adj_1219.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1220 (.I0(n30704), .I1(n16870), .I2(n35125), 
            .I3(n16587), .O(n6_adj_4423));
    defparam i1_2_lut_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1221 (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[5] [4]), 
            .I2(\data_out_frame[5] [3]), .I3(\data_out_frame[7] [5]), .O(n35057));
    defparam i1_2_lut_4_lut_adj_1221.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1222 (.I0(\data_out_frame[11] [6]), .I1(\data_out_frame[7] [5]), 
            .I2(\data_out_frame[5] [5]), .I3(\data_out_frame[11] [7]), .O(n35651));   // verilog/coms.v(84[17:28])
    defparam i2_3_lut_4_lut_adj_1222.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1223 (.I0(n37132), .I1(n35367), .I2(n35188), 
            .I3(\data_in_frame[21] [0]), .O(n14_adj_4281));
    defparam i5_3_lut_4_lut_adj_1223.LUT_INIT = 16'h9669;
    SB_LUT4 i13211_3_lut_4_lut (.I0(n10_adj_4424), .I1(n34995), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n17950));
    defparam i13211_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_3_lut_4_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n8_adj_4399), .I3(n38499), .O(n36526));   // verilog/coms.v(154[7:23])
    defparam i3_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 equal_109_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4425));   // verilog/coms.v(154[7:23])
    defparam equal_109_i10_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i4_4_lut_adj_1224 (.I0(\data_in_frame[15] [4]), .I1(n16645), 
            .I2(n35429), .I3(n6_adj_4259), .O(n31476));
    defparam i4_4_lut_adj_1224.LUT_INIT = 16'h6996;
    SB_LUT4 i20272_2_lut (.I0(n15886), .I1(n15963), .I2(GND_net), .I3(GND_net), 
            .O(n4498));
    defparam i20272_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1225 (.I0(r_SM_Main_2__N_3585[0]), .I1(tx_active), 
            .I2(GND_net), .I3(GND_net), .O(n101));
    defparam i1_2_lut_adj_1225.LUT_INIT = 16'heeee;
    SB_LUT4 i13212_3_lut_4_lut (.I0(n10_adj_4424), .I1(n34995), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n17951));
    defparam i13212_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13213_3_lut_4_lut (.I0(n10_adj_4424), .I1(n34995), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n17952));
    defparam i13213_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15025_3_lut (.I0(byte_transmit_counter[6]), .I1(n40622), .I2(n24918), 
            .I3(GND_net), .O(n18288));
    defparam i15025_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i13214_3_lut_4_lut (.I0(n10_adj_4424), .I1(n34995), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n17953));
    defparam i13214_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1226 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[7] [1]), 
            .I2(\data_out_frame[7] [2]), .I3(\data_out_frame[5] [1]), .O(n1286));   // verilog/coms.v(84[17:70])
    defparam i2_3_lut_4_lut_adj_1226.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1227 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[5] [4]), .I3(GND_net), .O(n16937));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_1227.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1228 (.I0(n30598), .I1(\data_out_frame[14] [4]), 
            .I2(\data_out_frame[14] [3]), .I3(GND_net), .O(n35422));
    defparam i1_2_lut_3_lut_adj_1228.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36855 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [4]), .I2(\data_out_frame[15] [4]), 
            .I3(\byte_transmit_counter[1] ), .O(n43703));
    defparam byte_transmit_counter_0__bdd_4_lut_36855.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1229 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[7] [3]), .I3(GND_net), .O(n35490));
    defparam i1_2_lut_3_lut_adj_1229.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1230 (.I0(n16239), .I1(\data_out_frame[5] [7]), 
            .I2(n35141), .I3(GND_net), .O(n14107));
    defparam i1_2_lut_3_lut_adj_1230.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1231 (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(\data_out_frame[15] [0]), .I3(GND_net), .O(n35654));
    defparam i1_2_lut_3_lut_adj_1231.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1232 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[6] [2]), .I3(GND_net), .O(n16239));
    defparam i1_2_lut_3_lut_adj_1232.LUT_INIT = 16'h9696;
    SB_LUT4 i13215_3_lut_4_lut (.I0(n10_adj_4424), .I1(n34995), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n17954));
    defparam i13215_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1233 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[6] [2]), .I3(GND_net), .O(n35141));
    defparam i1_2_lut_3_lut_adj_1233.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1234 (.I0(n30598), .I1(n16214), .I2(n35565), 
            .I3(\data_out_frame[16] [7]), .O(n35635));
    defparam i2_3_lut_4_lut_adj_1234.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1235 (.I0(\data_in_frame[10] [5]), .I1(\data_in_frame[10] [6]), 
            .I2(\data_in_frame[12] [7]), .I3(GND_net), .O(n35212));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1235.LUT_INIT = 16'h9696;
    SB_LUT4 n43703_bdd_4_lut (.I0(n43703), .I1(\data_out_frame[13] [4]), 
            .I2(\data_out_frame[12] [4]), .I3(\byte_transmit_counter[1] ), 
            .O(n43706));
    defparam n43703_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_3_lut_adj_1236 (.I0(\data_in_frame[9] [3]), .I1(n35249), 
            .I2(\data_in_frame[13] [5]), .I3(GND_net), .O(n30689));
    defparam i2_3_lut_adj_1236.LUT_INIT = 16'h9696;
    SB_LUT4 i3_3_lut_4_lut_adj_1237 (.I0(\data_out_frame[5] [7]), .I1(n35141), 
            .I2(n35475), .I3(n35596), .O(n8_adj_4426));
    defparam i3_3_lut_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1238 (.I0(n30558), .I1(\data_out_frame[13] [0]), 
            .I2(n35565), .I3(\data_out_frame[14] [7]), .O(n35475));
    defparam i1_2_lut_4_lut_adj_1238.LUT_INIT = 16'h9669;
    SB_LUT4 i12_4_lut_adj_1239 (.I0(\FRAME_MATCHER.state [17]), .I1(n24_adj_4421), 
            .I2(n18_adj_4420), .I3(\FRAME_MATCHER.state [20]), .O(n26_adj_4427));   // verilog/coms.v(151[5:27])
    defparam i12_4_lut_adj_1239.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_4_lut_adj_1240 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[6] [3]), 
            .I2(\data_out_frame[10] [6]), .I3(\data_out_frame[6] [4]), .O(n35596));
    defparam i2_3_lut_4_lut_adj_1240.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1241 (.I0(n30558), .I1(\data_out_frame[13] [0]), 
            .I2(n35565), .I3(GND_net), .O(n35566));
    defparam i1_2_lut_3_lut_adj_1241.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36850 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [5]), .I2(\data_out_frame[11] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n43697));
    defparam byte_transmit_counter_0__bdd_4_lut_36850.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1242 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[10] [5]), 
            .I2(\data_out_frame[12] [7]), .I3(GND_net), .O(n6_adj_4428));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_3_lut_adj_1242.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1243 (.I0(\data_out_frame[17] [4]), .I1(n35151), 
            .I2(\data_out_frame[20] [0]), .I3(GND_net), .O(n35530));
    defparam i1_2_lut_3_lut_adj_1243.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1244 (.I0(\data_in_frame[10] [5]), .I1(n16231), 
            .I2(n16645), .I3(\data_in_frame[12] [7]), .O(n35135));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1244.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_3_lut_4_lut (.I0(n16115), .I1(\data_in_frame[7] [6]), 
            .I2(\data_in_frame[7] [5]), .I3(\data_in_frame[9] [7]), .O(n16_adj_4429));
    defparam i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1245 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[8] [7]), .I3(\data_out_frame[6] [5]), .O(n7_adj_4430));
    defparam i1_3_lut_4_lut_adj_1245.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1246 (.I0(\data_out_frame[13] [4]), .I1(\data_out_frame[7] [0]), 
            .I2(n16772), .I3(GND_net), .O(n8_adj_4431));
    defparam i2_2_lut_3_lut_adj_1246.LUT_INIT = 16'h9696;
    SB_LUT4 i13216_3_lut_4_lut (.I0(n10_adj_4424), .I1(n34995), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n17955));
    defparam i13216_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n43697_bdd_4_lut (.I0(n43697), .I1(\data_out_frame[9] [5]), 
            .I2(\data_out_frame[8] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n43700));
    defparam n43697_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i13217_3_lut_4_lut (.I0(n10_adj_4424), .I1(n34995), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n17956));
    defparam i13217_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1247 (.I0(tx_transmit_N_3482), .I1(n101), 
            .I2(n15992), .I3(GND_net), .O(n3));   // verilog/coms.v(209[11:56])
    defparam i1_2_lut_3_lut_adj_1247.LUT_INIT = 16'h0e0e;
    SB_LUT4 i11_3_lut_adj_1248 (.I0(\FRAME_MATCHER.state [31]), .I1(n22_adj_4422), 
            .I2(\FRAME_MATCHER.state [24]), .I3(GND_net), .O(n25_adj_4433));   // verilog/coms.v(151[5:27])
    defparam i11_3_lut_adj_1248.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_1249 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[6] [6]), 
            .I2(n35432), .I3(\data_out_frame[11] [2]), .O(n16772));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_LUT4 i13218_3_lut_4_lut (.I0(n10_adj_4424), .I1(n34995), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n17957));
    defparam i13218_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut (.I0(\byte_transmit_counter[4] ), 
            .I1(\byte_transmit_counter[3] ), .I2(n38666), .I3(n38665), 
            .O(tx_data[1]));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 mux_1080_i9_3_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n4385), .I3(GND_net), .O(n4394));
    defparam mux_1080_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1250 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [2]), 
            .I2(n1286), .I3(n16714), .O(n30545));
    defparam i2_3_lut_4_lut_adj_1250.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1251 (.I0(\data_out_frame[7] [0]), .I1(\data_out_frame[7] [1]), 
            .I2(\data_out_frame[6] [6]), .I3(\data_out_frame[5] [0]), .O(n16714));   // verilog/coms.v(84[17:70])
    defparam i2_3_lut_4_lut_adj_1251.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1252 (.I0(\data_out_frame[13] [2]), .I1(n31254), 
            .I2(\data_out_frame[15] [4]), .I3(GND_net), .O(n35107));
    defparam i1_2_lut_3_lut_adj_1252.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1253 (.I0(n31610), .I1(n30653), .I2(\data_in_frame[16] [5]), 
            .I3(GND_net), .O(n17023));
    defparam i1_2_lut_3_lut_adj_1253.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1254 (.I0(n31455), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[17] [7]), .I3(GND_net), .O(n35081));
    defparam i1_2_lut_3_lut_adj_1254.LUT_INIT = 16'h9696;
    SB_LUT4 mux_1080_i8_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n4385), .I3(GND_net), .O(n4393));
    defparam mux_1080_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1080_i7_3_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n4385), .I3(GND_net), .O(n4392));
    defparam mux_1080_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1255 (.I0(\data_in_frame[17] [7]), .I1(n37314), 
            .I2(n31530), .I3(n35575), .O(n36755));
    defparam i2_3_lut_4_lut_adj_1255.LUT_INIT = 16'h6996;
    SB_LUT4 i13283_3_lut_4_lut (.I0(n8_adj_4407), .I1(n34984), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n18022));
    defparam i13283_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1256 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[18] [2]), 
            .I2(n16566), .I3(n36894), .O(n35285));
    defparam i2_3_lut_4_lut_adj_1256.LUT_INIT = 16'h9669;
    SB_LUT4 mux_1080_i6_3_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n4385), .I3(GND_net), .O(n4391));
    defparam mux_1080_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1080_i5_3_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n4385), .I3(GND_net), .O(n4390));
    defparam mux_1080_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1080_i4_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n4385), .I3(GND_net), .O(n4389));
    defparam mux_1080_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1257 (.I0(n31455), .I1(n35079), .I2(\data_out_frame[18] [2]), 
            .I3(n30516), .O(n35297));
    defparam i2_3_lut_4_lut_adj_1257.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1258 (.I0(\FRAME_MATCHER.state [0]), .I1(n63_adj_4315), 
            .I2(n63_c), .I3(n63), .O(\FRAME_MATCHER.state_31__N_2661[0] ));
    defparam i3_4_lut_adj_1258.LUT_INIT = 16'hbfff;
    SB_LUT4 i13284_3_lut_4_lut (.I0(n8_adj_4407), .I1(n34984), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n18023));
    defparam i13284_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1259 (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(n34984), .O(n34989));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1259.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_3_lut_adj_1260 (.I0(\data_out_frame[20] [2]), .I1(n16566), 
            .I2(n30667), .I3(GND_net), .O(n6_adj_4434));
    defparam i1_2_lut_3_lut_adj_1260.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1261 (.I0(n35081), .I1(\data_out_frame[18] [2]), 
            .I2(n30516), .I3(n35524), .O(n35525));
    defparam i1_2_lut_4_lut_adj_1261.LUT_INIT = 16'h9669;
    SB_LUT4 mux_1080_i3_3_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n4385), .I3(GND_net), .O(n4388));
    defparam mux_1080_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1262 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[20] [4]), 
            .I2(n31518), .I3(n35285), .O(n36347));
    defparam i2_3_lut_4_lut_adj_1262.LUT_INIT = 16'h6996;
    SB_LUT4 i36749_2_lut_3_lut (.I0(\FRAME_MATCHER.state[1] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n17348));
    defparam i36749_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i1_4_lut_3_lut (.I0(\FRAME_MATCHER.state [0]), .I1(\FRAME_MATCHER.state [2]), 
            .I2(n26), .I3(GND_net), .O(n5_adj_4435));
    defparam i1_4_lut_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i13285_3_lut_4_lut (.I0(n8_adj_4407), .I1(n34984), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n18024));
    defparam i13285_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1263 (.I0(n35671), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n15886), .I3(n15963), .O(n15861));
    defparam i1_3_lut_4_lut_adj_1263.LUT_INIT = 16'haaae;
    SB_LUT4 i1_3_lut_4_lut_adj_1264 (.I0(\FRAME_MATCHER.state[3] ), .I1(n10389), 
            .I2(n2774), .I3(n67), .O(n34333));
    defparam i1_3_lut_4_lut_adj_1264.LUT_INIT = 16'haa80;
    SB_LUT4 i1_2_lut_3_lut_adj_1265 (.I0(\data_in_frame[21] [0]), .I1(\data_in_frame[22] [7]), 
            .I2(\data_in_frame[22] [6]), .I3(GND_net), .O(n35493));
    defparam i1_2_lut_3_lut_adj_1265.LUT_INIT = 16'h9696;
    SB_LUT4 i77_2_lut_3_lut (.I0(n2957), .I1(n10389), .I2(n15957), .I3(GND_net), 
            .O(n46));   // verilog/coms.v(114[11:12])
    defparam i77_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i13286_3_lut_4_lut (.I0(n8_adj_4407), .I1(n34984), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n18025));
    defparam i13286_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1266 (.I0(n788), .I1(n10389), .I2(n15960), 
            .I3(GND_net), .O(n15_adj_4390));   // verilog/coms.v(114[11:12])
    defparam i1_2_lut_3_lut_adj_1266.LUT_INIT = 16'h0404;
    SB_LUT4 i13329_3_lut_4_lut (.I0(n8_adj_4399), .I1(n35006), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n18068));
    defparam i13329_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1267 (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[18] [6]), 
            .I2(\data_in_frame[19] [0]), .I3(GND_net), .O(n35188));
    defparam i1_2_lut_3_lut_adj_1267.LUT_INIT = 16'h9696;
    SB_LUT4 i13287_3_lut_4_lut (.I0(n8_adj_4407), .I1(n34984), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n18026));
    defparam i13287_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 \FRAME_MATCHER.state_31__I_0_3579_i64_1_lut_2_lut_3_lut  (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(n15963), .I2(n24738), .I3(GND_net), .O(\FRAME_MATCHER.i_31__N_2624 ));   // verilog/coms.v(207[5:16])
    defparam \FRAME_MATCHER.state_31__I_0_3579_i64_1_lut_2_lut_3_lut .LUT_INIT = 16'h1010;
    SB_LUT4 i1_3_lut_4_lut_adj_1268 (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[20] [6]), 
            .I2(n31558), .I3(n30721), .O(n7_adj_4436));
    defparam i1_3_lut_4_lut_adj_1268.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_4_lut_adj_1269 (.I0(n31476), .I1(\data_in_frame[17] [2]), 
            .I2(\data_in_frame[17] [3]), .I3(\data_in_frame[19] [6]), .O(n14_adj_4437));
    defparam i5_3_lut_4_lut_adj_1269.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1270 (.I0(n30588), .I1(\data_in_frame[20] [0]), 
            .I2(n15460), .I3(GND_net), .O(n6_adj_4438));
    defparam i1_2_lut_3_lut_adj_1270.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1271 (.I0(\data_in_frame[11] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(n10_adj_4439), .I3(\data_in_frame[11] [1]), .O(n37314));
    defparam i5_3_lut_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1272 (.I0(\data_in_frame[1] [7]), .I1(n35413), 
            .I2(n16142), .I3(n35091), .O(n6_adj_4440));   // verilog/coms.v(84[17:63])
    defparam i1_2_lut_4_lut_adj_1272.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i16_3_lut (.I0(\data_out_frame[16] [7]), 
            .I1(\data_out_frame[17] [7]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n16_adj_4406));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i17_3_lut (.I0(\data_out_frame[18] [7]), 
            .I1(\data_out_frame[19] [7]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n17_adj_4405));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34239_2_lut (.I0(\data_out_frame[22] [7]), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n40680));
    defparam i34239_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i19_3_lut (.I0(\data_out_frame[20] [7]), 
            .I1(\data_out_frame[21] [7]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4403));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19231_2_lut_3_lut_4_lut (.I0(n15992), .I1(\FRAME_MATCHER.state[3] ), 
            .I2(n15886), .I3(n15963), .O(n23947));
    defparam i19231_2_lut_3_lut_4_lut.LUT_INIT = 16'haaa2;
    SB_LUT4 i13288_3_lut_4_lut (.I0(n8_adj_4407), .I1(n34984), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n18027));
    defparam i13288_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1273 (.I0(n30689), .I1(n35082), .I2(GND_net), 
            .I3(GND_net), .O(n35575));
    defparam i1_2_lut_adj_1273.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1274 (.I0(\data_in_frame[17] [7]), .I1(n37314), 
            .I2(n30689), .I3(n35082), .O(n30588));
    defparam i1_2_lut_3_lut_4_lut_adj_1274.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut (.I0(\byte_transmit_counter[4] ), 
            .I1(\byte_transmit_counter[3] ), .I2(n38669), .I3(n38668), 
            .O(tx_data[2]));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i2_2_lut_3_lut_adj_1275 (.I0(\FRAME_MATCHER.state[3] ), .I1(n15886), 
            .I2(n15963), .I3(GND_net), .O(n63_adj_3));   // verilog/coms.v(196[5:24])
    defparam i2_2_lut_3_lut_adj_1275.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_3_lut_adj_1276 (.I0(\FRAME_MATCHER.state[3] ), .I1(n15963), 
            .I2(n24738), .I3(GND_net), .O(n15992));   // verilog/coms.v(207[5:16])
    defparam i1_2_lut_3_lut_adj_1276.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_adj_1277 (.I0(\data_in_frame[7] [1]), .I1(n16777), 
            .I2(GND_net), .I3(GND_net), .O(n35562));
    defparam i1_2_lut_adj_1277.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1278 (.I0(n16953), .I1(n35562), .I2(n30669), 
            .I3(\data_in_frame[6] [6]), .O(n12_adj_4442));
    defparam i5_4_lut_adj_1278.LUT_INIT = 16'h6996;
    SB_LUT4 i20017_2_lut_3_lut (.I0(\FRAME_MATCHER.state[1] ), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(GND_net), .O(n24738));
    defparam i20017_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_4_lut_adj_1279 (.I0(\data_in_frame[8] [6]), .I1(n16156), 
            .I2(\data_in_frame[6] [4]), .I3(\data_in_frame[6] [5]), .O(n16883));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1279.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1280 (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(n15963), .I2(\FRAME_MATCHER.state[1] ), .I3(n15958), .O(n15994));   // verilog/coms.v(246[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1280.LUT_INIT = 16'hffef;
    SB_LUT4 i13289_3_lut_4_lut (.I0(n8_adj_4407), .I1(n34984), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n18028));
    defparam i13289_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1281 (.I0(\FRAME_MATCHER.state[3] ), 
            .I1(n15963), .I2(\FRAME_MATCHER.state[1] ), .I3(\FRAME_MATCHER.state [0]), 
            .O(n43_adj_4416));   // verilog/coms.v(246[5:25])
    defparam i1_2_lut_3_lut_4_lut_adj_1281.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1282 (.I0(n37132), .I1(n30592), .I2(\data_in_frame[16] [2]), 
            .I3(n30807), .O(n35536));
    defparam i1_2_lut_3_lut_4_lut_adj_1282.LUT_INIT = 16'h9669;
    SB_LUT4 mux_1080_i1_3_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n4385), .I3(GND_net), .O(n4386));
    defparam mux_1080_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i13290_3_lut_4_lut (.I0(n8_adj_4407), .I1(n34984), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n18029));
    defparam i13290_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1283 (.I0(\data_in_frame[7] [0]), .I1(n12_adj_4442), 
            .I2(\data_in_frame[9] [2]), .I3(n35391), .O(n36539));
    defparam i6_4_lut_adj_1283.LUT_INIT = 16'h6996;
    SB_LUT4 i13203_3_lut_4_lut (.I0(n8_adj_4391), .I1(n34998), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n17942));
    defparam i13203_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i34261_2_lut (.I0(\byte_transmit_counter[2] ), .I1(\data_out_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n41108));   // verilog/coms.v(105[34:55])
    defparam i34261_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i5_3_lut (.I0(\data_out_frame[6] [7]), 
            .I1(\data_out_frame[7] [7]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4443));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1080_i24_3_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n4385), .I3(GND_net), .O(n4409));
    defparam mux_1080_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31803_4_lut (.I0(n5_adj_4443), .I1(n41108), .I2(n40522), 
            .I3(\byte_transmit_counter[0] ), .O(n38649));
    defparam i31803_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i31805_4_lut (.I0(n38649), .I1(n43784), .I2(\byte_transmit_counter[4] ), 
            .I3(\byte_transmit_counter[3] ), .O(n38651));
    defparam i31805_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31804_3_lut (.I0(n43670), .I1(n43664), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n38650));
    defparam i31804_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i19_3_lut (.I0(\data_out_frame[20] [6]), 
            .I1(\data_out_frame[21] [6]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4444));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34257_2_lut (.I0(\byte_transmit_counter[2] ), .I1(\data_out_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n41104));   // verilog/coms.v(105[34:55])
    defparam i34257_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i5_3_lut (.I0(\data_out_frame[6] [6]), 
            .I1(\data_out_frame[7] [6]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4445));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1284 (.I0(\data_in_frame[11] [3]), .I1(\data_in_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35067));
    defparam i1_2_lut_adj_1284.LUT_INIT = 16'h6666;
    SB_LUT4 i31849_4_lut (.I0(n19_adj_4444), .I1(\data_out_frame[22] [6]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n38695));
    defparam i31849_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31850_3_lut (.I0(n43808), .I1(n38695), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n38696));
    defparam i31850_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31833_4_lut (.I0(n5_adj_4445), .I1(n41104), .I2(n40522), 
            .I3(\byte_transmit_counter[0] ), .O(n38679));
    defparam i31833_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i31835_4_lut (.I0(n38679), .I1(n38696), .I2(\byte_transmit_counter[4] ), 
            .I3(\byte_transmit_counter[3] ), .O(n38681));
    defparam i31835_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31834_3_lut (.I0(n43682), .I1(n43676), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n38680));
    defparam i31834_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1285 (.I0(n35638), .I1(n31482), .I2(n35599), 
            .I3(n16246), .O(n14_adj_4446));
    defparam i6_4_lut_adj_1285.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1286 (.I0(n31474), .I1(n14_adj_4446), .I2(n10_adj_4311), 
            .I3(n35347), .O(n37080));
    defparam i7_4_lut_adj_1286.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i19_3_lut (.I0(\data_out_frame[20] [5]), 
            .I1(\data_out_frame[21] [5]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4447));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i6_3_lut (.I0(\data_out_frame[5] [5]), 
            .I1(\byte_transmit_counter[1] ), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n41099));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i6_3_lut.LUT_INIT = 16'ha3a3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i5_3_lut (.I0(\data_out_frame[6] [5]), 
            .I1(\data_out_frame[7] [5]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4448));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31846_4_lut (.I0(n19_adj_4447), .I1(\data_out_frame[22] [5]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n38692));
    defparam i31846_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31847_3_lut (.I0(n43802), .I1(n38692), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n38693));
    defparam i31847_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31830_4_lut (.I0(n5_adj_4448), .I1(\byte_transmit_counter[0] ), 
            .I2(n40522), .I3(n41099), .O(n38676));
    defparam i31830_4_lut.LUT_INIT = 16'haca0;
    SB_LUT4 i31832_4_lut (.I0(n38676), .I1(n38693), .I2(\byte_transmit_counter[4] ), 
            .I3(\byte_transmit_counter[3] ), .O(n38678));
    defparam i31832_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31831_3_lut (.I0(n43700), .I1(n43688), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n38677));
    defparam i31831_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i19_3_lut (.I0(\data_out_frame[20] [4]), 
            .I1(\data_out_frame[21] [4]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4449));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i6_4_lut (.I0(\data_out_frame[5] [4]), 
            .I1(\byte_transmit_counter[1] ), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n6_adj_4450));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i6_4_lut.LUT_INIT = 16'hac03;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i5_3_lut (.I0(\data_out_frame[6] [4]), 
            .I1(\data_out_frame[7] [4]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4451));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1287 (.I0(n25_adj_4433), .I1(\FRAME_MATCHER.state [28]), 
            .I2(n26_adj_4427), .I3(\FRAME_MATCHER.state [25]), .O(n24968));
    defparam i1_4_lut_adj_1287.LUT_INIT = 16'hfffe;
    SB_LUT4 i31843_4_lut (.I0(n19_adj_4449), .I1(\data_out_frame[22] [4]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n38689));
    defparam i31843_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i3_4_lut_adj_1288 (.I0(n36436), .I1(n35508), .I2(n35273), 
            .I3(Kp_23__N_1802), .O(n31474));
    defparam i3_4_lut_adj_1288.LUT_INIT = 16'h9669;
    SB_LUT4 i31844_3_lut (.I0(n43796), .I1(n38689), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n38690));
    defparam i31844_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31827_3_lut (.I0(n5_adj_4451), .I1(n6_adj_4450), .I2(n40522), 
            .I3(GND_net), .O(n38673));
    defparam i31827_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31829_4_lut (.I0(n38673), .I1(n38690), .I2(\byte_transmit_counter[4] ), 
            .I3(\byte_transmit_counter[3] ), .O(n38675));
    defparam i31829_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31828_3_lut (.I0(n43724), .I1(n43706), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n38674));
    defparam i31828_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1289 (.I0(n36539), .I1(n37597), .I2(GND_net), 
            .I3(GND_net), .O(n31457));
    defparam i1_2_lut_adj_1289.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1290 (.I0(n31528), .I1(\data_in_frame[20] [3]), 
            .I2(\data_in_frame[20] [2]), .I3(GND_net), .O(n35279));
    defparam i2_3_lut_adj_1290.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1291 (.I0(n16953), .I1(n35578), .I2(n35438), 
            .I3(n6_adj_4440), .O(n35164));   // verilog/coms.v(84[17:63])
    defparam i4_4_lut_adj_1291.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1292 (.I0(\data_in_frame[15] [5]), .I1(n35429), 
            .I2(n30529), .I3(n31457), .O(n10_adj_4439));
    defparam i4_4_lut_adj_1292.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1293 (.I0(n16115), .I1(n35164), .I2(\data_in_frame[6] [5]), 
            .I3(GND_net), .O(n31068));
    defparam i2_3_lut_adj_1293.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1294 (.I0(\data_in_frame[7] [0]), .I1(\data_in_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35472));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1294.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1295 (.I0(\data_in_frame[22] [4]), .I1(\data_in_frame[18] [0]), 
            .I2(n35279), .I3(n15460), .O(n35344));
    defparam i1_4_lut_adj_1295.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1296 (.I0(\data_in_frame[16] [6]), .I1(n30653), 
            .I2(GND_net), .I3(GND_net), .O(n35364));
    defparam i1_2_lut_adj_1296.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1297 (.I0(n16115), .I1(\data_in_frame[7] [6]), 
            .I2(\data_in_frame[10] [0]), .I3(GND_net), .O(n16812));
    defparam i1_2_lut_3_lut_adj_1297.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i19_3_lut (.I0(\data_out_frame[20] [3]), 
            .I1(\data_out_frame[21] [3]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4452));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i6_4_lut (.I0(\data_out_frame[5] [3]), 
            .I1(\byte_transmit_counter[1] ), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n6_adj_4453));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i6_4_lut.LUT_INIT = 16'haf03;
    SB_LUT4 i1_2_lut_adj_1298 (.I0(n15609), .I1(Kp_23__N_1768), .I2(GND_net), 
            .I3(GND_net), .O(n35176));
    defparam i1_2_lut_adj_1298.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i5_3_lut (.I0(\data_out_frame[6] [3]), 
            .I1(\data_out_frame[7] [3]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4454));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31840_4_lut (.I0(n19_adj_4452), .I1(\data_out_frame[22] [3]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n38686));
    defparam i31840_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31841_3_lut (.I0(n43790), .I1(n38686), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n38687));
    defparam i31841_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31824_3_lut (.I0(n5_adj_4454), .I1(n6_adj_4453), .I2(n40522), 
            .I3(GND_net), .O(n38670));
    defparam i31824_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut_adj_1299 (.I0(n31482), .I1(n30812), .I2(\data_in_frame[21] [7]), 
            .I3(n6_adj_4438), .O(Kp_23__N_1768));
    defparam i4_4_lut_adj_1299.LUT_INIT = 16'h6996;
    SB_LUT4 i31826_4_lut (.I0(n38670), .I1(n38687), .I2(\byte_transmit_counter[4] ), 
            .I3(\byte_transmit_counter[3] ), .O(n38672));
    defparam i31826_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31825_3_lut (.I0(n43736), .I1(n43730), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n38671));
    defparam i31825_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_4_lut_adj_1300 (.I0(n35511), .I1(Kp_23__N_1768), .I2(\data_in_frame[19] [4]), 
            .I3(\data_in_frame[22] [0]), .O(n15_adj_4455));
    defparam i6_4_lut_adj_1300.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1301 (.I0(\FRAME_MATCHER.state [10]), .I1(\FRAME_MATCHER.state [15]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4456));
    defparam i2_2_lut_adj_1301.LUT_INIT = 16'heeee;
    SB_LUT4 i8_4_lut_adj_1302 (.I0(n15_adj_4455), .I1(\data_in_frame[17] [4]), 
            .I2(n14_adj_4437), .I3(\data_in_frame[17] [5]), .O(n35157));
    defparam i8_4_lut_adj_1302.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1303 (.I0(\data_in_frame[22] [2]), .I1(\data_in_frame[22] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16659));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_adj_1303.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36845 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [5]), .I2(\data_out_frame[15] [5]), 
            .I3(\byte_transmit_counter[1] ), .O(n43685));
    defparam byte_transmit_counter_0__bdd_4_lut_36845.LUT_INIT = 16'he4aa;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i19_3_lut (.I0(\data_out_frame[20] [2]), 
            .I1(\data_out_frame[21] [2]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4457));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_4_lut_adj_1304 (.I0(\data_in_frame[22] [4]), .I1(\data_in_frame[22] [3]), 
            .I2(n16659), .I3(\data_in_frame[22] [5]), .O(n35599));
    defparam i3_4_lut_adj_1304.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i6_4_lut (.I0(\data_out_frame[5] [2]), 
            .I1(\byte_transmit_counter[0] ), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[1] ), .O(n6_adj_4458));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i6_4_lut.LUT_INIT = 16'hb0b3;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i5_3_lut (.I0(\data_out_frame[6] [2]), 
            .I1(\data_out_frame[7] [2]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4459));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31837_4_lut (.I0(n19_adj_4457), .I1(\data_out_frame[22] [2]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n38683));
    defparam i31837_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31838_3_lut (.I0(n43778), .I1(n38683), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n38684));
    defparam i31838_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31821_3_lut (.I0(n5_adj_4459), .I1(n6_adj_4458), .I2(n40522), 
            .I3(GND_net), .O(n38667));
    defparam i31821_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31823_4_lut (.I0(n38667), .I1(n38684), .I2(\byte_transmit_counter[4] ), 
            .I3(\byte_transmit_counter[3] ), .O(n38669));
    defparam i31823_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31822_3_lut (.I0(n43748), .I1(n43742), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n38668));
    defparam i31822_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n43685_bdd_4_lut (.I0(n43685), .I1(\data_out_frame[13] [5]), 
            .I2(\data_out_frame[12] [5]), .I3(\byte_transmit_counter[1] ), 
            .O(n43688));
    defparam n43685_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i6_4_lut_adj_1305 (.I0(\FRAME_MATCHER.state [8]), .I1(\FRAME_MATCHER.state [12]), 
            .I2(\FRAME_MATCHER.state [9]), .I3(\FRAME_MATCHER.state [14]), 
            .O(n14_adj_4460));
    defparam i6_4_lut_adj_1305.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1306 (.I0(\data_in_frame[19] [5]), .I1(n35173), 
            .I2(\data_in_frame[17] [3]), .I3(n37297), .O(n30812));
    defparam i3_4_lut_adj_1306.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i19_3_lut (.I0(\data_out_frame[20] [1]), 
            .I1(\data_out_frame[21] [1]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n19_adj_4461));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_adj_1307 (.I0(n36306), .I1(n31610), .I2(\data_in_frame[16] [4]), 
            .I3(GND_net), .O(n30721));
    defparam i2_3_lut_adj_1307.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i6_3_lut (.I0(\data_out_frame[5] [1]), 
            .I1(\byte_transmit_counter[0] ), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n6_adj_4462));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i6_3_lut.LUT_INIT = 16'hbcbc;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i5_3_lut (.I0(\data_out_frame[6] [1]), 
            .I1(\data_out_frame[7] [1]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n5_adj_4463));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31810_4_lut (.I0(n19_adj_4461), .I1(\data_out_frame[22] [1]), 
            .I2(\byte_transmit_counter[1] ), .I3(\byte_transmit_counter[0] ), 
            .O(n38656));
    defparam i31810_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i31811_3_lut (.I0(n43718), .I1(n38656), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n38657));
    defparam i31811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36836 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [6]), .I2(\data_out_frame[11] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n43679));
    defparam byte_transmit_counter_0__bdd_4_lut_36836.LUT_INIT = 16'he4aa;
    SB_LUT4 i31818_3_lut (.I0(n5_adj_4463), .I1(n6_adj_4462), .I2(n40522), 
            .I3(GND_net), .O(n38664));
    defparam i31818_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i31820_4_lut (.I0(n38664), .I1(n38657), .I2(\byte_transmit_counter[4] ), 
            .I3(\byte_transmit_counter[3] ), .O(n38666));
    defparam i31820_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_adj_1308 (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[20] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35546));
    defparam i1_2_lut_adj_1308.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1309 (.I0(\data_in_frame[20] [7]), .I1(n35602), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4464));
    defparam i2_2_lut_adj_1309.LUT_INIT = 16'h6666;
    SB_LUT4 i31819_3_lut (.I0(n43760), .I1(n43754), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n38665));
    defparam i31819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_4_lut_adj_1310 (.I0(n16202), .I1(n7_adj_4436), .I2(\data_in_frame[20] [2]), 
            .I3(n8_adj_4464), .O(n35273));
    defparam i5_4_lut_adj_1310.LUT_INIT = 16'h6996;
    SB_LUT4 n43679_bdd_4_lut (.I0(n43679), .I1(\data_out_frame[9] [6]), 
            .I2(\data_out_frame[8] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n43682));
    defparam n43679_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1311 (.I0(\data_in_frame[22] [7]), .I1(\data_in_frame[22] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n16246));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_adj_1311.LUT_INIT = 16'h6666;
    SB_LUT4 i13204_3_lut_4_lut (.I0(n8_adj_4391), .I1(n34998), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n17943));
    defparam i13204_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1312 (.I0(\data_in_frame[21] [4]), .I1(\data_in_frame[21] [1]), 
            .I2(\data_in_frame[21] [3]), .I3(\data_in_frame[21] [2]), .O(n35218));   // verilog/coms.v(84[17:63])
    defparam i1_4_lut_adj_1312.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1313 (.I0(n35472), .I1(n35590), .I2(\data_in_frame[9] [1]), 
            .I3(n35164), .O(n12_adj_4465));   // verilog/coms.v(73[16:43])
    defparam i5_4_lut_adj_1313.LUT_INIT = 16'h6996;
    SB_LUT4 i13250_3_lut_4_lut (.I0(n8_adj_4320), .I1(n34998), .I2(rx_data[7]), 
            .I3(\data_in_frame[6][7] ), .O(n17989));
    defparam i13250_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_adj_1314 (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[18] [7]), 
            .I2(\data_in_frame[17] [0]), .I3(GND_net), .O(n35037));   // verilog/coms.v(75[16:43])
    defparam i1_3_lut_adj_1314.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1315 (.I0(\data_in_frame[19] [1]), .I1(n35037), 
            .I2(\data_in_frame[19] [3]), .I3(GND_net), .O(n35407));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1315.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1316 (.I0(\data_in_frame[18] [0]), .I1(n30588), 
            .I2(GND_net), .I3(GND_net), .O(n35638));
    defparam i1_2_lut_adj_1316.LUT_INIT = 16'h6666;
    SB_LUT4 i13243_3_lut_4_lut (.I0(n8_adj_4320), .I1(n34998), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n17982));
    defparam i13243_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_110_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(GND_net), .O(n8_adj_4407));   // verilog/coms.v(154[7:23])
    defparam equal_110_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i13244_3_lut_4_lut (.I0(n8_adj_4320), .I1(n34998), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n17983));
    defparam i13244_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1317 (.I0(\data_in_frame[15] [0]), .I1(n30512), 
            .I2(n8_adj_4466), .I3(\data_in_frame[14] [6]), .O(n35511));
    defparam i1_4_lut_adj_1317.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1318 (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[19] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35410));
    defparam i1_2_lut_adj_1318.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1319 (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[19] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35515));
    defparam i1_2_lut_adj_1319.LUT_INIT = 16'h6666;
    SB_LUT4 i13245_3_lut_4_lut (.I0(n8_adj_4320), .I1(n34998), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n17984));
    defparam i13245_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1320 (.I0(\data_in_frame[12] [4]), .I1(\data_in_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n16486));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_adj_1320.LUT_INIT = 16'h6666;
    SB_LUT4 i13246_3_lut_4_lut (.I0(n8_adj_4320), .I1(n34998), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n17985));
    defparam i13246_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i41_4_lut (.I0(\data_in_frame[10] [3]), .I1(n35543), .I2(n35626), 
            .I3(n35357), .O(n98));
    defparam i41_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i39_4_lut (.I0(n30730), .I1(n35167), .I2(\data_in_frame[13] [4]), 
            .I3(n35388), .O(n96));
    defparam i39_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i40_4_lut (.I0(\data_in_frame[10] [4]), .I1(n35294), .I2(n35552), 
            .I3(Kp_23__N_805), .O(n97));
    defparam i40_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i19964_1_lut (.I0(n24684), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n2058));
    defparam i19964_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i13247_3_lut_4_lut (.I0(n8_adj_4320), .I1(n34998), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n17986));
    defparam i13247_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i38_4_lut (.I0(n35555), .I1(n16486), .I2(n35135), .I3(\data_in_frame[12] [3]), 
            .O(n95));
    defparam i38_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13248_3_lut_4_lut (.I0(n8_adj_4320), .I1(n34998), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n17987));
    defparam i13248_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i33_4_lut (.I0(\data_in_frame[16] [6]), .I1(n35309), .I2(n36306), 
            .I3(n31476), .O(n90));
    defparam i33_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1321 (.I0(\FRAME_MATCHER.state [31]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34323));
    defparam i1_2_lut_adj_1321.LUT_INIT = 16'h8888;
    SB_LUT4 i31_4_lut (.I0(n35515), .I1(n16835), .I2(n35188), .I3(n35575), 
            .O(n88));
    defparam i31_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1322 (.I0(\FRAME_MATCHER.state [28]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34379));
    defparam i1_2_lut_adj_1322.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1323 (.I0(\FRAME_MATCHER.state [27]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34341));
    defparam i1_2_lut_adj_1323.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1324 (.I0(\FRAME_MATCHER.state [26]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34337));
    defparam i1_2_lut_adj_1324.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_3_lut_adj_1325 (.I0(n30671), .I1(n16876), .I2(n17011), 
            .I3(GND_net), .O(n6_adj_4408));
    defparam i1_2_lut_3_lut_adj_1325.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1326 (.I0(\FRAME_MATCHER.state [24]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34345));
    defparam i1_2_lut_adj_1326.LUT_INIT = 16'h8888;
    SB_LUT4 i32_4_lut (.I0(n35407), .I1(\data_in_frame[17] [4]), .I2(n35341), 
            .I3(\data_in_frame[19] [5]), .O(n89));
    defparam i32_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut (.I0(\data_in_frame[19] [6]), .I1(n35354), .I2(\data_in_frame[20] [1]), 
            .I3(\data_in_frame[17] [6]), .O(n87));
    defparam i30_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1327 (.I0(\FRAME_MATCHER.state [23]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34347));
    defparam i1_2_lut_adj_1327.LUT_INIT = 16'h8888;
    SB_LUT4 i37_4_lut (.I0(\data_in_frame[13] [5]), .I1(n31457), .I2(n35463), 
            .I3(\data_in_frame[13] [3]), .O(n94));
    defparam i37_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1328 (.I0(\FRAME_MATCHER.state [22]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34349));
    defparam i1_2_lut_adj_1328.LUT_INIT = 16'h8888;
    SB_LUT4 i13249_3_lut_4_lut (.I0(n8_adj_4320), .I1(n34998), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n17988));
    defparam i13249_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i35_4_lut (.I0(n35511), .I1(n35303), .I2(n35315), .I3(\data_in_frame[14] [7]), 
            .O(n92));
    defparam i35_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i36_4_lut (.I0(n30592), .I1(n16272), .I2(n37527), .I3(\data_in_frame[13] [2]), 
            .O(n93));
    defparam i36_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1329 (.I0(\FRAME_MATCHER.state [20]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34381));
    defparam i1_2_lut_adj_1329.LUT_INIT = 16'h8888;
    SB_LUT4 i13205_3_lut_4_lut (.I0(n8_adj_4391), .I1(n34998), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n17944));
    defparam i13205_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i34_4_lut (.I0(n35367), .I1(\data_in_frame[13] [6]), .I2(n35147), 
            .I3(n37297), .O(n91));
    defparam i34_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1330 (.I0(\FRAME_MATCHER.state[1] ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n15963), .I3(n15958), .O(n15960));   // verilog/coms.v(151[5:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1330.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1331 (.I0(\FRAME_MATCHER.state[1] ), 
            .I1(\FRAME_MATCHER.state[3] ), .I2(n15963), .I3(n24190), .O(n15957));   // verilog/coms.v(151[5:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1331.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_adj_1332 (.I0(\FRAME_MATCHER.state [16]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34383));
    defparam i1_2_lut_adj_1332.LUT_INIT = 16'h8888;
    SB_LUT4 i42_4_lut (.I0(n35249), .I1(\data_in_frame[11] [1]), .I2(\data_in_frame[10] [2]), 
            .I3(\data_in_frame[10] [1]), .O(n99));
    defparam i42_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1333 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [3]), 
            .I2(n15845), .I3(\FRAME_MATCHER.i [2]), .O(n4_adj_4400));
    defparam i1_2_lut_4_lut_adj_1333.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1334 (.I0(\FRAME_MATCHER.state [15]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34385));
    defparam i1_2_lut_adj_1334.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1335 (.I0(\FRAME_MATCHER.state [14]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34351));
    defparam i1_2_lut_adj_1335.LUT_INIT = 16'h8888;
    SB_LUT4 i53_4_lut (.I0(n95), .I1(n97), .I2(n96), .I3(n98), .O(n110));
    defparam i53_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i51_4_lut (.I0(n87), .I1(n89), .I2(n88), .I3(n90), .O(n108));
    defparam i51_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1336 (.I0(\FRAME_MATCHER.state [13]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34387));
    defparam i1_2_lut_adj_1336.LUT_INIT = 16'h8888;
    SB_LUT4 i52_4_lut (.I0(n91), .I1(n93), .I2(n92), .I3(n94), .O(n109));
    defparam i52_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1337 (.I0(\FRAME_MATCHER.state [12]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34339));
    defparam i1_2_lut_adj_1337.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1338 (.I0(\FRAME_MATCHER.state [11]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34389));
    defparam i1_2_lut_adj_1338.LUT_INIT = 16'h8888;
    SB_LUT4 i50_4_lut (.I0(n99), .I1(\data_in_frame[10] [0]), .I2(n86), 
            .I3(\data_in_frame[18] [2]), .O(n107));
    defparam i50_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i13206_3_lut_4_lut (.I0(n8_adj_4391), .I1(n34998), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n17945));
    defparam i13206_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1339 (.I0(\FRAME_MATCHER.state [10]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34401));
    defparam i1_2_lut_adj_1339.LUT_INIT = 16'h8888;
    SB_LUT4 i56_4_lut (.I0(n107), .I1(n109), .I2(n108), .I3(n110), .O(n35602));
    defparam i56_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20245_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), .I1(\byte_transmit_counter[1] ), 
            .I2(\byte_transmit_counter[4] ), .I3(\byte_transmit_counter[3] ), 
            .O(n24966));
    defparam i20245_3_lut_4_lut.LUT_INIT = 16'hf080;
    SB_LUT4 i1_2_lut_adj_1340 (.I0(\FRAME_MATCHER.state [9]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34335));
    defparam i1_2_lut_adj_1340.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1341 (.I0(\FRAME_MATCHER.state [8]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34391));
    defparam i1_2_lut_adj_1341.LUT_INIT = 16'h8888;
    SB_LUT4 i13339_3_lut_4_lut (.I0(n10_adj_4425), .I1(n34995), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n18078));
    defparam i13339_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1342 (.I0(\FRAME_MATCHER.state [7]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34393));
    defparam i1_2_lut_adj_1342.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1343 (.I0(\FRAME_MATCHER.state [6]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34395));
    defparam i1_2_lut_adj_1343.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1344 (.I0(\FRAME_MATCHER.state [5]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34397));
    defparam i1_2_lut_adj_1344.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_1345 (.I0(n13144), .I1(n13181), .I2(n15958), 
            .I3(n24190), .O(n9_adj_4401));
    defparam i1_4_lut_adj_1345.LUT_INIT = 16'hce0a;
    SB_LUT4 i1_2_lut_adj_1346 (.I0(\FRAME_MATCHER.state [4]), .I1(n12_adj_4402), 
            .I2(GND_net), .I3(GND_net), .O(n34331));
    defparam i1_2_lut_adj_1346.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_1347 (.I0(n31476), .I1(\data_in_frame[19] [7]), 
            .I2(\data_in_frame[17] [5]), .I3(n16272), .O(n31482));
    defparam i2_3_lut_4_lut_adj_1347.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1348 (.I0(n2957), .I1(n10389), .I2(GND_net), 
            .I3(GND_net), .O(n13181));   // verilog/coms.v(222[6] 224[9])
    defparam i1_2_lut_adj_1348.LUT_INIT = 16'h4444;
    SB_LUT4 i1_2_lut_adj_1349 (.I0(n788), .I1(n10389), .I2(GND_net), .I3(GND_net), 
            .O(n13144));   // verilog/coms.v(157[6] 159[9])
    defparam i1_2_lut_adj_1349.LUT_INIT = 16'h4444;
    SB_LUT4 i1_3_lut_adj_1350 (.I0(n15994), .I1(n3894), .I2(n10389), .I3(GND_net), 
            .O(n67));   // verilog/coms.v(246[5:25])
    defparam i1_3_lut_adj_1350.LUT_INIT = 16'h1010;
    SB_LUT4 i55_2_lut (.I0(n10389), .I1(n2774), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i13207_3_lut_4_lut (.I0(n8_adj_4391), .I1(n34998), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n17946));
    defparam i13207_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i80_4_lut (.I0(n46), .I1(\FRAME_MATCHER.state[3] ), .I2(n15_adj_4390), 
            .I3(n70), .O(n65));   // verilog/coms.v(114[11:12])
    defparam i80_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i81_4_lut (.I0(n65), .I1(\FRAME_MATCHER.state [2]), .I2(n43_adj_4416), 
            .I3(\FRAME_MATCHER.state_31__N_2725 [3]), .O(n10_adj_4385));   // verilog/coms.v(114[11:12])
    defparam i81_4_lut.LUT_INIT = 16'habaa;
    SB_LUT4 i13208_3_lut_4_lut (.I0(n8_adj_4391), .I1(n34998), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n17947));
    defparam i13208_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13340_3_lut_4_lut (.I0(n10_adj_4425), .I1(n34995), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n18079));
    defparam i13340_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i28992_2_lut (.I0(n15994), .I1(n3894), .I2(GND_net), .I3(GND_net), 
            .O(n35746));
    defparam i28992_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1351 (.I0(n30730), .I1(n30622), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4467));
    defparam i1_2_lut_adj_1351.LUT_INIT = 16'h6666;
    SB_LUT4 i13341_3_lut_4_lut (.I0(n10_adj_4425), .I1(n34995), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n18080));
    defparam i13341_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i19462_2_lut (.I0(n23[1]), .I1(n63), .I2(GND_net), .I3(GND_net), 
            .O(\FRAME_MATCHER.state_31__N_2661 [1]));   // verilog/coms.v(142[4] 144[7])
    defparam i19462_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 select_368_Select_1_i5_4_lut (.I0(n63), .I1(n15957), .I2(n2957), 
            .I3(n23[1]), .O(n5_adj_4468));
    defparam select_368_Select_1_i5_4_lut.LUT_INIT = 16'h3331;
    SB_LUT4 i4_4_lut_adj_1352 (.I0(\data_in_frame[12] [3]), .I1(\data_in_frame[12] [4]), 
            .I2(\data_in_frame[14] [5]), .I3(n6_adj_4467), .O(n37403));
    defparam i4_4_lut_adj_1352.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1353 (.I0(n63_adj_3), .I1(n23[1]), .I2(n15960), 
            .I3(n9015), .O(n5_adj_4469));
    defparam i1_4_lut_adj_1353.LUT_INIT = 16'h5d5f;
    SB_LUT4 i3_4_lut_adj_1354 (.I0(n5_adj_4469), .I1(\FRAME_MATCHER.state_31__N_2661 [1]), 
            .I2(n5_adj_4468), .I3(n35746), .O(n44032));
    defparam i3_4_lut_adj_1354.LUT_INIT = 16'hfafe;
    SB_LUT4 i13342_3_lut_4_lut (.I0(n10_adj_4425), .I1(n34995), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n18081));
    defparam i13342_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1355 (.I0(n37403), .I1(\data_in_frame[16] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35315));
    defparam i1_2_lut_adj_1355.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1356 (.I0(\data_in_frame[12] [4]), .I1(n30512), 
            .I2(\data_in_frame[14] [6]), .I3(\data_in_frame[12] [5]), .O(n31470));
    defparam i3_4_lut_adj_1356.LUT_INIT = 16'h6996;
    SB_LUT4 i13209_3_lut_4_lut (.I0(n8_adj_4391), .I1(n34998), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n17948));
    defparam i13209_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13343_3_lut_4_lut (.I0(n10_adj_4425), .I1(n34995), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n18082));
    defparam i13343_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1357 (.I0(n35129), .I1(\data_in_frame[10] [3]), 
            .I2(n16642), .I3(GND_net), .O(n30730));
    defparam i2_3_lut_adj_1357.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1358 (.I0(\data_in_frame[14] [7]), .I1(n30730), 
            .I2(GND_net), .I3(GND_net), .O(n35336));
    defparam i1_2_lut_adj_1358.LUT_INIT = 16'h6666;
    SB_LUT4 i36779_3_lut (.I0(n15963), .I1(n15886), .I2(n15861), .I3(GND_net), 
            .O(n37152));
    defparam i36779_3_lut.LUT_INIT = 16'h0101;
    SB_LUT4 i5_4_lut_adj_1359 (.I0(\data_in_frame[12] [5]), .I1(n35617), 
            .I2(n35212), .I3(n35336), .O(n12_adj_4470));
    defparam i5_4_lut_adj_1359.LUT_INIT = 16'h6996;
    SB_LUT4 i13344_3_lut_4_lut (.I0(n10_adj_4425), .I1(n34995), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n18083));
    defparam i13344_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i6_4_lut_adj_1360 (.I0(\data_in_frame[13] [0]), .I1(n12_adj_4470), 
            .I2(\data_in_frame[15] [1]), .I3(n35533), .O(n37297));
    defparam i6_4_lut_adj_1360.LUT_INIT = 16'h6996;
    SB_LUT4 i36760_4_lut (.I0(n15861), .I1(n4498), .I2(n5_adj_4435), .I3(n6_adj_4314), 
            .O(n34927));
    defparam i36760_4_lut.LUT_INIT = 16'h1115;
    SB_LUT4 i13345_3_lut_4_lut (.I0(n10_adj_4425), .I1(n34995), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n18084));
    defparam i13345_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13346_3_lut_4_lut (.I0(n10_adj_4425), .I1(n34995), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n18085));
    defparam i13346_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1361 (.I0(\FRAME_MATCHER.i [0]), .I1(n7_adj_4404), 
            .I2(n161), .I3(n24684), .O(n34995));   // verilog/coms.v(154[7:23])
    defparam i1_2_lut_3_lut_4_lut_adj_1361.LUT_INIT = 16'hffef;
    SB_LUT4 i1_2_lut_adj_1362 (.I0(\data_in_frame[17] [2]), .I1(n37297), 
            .I2(GND_net), .I3(GND_net), .O(n31460));
    defparam i1_2_lut_adj_1362.LUT_INIT = 16'h9999;
    SB_LUT4 i3_4_lut_adj_1363 (.I0(\data_out_frame[20] [3]), .I1(n35285), 
            .I2(\data_out_frame[20] [4]), .I3(n35525), .O(n36345));
    defparam i3_4_lut_adj_1363.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1364 (.I0(n31017), .I1(n35382), .I2(GND_net), 
            .I3(GND_net), .O(n35383));
    defparam i1_2_lut_adj_1364.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1365 (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[18] [1]), 
            .I2(n35318), .I3(n6_adj_4434), .O(n36260));
    defparam i4_4_lut_adj_1365.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1366 (.I0(n36368), .I1(n35351), .I2(\data_out_frame[20] [1]), 
            .I3(GND_net), .O(n36143));
    defparam i2_3_lut_adj_1366.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1367 (.I0(n14129), .I1(\data_out_frame[19] [7]), 
            .I2(n16020), .I3(\data_out_frame[17] [5]), .O(n10_adj_4471));
    defparam i4_4_lut_adj_1367.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1368 (.I0(\data_out_frame[13] [2]), .I1(\data_out_frame[13] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16020));   // verilog/coms.v(84[17:63])
    defparam i1_2_lut_adj_1368.LUT_INIT = 16'h6666;
    SB_LUT4 i13330_3_lut_4_lut (.I0(n8_adj_4399), .I1(n35006), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n18069));
    defparam i13330_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1369 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4472));
    defparam i1_2_lut_adj_1369.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1370 (.I0(\data_out_frame[13] [3]), .I1(n7_adj_4472), 
            .I2(n30582), .I3(n8_adj_4313), .O(n16566));
    defparam i5_4_lut_adj_1370.LUT_INIT = 16'h6996;
    SB_LUT4 i13210_3_lut_4_lut (.I0(n8_adj_4391), .I1(n34998), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n17949));
    defparam i13210_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7_4_lut_adj_1371 (.I0(\FRAME_MATCHER.state [13]), .I1(n14_adj_4460), 
            .I2(n10_adj_4456), .I3(\FRAME_MATCHER.state [11]), .O(n24910));
    defparam i7_4_lut_adj_1371.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1372 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35549));
    defparam i1_2_lut_adj_1372.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1373 (.I0(\data_in_frame[5] [6]), .I1(n35518), 
            .I2(n35629), .I3(n35394), .O(n22_adj_4473));
    defparam i9_4_lut_adj_1373.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut_adj_1374 (.I0(n31068), .I1(\data_in_frame[10] [1]), 
            .I2(n35472), .I3(GND_net), .O(n20_adj_4474));
    defparam i7_3_lut_adj_1374.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut_adj_1375 (.I0(Kp_23__N_949), .I1(n22_adj_4473), .I2(n16_adj_4429), 
            .I3(\data_in_frame[8] [3]), .O(n24_adj_4475));
    defparam i11_4_lut_adj_1375.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1376 (.I0(n35122), .I1(n24_adj_4475), .I2(n20_adj_4474), 
            .I3(n16782), .O(n30622));
    defparam i12_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i12853_3_lut_4_lut (.I0(n8_adj_4399), .I1(n34998), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n17592));
    defparam i12853_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1377 (.I0(\data_in_frame[8] [1]), .I1(n16464), 
            .I2(n35091), .I3(\data_in_frame[7] [7]), .O(n35129));
    defparam i3_4_lut_adj_1377.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36831 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [6]), .I2(\data_out_frame[15] [6]), 
            .I3(\byte_transmit_counter[1] ), .O(n43673));
    defparam byte_transmit_counter_0__bdd_4_lut_36831.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_adj_1378 (.I0(\data_in_frame[10] [2]), .I1(n16386), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4476));
    defparam i1_2_lut_adj_1378.LUT_INIT = 16'h6666;
    SB_LUT4 n43673_bdd_4_lut (.I0(n43673), .I1(\data_out_frame[13] [6]), 
            .I2(\data_out_frame[12] [6]), .I3(\byte_transmit_counter[1] ), 
            .O(n43676));
    defparam n43673_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1379 (.I0(n16566), .I1(n30667), .I2(GND_net), 
            .I3(GND_net), .O(n35521));
    defparam i1_2_lut_adj_1379.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1380 (.I0(n35129), .I1(n6_adj_4296), .I2(n35454), 
            .I3(n6_adj_4476), .O(n35185));
    defparam i4_4_lut_adj_1380.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1381 (.I0(\data_in_frame[12] [3]), .I1(n35502), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4477));
    defparam i1_2_lut_adj_1381.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1382 (.I0(\data_out_frame[18] [4]), .I1(n30516), 
            .I2(\data_out_frame[18] [3]), .I3(n31552), .O(n31518));
    defparam i3_4_lut_adj_1382.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1383 (.I0(n31518), .I1(n35285), .I2(GND_net), 
            .I3(GND_net), .O(n30681));
    defparam i1_2_lut_adj_1383.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1384 (.I0(\data_in_frame[14] [4]), .I1(\data_in_frame[12] [2]), 
            .I2(n35185), .I3(n6_adj_4477), .O(n30653));
    defparam i4_4_lut_adj_1384.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1385 (.I0(n30653), .I1(\data_in_frame[16] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n35303));
    defparam i1_2_lut_adj_1385.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1386 (.I0(n16184), .I1(n35614), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4478));
    defparam i1_2_lut_adj_1386.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1387 (.I0(\data_out_frame[15] [2]), .I1(n31504), 
            .I2(n35530), .I3(n6_adj_4478), .O(n35351));
    defparam i4_4_lut_adj_1387.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1388 (.I0(n31017), .I1(n36368), .I2(n30681), 
            .I3(n6_adj_4479), .O(n35271));
    defparam i4_4_lut_adj_1388.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1389 (.I0(n35271), .I1(n35351), .I2(GND_net), 
            .I3(GND_net), .O(n35353));
    defparam i1_2_lut_adj_1389.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1390 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35382));
    defparam i1_2_lut_adj_1390.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1391 (.I0(\data_out_frame[20] [5]), .I1(\data_out_frame[20] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35070));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1391.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1392 (.I0(\data_out_frame[15] [3]), .I1(n31140), 
            .I2(GND_net), .I3(GND_net), .O(n31595));
    defparam i1_2_lut_adj_1392.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1393 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [6]), 
            .I2(n35081), .I3(n31595), .O(n35614));
    defparam i3_4_lut_adj_1393.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1394 (.I0(\data_out_frame[18] [3]), .I1(\data_out_frame[18] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16163));
    defparam i1_2_lut_adj_1394.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1395 (.I0(n35033), .I1(\data_out_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n18_adj_4480));
    defparam i1_2_lut_adj_1395.LUT_INIT = 16'h6666;
    SB_LUT4 i13_4_lut_adj_1396 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[15] [7]), 
            .I2(n17033), .I3(n18_adj_4480), .O(n30_adj_4481));
    defparam i13_4_lut_adj_1396.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1397 (.I0(\data_out_frame[5] [6]), .I1(\data_out_frame[16] [1]), 
            .I2(\data_out_frame[11] [7]), .I3(n35505), .O(n28_adj_4482));
    defparam i11_4_lut_adj_1397.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1398 (.I0(n35288), .I1(n17080), .I2(n35141), 
            .I3(\data_out_frame[13] [5]), .O(n29_adj_4483));
    defparam i12_4_lut_adj_1398.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1399 (.I0(n35397), .I1(n35587), .I2(\data_out_frame[13] [7]), 
            .I3(n35262), .O(n27_adj_4484));
    defparam i10_4_lut_adj_1399.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1400 (.I0(n27_adj_4484), .I1(n29_adj_4483), .I2(n28_adj_4482), 
            .I3(n30_adj_4481), .O(n30516));
    defparam i16_4_lut_adj_1400.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1401 (.I0(n30622), .I1(n35549), .I2(n35370), 
            .I3(n16812), .O(n12_adj_4485));
    defparam i5_4_lut_adj_1401.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1402 (.I0(\data_in_frame[14] [3]), .I1(n35502), 
            .I2(n12_adj_4485), .I3(n8_adj_4312), .O(n31610));
    defparam i1_4_lut_adj_1402.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1403 (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[20] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4486));   // verilog/coms.v(69[16:27])
    defparam i1_2_lut_adj_1403.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1404 (.I0(\data_in_frame[18] [5]), .I1(n17023), 
            .I2(n31558), .I3(n6_adj_4486), .O(n35276));   // verilog/coms.v(69[16:27])
    defparam i4_4_lut_adj_1404.LUT_INIT = 16'h9669;
    SB_LUT4 i13196_3_lut_4_lut (.I0(n8_adj_4399), .I1(n34998), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n17935));
    defparam i13196_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1405 (.I0(n24910), .I1(n24968), .I2(n24686), 
            .I3(GND_net), .O(n15963));   // verilog/coms.v(151[5:27])
    defparam i2_3_lut_adj_1405.LUT_INIT = 16'hfefe;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36826 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[10] [7]), .I2(\data_out_frame[11] [7]), 
            .I3(\byte_transmit_counter[1] ), .O(n43667));
    defparam byte_transmit_counter_0__bdd_4_lut_36826.LUT_INIT = 16'he4aa;
    SB_LUT4 n43667_bdd_4_lut (.I0(n43667), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[8] [7]), .I3(\byte_transmit_counter[1] ), 
            .O(n43670));
    defparam n43667_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1406 (.I0(\FRAME_MATCHER.state[3] ), .I1(n15963), 
            .I2(GND_net), .I3(GND_net), .O(n15722));   // verilog/coms.v(151[5:27])
    defparam i1_2_lut_adj_1406.LUT_INIT = 16'heeee;
    SB_LUT4 select_340_Select_31_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [31]), .O(n3_adj_4384));
    defparam select_340_Select_31_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i13197_3_lut_4_lut (.I0(n8_adj_4399), .I1(n34998), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n17936));
    defparam i13197_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1407 (.I0(n30807), .I1(n31530), .I2(GND_net), 
            .I3(GND_net), .O(n35309));
    defparam i1_2_lut_adj_1407.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_adj_1408 (.I0(n30669), .I1(\data_in_frame[7] [2]), 
            .I2(\data_in_frame[13] [6]), .I3(GND_net), .O(n9_adj_4393));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1408.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_1409 (.I0(n30545), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[11] [4]), .I3(GND_net), .O(n35376));
    defparam i2_3_lut_adj_1409.LUT_INIT = 16'h9696;
    SB_LUT4 i13198_3_lut_4_lut (.I0(n8_adj_4399), .I1(n34998), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n17937));
    defparam i13198_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_340_Select_30_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [30]), .O(n3_adj_4382));
    defparam select_340_Select_30_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_340_Select_29_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [29]), .O(n3_adj_4380));
    defparam select_340_Select_29_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36821 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[14] [7]), .I2(\data_out_frame[15] [7]), 
            .I3(\byte_transmit_counter[1] ), .O(n43661));
    defparam byte_transmit_counter_0__bdd_4_lut_36821.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1410 (.I0(n24684), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(n10_adj_4424), 
            .O(n34998));
    defparam i1_2_lut_3_lut_4_lut_adj_1410.LUT_INIT = 16'hfffb;
    SB_LUT4 i3_4_lut_adj_1411 (.I0(\data_out_frame[15] [5]), .I1(n30582), 
            .I2(n31510), .I3(n16029), .O(n16184));
    defparam i3_4_lut_adj_1411.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1412 (.I0(n16184), .I1(\data_out_frame[18] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n35524));
    defparam i1_2_lut_adj_1412.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1413 (.I0(\data_out_frame[13] [3]), .I1(\data_out_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n16029));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1413.LUT_INIT = 16'h6666;
    SB_LUT4 select_340_Select_28_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [28]), .O(n3_adj_4378));
    defparam select_340_Select_28_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i13199_3_lut_4_lut (.I0(n8_adj_4399), .I1(n34998), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n17938));
    defparam i13199_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_340_Select_27_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [27]), .O(n3_adj_4376));
    defparam select_340_Select_27_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i3_4_lut_adj_1414 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[6] [7]), 
            .I2(\data_out_frame[6] [4]), .I3(\data_out_frame[9] [0]), .O(n12_adj_4487));
    defparam i3_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1415 (.I0(n35478), .I1(\data_out_frame[9] [1]), 
            .I2(\data_out_frame[8] [4]), .I3(n35196), .O(n16_adj_4488));
    defparam i7_4_lut_adj_1415.LUT_INIT = 16'h6996;
    SB_LUT4 select_340_Select_26_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [26]), .O(n3_adj_4374));
    defparam select_340_Select_26_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i13200_3_lut_4_lut (.I0(n8_adj_4399), .I1(n34998), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n17939));
    defparam i13200_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i8_4_lut_adj_1416 (.I0(n35379), .I1(n16_adj_4488), .I2(n12_adj_4487), 
            .I3(\data_out_frame[11] [1]), .O(n31510));
    defparam i8_4_lut_adj_1416.LUT_INIT = 16'h6996;
    SB_LUT4 select_340_Select_25_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [25]), .O(n3_adj_4372));
    defparam select_340_Select_25_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 n43661_bdd_4_lut (.I0(n43661), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[12] [7]), .I3(\byte_transmit_counter[1] ), 
            .O(n43664));
    defparam n43661_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_adj_1417 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n35265));   // verilog/coms.v(84[17:70])
    defparam i1_2_lut_adj_1417.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1418 (.I0(\FRAME_MATCHER.state [2]), .I1(\FRAME_MATCHER.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n15958));   // verilog/coms.v(246[5:25])
    defparam i1_2_lut_adj_1418.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_1419 (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n35288));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1419.LUT_INIT = 16'h6666;
    SB_LUT4 select_340_Select_24_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [24]), .O(n3_adj_4370));
    defparam select_340_Select_24_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i13201_3_lut_4_lut (.I0(n8_adj_4399), .I1(n34998), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n17940));
    defparam i13201_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1420 (.I0(\data_out_frame[7] [0]), .I1(n16772), 
            .I2(GND_net), .I3(GND_net), .O(n35379));
    defparam i1_2_lut_adj_1420.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1421 (.I0(n30545), .I1(n7_adj_4430), .I2(n16949), 
            .I3(n8_adj_4431), .O(n31455));
    defparam i5_4_lut_adj_1421.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1422 (.I0(\data_out_frame[15] [6]), .I1(\data_out_frame[17] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35079));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_1422.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1423 (.I0(n31510), .I1(n35107), .I2(\data_out_frame[13] [3]), 
            .I3(GND_net), .O(n30667));
    defparam i2_3_lut_adj_1423.LUT_INIT = 16'h6969;
    SB_LUT4 select_340_Select_23_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [23]), .O(n3_adj_4368));
    defparam select_340_Select_23_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_340_Select_22_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [22]), .O(n3_adj_4366));
    defparam select_340_Select_22_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_340_Select_21_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [21]), .O(n3_adj_4364));
    defparam select_340_Select_21_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_340_Select_20_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [20]), .O(n3_adj_4362));
    defparam select_340_Select_20_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i6_4_lut_adj_1424 (.I0(n16876), .I1(n12_adj_4465), .I2(n35641), 
            .I3(n15568), .O(n31118));   // verilog/coms.v(73[16:43])
    defparam i6_4_lut_adj_1424.LUT_INIT = 16'h6996;
    SB_LUT4 select_340_Select_19_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [19]), .O(n3_adj_4360));
    defparam select_340_Select_19_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_340_Select_18_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [18]), .O(n3_adj_4358));
    defparam select_340_Select_18_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_340_Select_17_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [17]), .O(n3_adj_4356));
    defparam select_340_Select_17_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_340_Select_16_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [16]), .O(n3_adj_4354));
    defparam select_340_Select_16_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i13202_3_lut_4_lut (.I0(n8_adj_4399), .I1(n34998), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n17941));
    defparam i13202_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_340_Select_15_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [15]), .O(n3_adj_4352));
    defparam select_340_Select_15_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_adj_1425 (.I0(\data_in_frame[13] [3]), .I1(n31118), 
            .I2(GND_net), .I3(GND_net), .O(n35429));
    defparam i1_2_lut_adj_1425.LUT_INIT = 16'h6666;
    SB_LUT4 select_340_Select_14_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [14]), .O(n3_adj_4350));
    defparam select_340_Select_14_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i13323_3_lut_4_lut (.I0(n8_adj_4399), .I1(n35006), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n18062));
    defparam i13323_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_340_Select_13_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [13]), .O(n3_adj_4348));
    defparam select_340_Select_13_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 select_340_Select_12_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [12]), .O(n3_adj_4346));
    defparam select_340_Select_12_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i3_3_lut_4_lut_adj_1426 (.I0(\data_in_frame[10] [5]), .I1(n35167), 
            .I2(n35336), .I3(n16486), .O(n8_adj_4466));   // verilog/coms.v(74[16:43])
    defparam i3_3_lut_4_lut_adj_1426.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1427 (.I0(n35060), .I1(\data_out_frame[13] [7]), 
            .I2(\data_out_frame[9] [4]), .I3(\data_out_frame[13] [6]), .O(n36548));   // verilog/coms.v(84[17:28])
    defparam i3_4_lut_adj_1427.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1428 (.I0(n30667), .I1(n35079), .I2(\data_out_frame[17] [6]), 
            .I3(n31455), .O(n31140));   // verilog/coms.v(77[16:27])
    defparam i3_4_lut_adj_1428.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1429 (.I0(\data_in_frame[10] [6]), .I1(\data_in_frame[11] [0]), 
            .I2(n16883), .I3(\data_in_frame[11] [2]), .O(n35357));
    defparam i3_4_lut_adj_1429.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1430 (.I0(n35404), .I1(n16029), .I2(n30558), 
            .I3(n35647), .O(n52));
    defparam i18_4_lut_adj_1430.LUT_INIT = 16'h6996;
    SB_LUT4 i25_4_lut_adj_1431 (.I0(n35475), .I1(n35484), .I2(\data_out_frame[14] [5]), 
            .I3(n35426), .O(n59));
    defparam i25_4_lut_adj_1431.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1432 (.I0(\data_out_frame[13] [3]), .I1(n35524), 
            .I2(n35608), .I3(n31504), .O(n40_adj_4489));
    defparam i16_4_lut_adj_1432.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1433 (.I0(n35448), .I1(\data_out_frame[19] [4]), 
            .I2(\data_out_frame[17] [7]), .I3(n35527), .O(n38));
    defparam i14_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1434 (.I0(n35236), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[17] [5]), .I3(n31478), .O(n39_adj_4490));
    defparam i15_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1435 (.I0(n31478), .I1(n35614), .I2(n31510), 
            .I3(\data_out_frame[17] [4]), .O(n37));
    defparam i13_4_lut_adj_1435.LUT_INIT = 16'h9669;
    SB_LUT4 i22_4_lut (.I0(n35400), .I1(n35230), .I2(n35306), .I3(n35064), 
            .O(n56));
    defparam i22_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(n35376), .I1(\data_out_frame[15] [1]), .I2(n35107), 
            .I3(\data_out_frame[15] [2]), .O(n54));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i21_4_lut (.I0(n35054), .I1(\data_out_frame[9] [1]), .I2(\data_out_frame[12] [2]), 
            .I3(n35460), .O(n55));
    defparam i21_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i19_4_lut_adj_1436 (.I0(n35265), .I1(\data_out_frame[16] [6]), 
            .I2(n14107), .I3(n35587), .O(n53));
    defparam i19_4_lut_adj_1436.LUT_INIT = 16'h6996;
    SB_LUT4 i24_4_lut_adj_1437 (.I0(n30516), .I1(n35565), .I2(\data_out_frame[15] [3]), 
            .I3(n16214), .O(n58));
    defparam i24_4_lut_adj_1437.LUT_INIT = 16'h6996;
    SB_LUT4 i30_4_lut_adj_1438 (.I0(n59), .I1(\data_out_frame[14] [6]), 
            .I2(n52), .I3(\data_out_frame[14] [0]), .O(n64));
    defparam i30_4_lut_adj_1438.LUT_INIT = 16'h6996;
    SB_LUT4 i23_4_lut (.I0(\data_out_frame[13] [6]), .I1(\data_out_frame[16] [0]), 
            .I2(\data_out_frame[14] [4]), .I3(n16729), .O(n57));
    defparam i23_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i31_4_lut_adj_1439 (.I0(n53), .I1(n55), .I2(n54), .I3(n56), 
            .O(n65_adj_4491));
    defparam i31_4_lut_adj_1439.LUT_INIT = 16'h6996;
    SB_LUT4 i33_4_lut_adj_1440 (.I0(n65_adj_4491), .I1(n57), .I2(n64), 
            .I3(n58), .O(n37570));
    defparam i33_4_lut_adj_1440.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1441 (.I0(\data_out_frame[17] [2]), .I1(\data_out_frame[15] [4]), 
            .I2(\data_out_frame[18] [5]), .I3(n16163), .O(n42_adj_4492));
    defparam i18_4_lut_adj_1441.LUT_INIT = 16'h6996;
    SB_LUT4 i22_4_lut_adj_1442 (.I0(n37), .I1(n39_adj_4490), .I2(n38), 
            .I3(n40_adj_4489), .O(n46_adj_4493));
    defparam i22_4_lut_adj_1442.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1443 (.I0(\data_out_frame[19] [1]), .I1(n37570), 
            .I2(\data_out_frame[18] [0]), .I3(\data_out_frame[17] [3]), 
            .O(n41_adj_4494));
    defparam i17_4_lut_adj_1443.LUT_INIT = 16'h9669;
    SB_LUT4 i2_4_lut_adj_1444 (.I0(n35321), .I1(n41_adj_4494), .I2(n46_adj_4493), 
            .I3(n42_adj_4492), .O(n35322));
    defparam i2_4_lut_adj_1444.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1445 (.I0(n35070), .I1(\data_out_frame[20] [1]), 
            .I2(n35322), .I3(n35382), .O(n10_adj_4495));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1445.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_1446 (.I0(\data_out_frame[20] [4]), .I1(n10_adj_4495), 
            .I2(\data_out_frame[20] [7]), .I3(GND_net), .O(n31178));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_adj_1446.LUT_INIT = 16'h9696;
    SB_LUT4 i3_2_lut_adj_1447 (.I0(n35611), .I1(n35330), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4496));
    defparam i3_2_lut_adj_1447.LUT_INIT = 16'h6666;
    SB_LUT4 select_340_Select_11_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [11]), .O(n3_adj_4344));
    defparam select_340_Select_11_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i5_4_lut_adj_1448 (.I0(n31178), .I1(n35530), .I2(n31504), 
            .I3(n31140), .O(n13_adj_4497));
    defparam i5_4_lut_adj_1448.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1449 (.I0(n13_adj_4497), .I1(n11_adj_4496), .I2(\data_out_frame[19] [5]), 
            .I3(n31595), .O(n36904));
    defparam i7_4_lut_adj_1449.LUT_INIT = 16'h9669;
    SB_LUT4 equal_122_i10_2_lut_3_lut (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(GND_net), .O(n10_adj_4424));   // verilog/coms.v(154[7:23])
    defparam equal_122_i10_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_adj_1450 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[6] [1]), 
            .I2(\data_out_frame[5] [7]), .I3(GND_net), .O(n35478));
    defparam i2_3_lut_adj_1450.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1451 (.I0(\data_out_frame[6] [6]), .I1(n35432), 
            .I2(GND_net), .I3(GND_net), .O(n35041));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1451.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1452 (.I0(n35041), .I1(n35113), .I2(n35478), 
            .I3(n6_adj_4498), .O(n31254));   // verilog/coms.v(70[16:27])
    defparam i4_4_lut_adj_1452.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1453 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[19] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n35448));
    defparam i1_2_lut_adj_1453.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1454 (.I0(\data_out_frame[13] [2]), .I1(n31254), 
            .I2(GND_net), .I3(GND_net), .O(n31504));
    defparam i1_2_lut_adj_1454.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1455 (.I0(\data_in_frame[9] [0]), .I1(n31068), 
            .I2(n16142), .I3(\data_in_frame[8] [6]), .O(n37407));
    defparam i3_4_lut_adj_1455.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1456 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(n38499), .I3(GND_net), .O(n34984));   // verilog/coms.v(154[7:23])
    defparam i2_2_lut_3_lut_adj_1456.LUT_INIT = 16'hefef;
    SB_LUT4 select_340_Select_10_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [10]), .O(n3_adj_4342));
    defparam select_340_Select_10_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_3_lut_adj_1457 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [4]), 
            .I2(\data_in_frame[6] [6]), .I3(GND_net), .O(n35590));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_3_lut_adj_1457.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1458 (.I0(\data_out_frame[17] [4]), .I1(n35151), 
            .I2(GND_net), .I3(GND_net), .O(n16982));
    defparam i1_2_lut_adj_1458.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1459 (.I0(n30618), .I1(n35119), .I2(GND_net), 
            .I3(GND_net), .O(n7_adj_4499));
    defparam i2_2_lut_adj_1459.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1460 (.I0(n7_adj_4499), .I1(n16982), .I2(n31504), 
            .I3(n35448), .O(n37556));
    defparam i4_4_lut_adj_1460.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1461 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [4]), 
            .I2(n16782), .I3(n16555), .O(Kp_23__N_1186));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_4_lut_adj_1461.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1462 (.I0(\data_in_frame[6] [3]), .I1(n17042), 
            .I2(\data_in_frame[8] [4]), .I3(GND_net), .O(n35122));   // verilog/coms.v(72[16:42])
    defparam i1_2_lut_3_lut_adj_1462.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1463 (.I0(\data_out_frame[8] [6]), .I1(n16530), 
            .I2(n35196), .I3(n6_adj_4428), .O(n14129));   // verilog/coms.v(74[16:27])
    defparam i4_4_lut_adj_1463.LUT_INIT = 16'h6996;
    SB_LUT4 select_340_Select_9_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [9]), .O(n3_adj_4340));
    defparam select_340_Select_9_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i4_4_lut_adj_1464 (.I0(\data_out_frame[10] [4]), .I1(n1608), 
            .I2(\data_out_frame[13] [0]), .I3(n35596), .O(n10_adj_4310));
    defparam i4_4_lut_adj_1464.LUT_INIT = 16'h6996;
    SB_LUT4 select_340_Select_8_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [8]), .O(n3_adj_4338));
    defparam select_340_Select_8_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i2_3_lut_adj_1465 (.I0(\data_out_frame[13] [1]), .I1(n35151), 
            .I2(n14129), .I3(GND_net), .O(n16729));
    defparam i2_3_lut_adj_1465.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1466 (.I0(\data_out_frame[15] [2]), .I1(\data_out_frame[19] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35119));
    defparam i1_2_lut_adj_1466.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_adj_1467 (.I0(n16729), .I1(\data_out_frame[17] [3]), 
            .I2(n35161), .I3(GND_net), .O(n35330));
    defparam i1_3_lut_adj_1467.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1468 (.I0(n16806), .I1(n35330), .I2(n35119), 
            .I3(\data_out_frame[19] [3]), .O(n36199));
    defparam i3_4_lut_adj_1468.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1469 (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[12] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35481));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_adj_1469.LUT_INIT = 16'h6666;
    SB_LUT4 i804_2_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1608));   // verilog/coms.v(70[16:27])
    defparam i804_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1470 (.I0(\data_out_frame[11] [5]), .I1(n16949), 
            .I2(\data_out_frame[7] [0]), .I3(\data_out_frame[11] [3]), .O(n35054));
    defparam i3_4_lut_adj_1470.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1471 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[8] [6]), 
            .I2(\data_out_frame[8] [7]), .I3(GND_net), .O(n35432));
    defparam i2_3_lut_adj_1471.LUT_INIT = 16'h9696;
    SB_LUT4 select_340_Select_7_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [7]), .O(n3_adj_4336));
    defparam select_340_Select_7_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i2_3_lut_adj_1472 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[11] [0]), 
            .I2(\data_out_frame[10] [6]), .I3(GND_net), .O(n35593));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1472.LUT_INIT = 16'h9696;
    SB_LUT4 i10_4_lut_adj_1473 (.I0(\data_out_frame[10] [4]), .I1(n35076), 
            .I2(n35125), .I3(n35593), .O(n28_adj_4306));
    defparam i10_4_lut_adj_1473.LUT_INIT = 16'h6996;
    SB_LUT4 i8_3_lut (.I0(n1205), .I1(n31464), .I2(n4_c), .I3(GND_net), 
            .O(n26_adj_4500));
    defparam i8_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1474 (.I0(\data_in_frame[6] [3]), .I1(n17042), 
            .I2(n37407), .I3(n35327), .O(n37597));   // verilog/coms.v(72[16:42])
    defparam i2_3_lut_4_lut_adj_1474.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1475 (.I0(\data_out_frame[10] [7]), .I1(n35651), 
            .I2(n16006), .I3(n35572), .O(n30_adj_4501));
    defparam i12_4_lut_adj_1475.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1476 (.I0(n35432), .I1(n32), .I2(n26_adj_4500), 
            .I3(n35054), .O(n34));
    defparam i16_4_lut_adj_1476.LUT_INIT = 16'h6996;
    SB_LUT4 i11_4_lut_adj_1477 (.I0(\data_out_frame[10] [1]), .I1(n35490), 
            .I2(n35657), .I3(\data_out_frame[11] [2]), .O(n29_adj_4502));
    defparam i11_4_lut_adj_1477.LUT_INIT = 16'h6996;
    SB_LUT4 i2_4_lut_adj_1478 (.I0(n35469), .I1(n29_adj_4502), .I2(n34), 
            .I3(n30_adj_4501), .O(n10_adj_4503));
    defparam i2_4_lut_adj_1478.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1479 (.I0(\data_out_frame[12] [5]), .I1(n17071), 
            .I2(n35209), .I3(n30704), .O(n14_adj_4504));
    defparam i6_4_lut_adj_1479.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1480 (.I0(n1608), .I1(n14_adj_4504), .I2(n10_adj_4503), 
            .I3(n35206), .O(n30558));
    defparam i7_4_lut_adj_1480.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1481 (.I0(n30558), .I1(\data_out_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35397));
    defparam i1_2_lut_adj_1481.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1482 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n35657));
    defparam i1_2_lut_adj_1482.LUT_INIT = 16'h6666;
    SB_LUT4 select_340_Select_6_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [6]), .O(n3_adj_4334));
    defparam select_340_Select_6_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_4_lut_adj_1483 (.I0(\data_out_frame[15] [1]), .I1(n30558), 
            .I2(n8_adj_4426), .I3(n35481), .O(n35161));
    defparam i1_4_lut_adj_1483.LUT_INIT = 16'h9669;
    SB_LUT4 i4_4_lut_adj_1484 (.I0(n35584), .I1(n35161), .I2(n14123), 
            .I3(n35654), .O(n10_adj_4505));
    defparam i4_4_lut_adj_1484.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1485 (.I0(\data_out_frame[17] [2]), .I1(n35469), 
            .I2(n10_adj_4505), .I3(\data_out_frame[14] [6]), .O(n30618));
    defparam i1_4_lut_adj_1485.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1486 (.I0(\data_out_frame[19] [3]), .I1(\data_out_frame[19] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35236));
    defparam i1_2_lut_adj_1486.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1487 (.I0(n14180), .I1(n35236), .I2(n16806), 
            .I3(n30618), .O(n36181));
    defparam i3_4_lut_adj_1487.LUT_INIT = 16'h6996;
    SB_LUT4 select_340_Select_5_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [5]), .O(n3_adj_4332));
    defparam select_340_Select_5_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i2_3_lut_adj_1488 (.I0(\data_out_frame[19] [1]), .I1(n35291), 
            .I2(\data_out_frame[19] [2]), .I3(GND_net), .O(n36758));
    defparam i2_3_lut_adj_1488.LUT_INIT = 16'h6969;
    SB_LUT4 select_340_Select_4_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [4]), .O(n3_adj_4330));
    defparam select_340_Select_4_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i2_3_lut_adj_1489 (.I0(n16345), .I1(\data_out_frame[10] [2]), 
            .I2(\data_out_frame[10] [3]), .I3(GND_net), .O(n35572));
    defparam i2_3_lut_adj_1489.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1490 (.I0(n16870), .I1(n35064), .I2(GND_net), 
            .I3(GND_net), .O(n14123));
    defparam i1_2_lut_adj_1490.LUT_INIT = 16'h6666;
    SB_LUT4 i2_2_lut_adj_1491 (.I0(n35457), .I1(\data_out_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4506));
    defparam i2_2_lut_adj_1491.LUT_INIT = 16'h6666;
    SB_LUT4 select_340_Select_3_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [3]), .O(n3_adj_4328));
    defparam select_340_Select_3_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i6_4_lut_adj_1492 (.I0(n35635), .I1(n14123), .I2(n35324), 
            .I3(\data_out_frame[19] [0]), .O(n14_adj_4507));
    defparam i6_4_lut_adj_1492.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1493 (.I0(\data_out_frame[19] [1]), .I1(n14_adj_4507), 
            .I2(n10_adj_4506), .I3(\data_out_frame[12] [4]), .O(n37044));
    defparam i7_4_lut_adj_1493.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1494 (.I0(n2774), .I1(n3), .I2(n23[1]), 
            .I3(n63), .O(n34329));
    defparam i1_2_lut_3_lut_4_lut_adj_1494.LUT_INIT = 16'he0ee;
    SB_LUT4 i1_2_lut_adj_1495 (.I0(\data_out_frame[16] [3]), .I1(n30630), 
            .I2(GND_net), .I3(GND_net), .O(n31552));
    defparam i1_2_lut_adj_1495.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1496 (.I0(n2774), .I1(n3), .I2(n15994), 
            .I3(n3894), .O(n5_adj_4));
    defparam i1_2_lut_3_lut_4_lut_adj_1496.LUT_INIT = 16'heeef;
    SB_LUT4 i1_2_lut_adj_1497 (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[12] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n17071));
    defparam i1_2_lut_adj_1497.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1498 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[12] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17033));
    defparam i1_2_lut_adj_1498.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1499 (.I0(\data_out_frame[7] [7]), .I1(n30584), 
            .I2(\data_out_frame[10] [4]), .I3(\data_out_frame[10] [3]), 
            .O(n35262));
    defparam i3_4_lut_adj_1499.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1500 (.I0(n24684), .I1(rx_data_ready), 
            .I2(\FRAME_MATCHER.rx_data_ready_prev ), .I3(n10_adj_4425), 
            .O(n35006));
    defparam i1_2_lut_3_lut_4_lut_adj_1500.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1501 (.I0(n16239), .I1(n16716), .I2(\data_out_frame[8] [5]), 
            .I3(\data_out_frame[10] [7]), .O(n35196));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1501.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1502 (.I0(n16239), .I1(n16716), .I2(\data_out_frame[8] [5]), 
            .I3(n35593), .O(n6_adj_4498));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1502.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1503 (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[17] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4509));
    defparam i1_2_lut_adj_1503.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1504 (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[14] [6]), 
            .I2(n35451), .I3(n6_adj_4509), .O(n35457));
    defparam i4_4_lut_adj_1504.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1505 (.I0(\data_out_frame[12] [5]), .I1(n16716), 
            .I2(n35262), .I3(n16445), .O(n35565));
    defparam i3_4_lut_adj_1505.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1506 (.I0(\data_out_frame[17] [0]), .I1(\data_out_frame[18] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35608));
    defparam i1_2_lut_adj_1506.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1507 (.I0(n35457), .I1(n35584), .I2(n35132), 
            .I3(GND_net), .O(n14180));
    defparam i2_3_lut_adj_1507.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1508 (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[15] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35647));
    defparam i1_2_lut_adj_1508.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1509 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35113));
    defparam i1_2_lut_adj_1509.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1510 (.I0(\data_out_frame[5] [7]), .I1(n35141), 
            .I2(GND_net), .I3(GND_net), .O(n16716));
    defparam i1_2_lut_adj_1510.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1511 (.I0(n14107), .I1(n35654), .I2(\data_out_frame[14] [5]), 
            .I3(\data_out_frame[17] [1]), .O(n35132));
    defparam i3_4_lut_adj_1511.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1512 (.I0(\data_out_frame[7] [7]), .I1(n17033), 
            .I2(n17071), .I3(\data_out_frame[16] [7]), .O(n35460));
    defparam i3_4_lut_adj_1512.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1513 (.I0(n16587), .I1(n35460), .I2(n35132), 
            .I3(\data_out_frame[12] [4]), .O(n16806));
    defparam i3_4_lut_adj_1513.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1514 (.I0(\data_out_frame[16] [5]), .I1(n14180), 
            .I2(n35635), .I3(n35608), .O(n10_adj_4510));
    defparam i4_4_lut_adj_1514.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1515 (.I0(\data_out_frame[14] [5]), .I1(n10_adj_4510), 
            .I2(\data_out_frame[14] [6]), .I3(GND_net), .O(n35291));
    defparam i5_3_lut_adj_1515.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1516 (.I0(\data_out_frame[19] [0]), .I1(n35611), 
            .I2(GND_net), .I3(GND_net), .O(n35321));
    defparam i1_2_lut_adj_1516.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1517 (.I0(\data_out_frame[20] [7]), .I1(n35321), 
            .I2(n35291), .I3(n16806), .O(n36416));
    defparam i3_4_lut_adj_1517.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1518 (.I0(\data_out_frame[11] [4]), .I1(\data_out_frame[9] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n16949));
    defparam i1_2_lut_adj_1518.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1519 (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[14] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35484));
    defparam i1_2_lut_adj_1519.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1520 (.I0(n30598), .I1(\data_out_frame[11] [6]), 
            .I2(n35230), .I3(n16482), .O(n35206));
    defparam i3_4_lut_adj_1520.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1521 (.I0(\data_out_frame[6] [6]), .I1(\data_out_frame[6] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35242));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1521.LUT_INIT = 16'h6666;
    SB_LUT4 select_340_Select_2_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [2]), .O(n3_adj_4326));
    defparam select_340_Select_2_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_adj_1522 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35496));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1522.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1523 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16530));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1523.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1524 (.I0(n16530), .I1(n35496), .I2(n35242), 
            .I3(\data_out_frame[6] [4]), .O(n1205));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_1524.LUT_INIT = 16'h6996;
    SB_LUT4 i31734_2_lut_3_lut_4_lut (.I0(n24684), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(\FRAME_MATCHER.i [3]), .O(n38499));
    defparam i31734_2_lut_3_lut_4_lut.LUT_INIT = 16'h0400;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1525 (.I0(\data_out_frame[18] [5]), .I1(n37560), 
            .I2(\data_out_frame[16] [3]), .I3(n30630), .O(n35611));
    defparam i1_2_lut_3_lut_4_lut_adj_1525.LUT_INIT = 16'h6996;
    SB_LUT4 select_340_Select_1_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [1]), .O(n3_adj_4324));
    defparam select_340_Select_1_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i19337_3_lut_4_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(n15765), .I3(\FRAME_MATCHER.i [31]), .O(n2957));
    defparam i19337_3_lut_4_lut.LUT_INIT = 16'h00f8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1526 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[7] [4]), .I3(n35605), .O(n16482));
    defparam i1_2_lut_3_lut_4_lut_adj_1526.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1527 (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[14] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n16214));
    defparam i1_2_lut_adj_1527.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1528 (.I0(\data_out_frame[12] [1]), .I1(n35209), 
            .I2(\data_out_frame[11] [7]), .I3(\data_out_frame[10] [0]), 
            .O(n10_adj_4511));
    defparam i4_4_lut_adj_1528.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1529 (.I0(n16482), .I1(n10_adj_4511), .I2(n16821), 
            .I3(GND_net), .O(n30598));
    defparam i5_3_lut_adj_1529.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1530 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35060));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_adj_1530.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1531 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(n35499), .O(n16360));
    defparam i1_2_lut_3_lut_4_lut_adj_1531.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1532 (.I0(\data_out_frame[5] [6]), .I1(n16252), 
            .I2(n35060), .I3(n6_adj_4308), .O(n16445));   // verilog/coms.v(84[17:28])
    defparam i4_4_lut_adj_1532.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1533 (.I0(n16937), .I1(n35057), .I2(\data_out_frame[12] [3]), 
            .I3(\data_out_frame[10] [2]), .O(n12_adj_4512));
    defparam i5_4_lut_adj_1533.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1534 (.I0(n31464), .I1(n12_adj_4512), .I2(n35422), 
            .I3(n16445), .O(n31478));
    defparam i6_4_lut_adj_1534.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1535 (.I0(n35206), .I1(n35484), .I2(\data_out_frame[13] [7]), 
            .I3(GND_net), .O(n30630));
    defparam i2_3_lut_adj_1535.LUT_INIT = 16'h9696;
    SB_LUT4 select_340_Select_0_i3_2_lut_4_lut (.I0(n24684), .I1(n15722), 
            .I2(n15886), .I3(\FRAME_MATCHER.i [0]), .O(n3_c));
    defparam select_340_Select_0_i3_2_lut_4_lut.LUT_INIT = 16'ha800;
    SB_LUT4 i1_2_lut_adj_1536 (.I0(\data_out_frame[7] [1]), .I1(\data_out_frame[7] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n35076));   // verilog/coms.v(84[17:70])
    defparam i1_2_lut_adj_1536.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1537 (.I0(\FRAME_MATCHER.state[1] ), .I1(\FRAME_MATCHER.state [0]), 
            .I2(\FRAME_MATCHER.state [2]), .I3(GND_net), .O(n15886));
    defparam i1_2_lut_3_lut_adj_1537.LUT_INIT = 16'hfefe;
    SB_LUT4 i2_3_lut_4_lut_adj_1538 (.I0(\FRAME_MATCHER.state[1] ), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n15722), .I3(\FRAME_MATCHER.state [2]), .O(n15950));
    defparam i2_3_lut_4_lut_adj_1538.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_adj_1539 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[9] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n16006));   // verilog/coms.v(84[17:63])
    defparam i1_2_lut_adj_1539.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1540 (.I0(\data_out_frame[7] [2]), .I1(\data_out_frame[7] [3]), 
            .I2(\data_out_frame[9] [6]), .I3(\data_out_frame[7] [4]), .O(n35400));
    defparam i1_2_lut_3_lut_4_lut_adj_1540.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1541 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[11] [5]), 
            .I2(n1286), .I3(GND_net), .O(n35230));
    defparam i2_3_lut_adj_1541.LUT_INIT = 16'h9696;
    SB_LUT4 i13331_3_lut_4_lut (.I0(n8_adj_4391), .I1(n35006), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n18070));
    defparam i13331_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1542 (.I0(n4_c), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[6] [0]), .I3(n35057), .O(n16587));
    defparam i1_2_lut_3_lut_4_lut_adj_1542.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1543 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[7] [0]), .I3(n35230), .O(n10_adj_4513));
    defparam i4_4_lut_adj_1543.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1544 (.I0(\data_out_frame[9] [1]), .I1(n10_adj_4513), 
            .I2(\data_out_frame[14] [0]), .I3(n35221), .O(n35505));
    defparam i5_4_lut_adj_1544.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1545 (.I0(\data_out_frame[9] [5]), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n35605));
    defparam i1_2_lut_adj_1545.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1546 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[9] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n35256));   // verilog/coms.v(84[17:63])
    defparam i1_2_lut_adj_1546.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1547 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17080));
    defparam i1_2_lut_adj_1547.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1548 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [6]), 
            .I2(\data_in_frame[1] [0]), .I3(\data_in_frame[3] [2]), .O(n6_adj_4286));
    defparam i1_2_lut_3_lut_4_lut_adj_1548.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1549 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[7] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35032));   // verilog/coms.v(84[17:63])
    defparam i1_2_lut_adj_1549.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1550 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[10] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35404));
    defparam i1_2_lut_adj_1550.LUT_INIT = 16'h6666;
    SB_LUT4 i13332_3_lut_4_lut (.I0(n8_adj_4391), .I1(n35006), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n18071));
    defparam i13332_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1551 (.I0(\data_out_frame[5] [4]), .I1(\data_out_frame[5] [3]), 
            .I2(\data_out_frame[7] [5]), .I3(GND_net), .O(n16821));
    defparam i2_3_lut_adj_1551.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1552 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4309));   // verilog/coms.v(84[17:70])
    defparam i1_2_lut_adj_1552.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1553 (.I0(n4_c), .I1(\data_out_frame[5] [5]), 
            .I2(\data_out_frame[6] [0]), .I3(n35572), .O(n35064));
    defparam i1_2_lut_3_lut_4_lut_adj_1553.LUT_INIT = 16'h6996;
    SB_LUT4 i13333_3_lut_4_lut (.I0(n8_adj_4391), .I1(n35006), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n18072));
    defparam i13333_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1554 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[5] [5]), .I3(\data_out_frame[5] [4]), .O(n16870));
    defparam i1_2_lut_3_lut_4_lut_adj_1554.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1555 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n16252));   // verilog/coms.v(84[17:28])
    defparam i1_2_lut_adj_1555.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1556 (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(n35404), .I3(n35032), .O(n35125));
    defparam i3_4_lut_adj_1556.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1557 (.I0(\data_in_frame[18] [2]), .I1(n30807), 
            .I2(n31530), .I3(GND_net), .O(n31528));
    defparam i1_2_lut_3_lut_adj_1557.LUT_INIT = 16'h6969;
    SB_LUT4 i3_4_lut_adj_1558 (.I0(n16252), .I1(n35651), .I2(n35400), 
            .I3(\data_out_frame[5] [0]), .O(n35033));   // verilog/coms.v(84[17:63])
    defparam i3_4_lut_adj_1558.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1559 (.I0(n16870), .I1(n35125), .I2(n16587), 
            .I3(GND_net), .O(n35451));   // verilog/coms.v(72[16:42])
    defparam i2_3_lut_adj_1559.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1560 (.I0(n35033), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[12] [0]), .I3(GND_net), .O(n30704));   // verilog/coms.v(84[17:63])
    defparam i2_3_lut_adj_1560.LUT_INIT = 16'h9696;
    SB_LUT4 i13334_3_lut_4_lut (.I0(n8_adj_4391), .I1(n35006), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n18073));
    defparam i13334_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1561 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[14] [3]), 
            .I2(\data_out_frame[14] [2]), .I3(n6_adj_4423), .O(n37560));
    defparam i4_4_lut_adj_1561.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1562 (.I0(n35605), .I1(\data_out_frame[16] [2]), 
            .I2(\data_out_frame[14] [1]), .I3(n35505), .O(n15_adj_4514));
    defparam i6_4_lut_adj_1562.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1563 (.I0(n15_adj_4514), .I1(n35242), .I2(n14_adj_4419), 
            .I3(n16949), .O(n36894));
    defparam i8_4_lut_adj_1563.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1564 (.I0(\data_out_frame[16] [5]), .I1(n37560), 
            .I2(GND_net), .I3(GND_net), .O(n35324));
    defparam i1_2_lut_adj_1564.LUT_INIT = 16'h9999;
    SB_LUT4 i19991_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n24712));
    defparam i19991_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i13335_3_lut_4_lut (.I0(n8_adj_4391), .I1(n35006), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n18074));
    defparam i13335_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1565 (.I0(n30630), .I1(\data_out_frame[16] [3]), 
            .I2(n6_adj_4418), .I3(n31478), .O(n35306));
    defparam i1_4_lut_adj_1565.LUT_INIT = 16'h6996;
    SB_LUT4 i13324_3_lut_4_lut (.I0(n8_adj_4399), .I1(n35006), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n18063));
    defparam i13324_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13336_3_lut_4_lut (.I0(n8_adj_4391), .I1(n35006), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n18075));
    defparam i13336_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1566 (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n35527));
    defparam i1_2_lut_adj_1566.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1567 (.I0(\FRAME_MATCHER.state[1] ), .I1(n15963), 
            .I2(n34898), .I3(GND_net), .O(n17205));   // verilog/coms.v(127[12] 295[6])
    defparam i2_3_lut_adj_1567.LUT_INIT = 16'h1010;
    SB_LUT4 i13337_3_lut_4_lut (.I0(n8_adj_4391), .I1(n35006), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n18076));
    defparam i13337_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1568 (.I0(\data_out_frame[20] [7]), .I1(n35527), 
            .I2(n35306), .I3(\data_out_frame[20] [6]), .O(n36265));
    defparam i3_4_lut_adj_1568.LUT_INIT = 16'h6996;
    SB_LUT4 i13338_3_lut_4_lut (.I0(n8_adj_4391), .I1(n35006), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n18077));
    defparam i13338_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1569 (.I0(\data_in_frame[22] [5]), .I1(\data_in_frame[20] [3]), 
            .I2(\data_in_frame[20] [4]), .I3(GND_net), .O(n6_adj_4304));
    defparam i1_2_lut_3_lut_adj_1569.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1570 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[1] [1]), 
            .I2(n35581), .I3(\data_in_frame[1] [3]), .O(n16115));   // verilog/coms.v(72[16:34])
    defparam i2_3_lut_4_lut_adj_1570.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1571 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[2] [6]), 
            .I2(\data_in_frame[3] [0]), .I3(\data_in_frame[0] [5]), .O(n35245));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_4_lut_adj_1571.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1572 (.I0(\data_in_frame[5] [5]), .I1(\data_in_frame[3] [3]), 
            .I2(\data_in_frame[3] [4]), .I3(GND_net), .O(n35581));   // verilog/coms.v(72[16:34])
    defparam i1_2_lut_3_lut_adj_1572.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1573 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[1] [5]), .I3(n35098), .O(n35416));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_4_lut_adj_1573.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_4_lut_adj_1574 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [4]), 
            .I2(\data_in_frame[1] [2]), .I3(\data_in_frame[1] [7]), .O(n8_adj_4290));   // verilog/coms.v(77[16:27])
    defparam i3_3_lut_4_lut_adj_1574.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1575 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n6_adj_4289));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1575.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1576 (.I0(\data_in_frame[4] [6]), .I1(n5_adj_4288), 
            .I2(n6_adj_4289), .I3(GND_net), .O(n16876));
    defparam i1_2_lut_3_lut_adj_1576.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1577 (.I0(\data_in_frame[4] [3]), .I1(\data_in_frame[0] [1]), 
            .I2(\data_in_frame[2] [2]), .I3(\data_in_frame[2] [1]), .O(n35413));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_4_lut_adj_1577.LUT_INIT = 16'h6996;
    SB_LUT4 equal_105_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4399));   // verilog/coms.v(154[7:23])
    defparam equal_105_i8_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 equal_104_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4391));   // verilog/coms.v(154[7:23])
    defparam equal_104_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 equal_107_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4320));
    defparam equal_107_i8_2_lut_3_lut.LUT_INIT = 16'hf7f7;
    SB_LUT4 i1_2_lut_4_lut_adj_1578 (.I0(n31480), .I1(\data_out_frame[20] [4]), 
            .I2(n10_adj_4495), .I3(\data_out_frame[20] [7]), .O(n6_adj_4479));
    defparam i1_2_lut_4_lut_adj_1578.LUT_INIT = 16'h6996;
    SB_LUT4 i13262_3_lut_4_lut (.I0(n8_adj_4399), .I1(n34984), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n18001));
    defparam i13262_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13263_3_lut_4_lut (.I0(n8_adj_4399), .I1(n34984), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n18002));
    defparam i13263_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13264_3_lut_4_lut (.I0(n8_adj_4399), .I1(n34984), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n18003));
    defparam i13264_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13265_3_lut_4_lut (.I0(n8_adj_4399), .I1(n34984), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n18004));
    defparam i13265_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13266_3_lut_4_lut (.I0(n8_adj_4399), .I1(n34984), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n18005));
    defparam i13266_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1579 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[3] [5]), 
            .I2(\data_in_frame[5] [7]), .I3(GND_net), .O(n35110));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1579.LUT_INIT = 16'h9696;
    SB_LUT4 i4_3_lut_4_lut (.I0(\data_in_frame[23] [5]), .I1(n8_adj_4278), 
            .I2(n31610), .I3(n35303), .O(n36394));   // verilog/coms.v(75[16:43])
    defparam i4_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_4_lut_adj_1580 (.I0(\data_in_frame[17] [2]), .I1(n37297), 
            .I2(\data_in_frame[20] [0]), .I3(n35259), .O(n18));
    defparam i5_3_lut_4_lut_adj_1580.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1581 (.I0(\data_in_frame[5] [3]), .I1(n15531), 
            .I2(\data_in_frame[9] [4]), .I3(\data_in_frame[9] [3]), .O(n35552));
    defparam i2_3_lut_4_lut_adj_1581.LUT_INIT = 16'h6996;
    SB_LUT4 i13260_3_lut_4_lut (.I0(n8_adj_4399), .I1(n34984), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n17999));
    defparam i13260_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1582 (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[17] [3]), 
            .I2(\data_in_frame[23] [6]), .I3(n37527), .O(n12_adj_4273));
    defparam i2_3_lut_4_lut_adj_1582.LUT_INIT = 16'h9669;
    SB_LUT4 i13261_3_lut_4_lut (.I0(n8_adj_4399), .I1(n34984), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n18000));
    defparam i13261_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1583 (.I0(\data_in_frame[10] [7]), .I1(n37006), 
            .I2(n35518), .I3(GND_net), .O(n30529));
    defparam i1_2_lut_3_lut_adj_1583.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_3_lut_adj_1584 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[6] [2]), 
            .I2(\data_in_frame[8] [3]), .I3(GND_net), .O(n35224));   // verilog/coms.v(71[16:41])
    defparam i1_2_lut_3_lut_adj_1584.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1585 (.I0(n16552), .I1(\data_in_frame[5] [6]), 
            .I2(Kp_23__N_949), .I3(GND_net), .O(n35154));   // verilog/coms.v(70[16:27])
    defparam i2_2_lut_3_lut_adj_1585.LUT_INIT = 16'h9696;
    SB_LUT4 i13259_3_lut_4_lut (.I0(n8_adj_4399), .I1(n34984), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n17998));
    defparam i13259_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1586 (.I0(n15957), .I1(\FRAME_MATCHER.state [2]), 
            .I2(\FRAME_MATCHER.state [0]), .I3(n15722), .O(n24684));
    defparam i2_3_lut_4_lut_adj_1586.LUT_INIT = 16'haa8a;
    SB_LUT4 i1_2_lut_4_lut_adj_1587 (.I0(\data_in_frame[6][7] ), .I1(n21), 
            .I2(n19_adj_4263), .I3(n20), .O(n35578));   // verilog/coms.v(84[17:63])
    defparam i1_2_lut_4_lut_adj_1587.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1588 (.I0(\data_in_frame[4] [4]), .I1(n35104), 
            .I2(n17042), .I3(GND_net), .O(n16156));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_adj_1588.LUT_INIT = 16'h9696;
    SB_LUT4 i13251_3_lut_4_lut (.I0(n24712), .I1(n34998), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n17990));
    defparam i13251_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i5_3_lut_4_lut_adj_1589 (.I0(n31254), .I1(n10_adj_4471), .I2(\data_out_frame[15] [3]), 
            .I3(n31140), .O(n35318));
    defparam i5_3_lut_4_lut_adj_1589.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1590 (.I0(\data_in_frame[8] [2]), .I1(\data_in_frame[7] [2]), 
            .I2(\data_in_frame[7] [1]), .I3(\data_in_frame[8] [1]), .O(n35629));
    defparam i2_3_lut_4_lut_adj_1590.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1591 (.I0(n16115), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n35091));   // verilog/coms.v(73[16:43])
    defparam i1_2_lut_adj_1591.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1592 (.I0(n16231), .I1(n35533), .I2(\data_in_frame[13] [0]), 
            .I3(\data_in_frame[13] [1]), .O(n35555));   // verilog/coms.v(73[16:43])
    defparam i2_3_lut_4_lut_adj_1592.LUT_INIT = 16'h6996;
    SB_LUT4 i13252_3_lut_4_lut (.I0(n24712), .I1(n34998), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n17991));
    defparam i13252_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13253_3_lut_4_lut (.I0(n24712), .I1(n34998), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n17992));
    defparam i13253_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13254_3_lut_4_lut (.I0(n24712), .I1(n34998), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n17993));
    defparam i13254_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13255_3_lut_4_lut (.I0(n24712), .I1(n34998), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n17994));
    defparam i13255_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13256_3_lut_4_lut (.I0(n24712), .I1(n34998), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n17995));
    defparam i13256_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13257_3_lut_4_lut (.I0(n24712), .I1(n34998), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n17996));
    defparam i13257_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13258_3_lut_4_lut (.I0(n24712), .I1(n34998), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n17997));
    defparam i13258_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i2_3_lut_4_lut_adj_1593 (.I0(n31518), .I1(\data_out_frame[20] [5]), 
            .I2(\data_out_frame[20] [6]), .I3(n31480), .O(n37510));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1593.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1594 (.I0(n31470), .I1(n37403), .I2(\data_in_frame[16] [7]), 
            .I3(GND_net), .O(n16838));
    defparam i1_2_lut_3_lut_adj_1594.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_4_lut_adj_1595 (.I0(Kp_23__N_805), .I1(n16812), .I2(n30578), 
            .I3(n16360), .O(n35502));
    defparam i2_3_lut_4_lut_adj_1595.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1596 (.I0(\data_in_frame[17] [1]), .I1(n31470), 
            .I2(n37403), .I3(\data_in_frame[16] [7]), .O(n35259));
    defparam i1_2_lut_3_lut_4_lut_adj_1596.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1597 (.I0(n16239), .I1(\data_out_frame[5] [7]), 
            .I2(n35141), .I3(\data_out_frame[12] [4]), .O(n35469));
    defparam i1_2_lut_3_lut_4_lut_adj_1597.LUT_INIT = 16'h6996;
    SB_LUT4 i13382_3_lut_4_lut (.I0(n24712), .I1(n35006), .I2(rx_data[3]), 
            .I3(\data_in_frame[23] [3]), .O(n18121));
    defparam i13382_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1598 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[9] [7]), 
            .I2(\data_out_frame[5] [5]), .I3(\data_out_frame[5] [4]), .O(n35209));
    defparam i1_2_lut_3_lut_4_lut_adj_1598.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1599 (.I0(\data_in_frame[15] [3]), .I1(\data_in_frame[11] [1]), 
            .I2(n16231), .I3(n35212), .O(n12));   // verilog/coms.v(74[16:43])
    defparam i5_4_lut_adj_1599.LUT_INIT = 16'h6996;
    SB_LUT4 i13381_3_lut_4_lut (.I0(n24712), .I1(n35006), .I2(rx_data[2]), 
            .I3(\data_in_frame[23] [2]), .O(n18120));
    defparam i13381_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i20197_3_lut_4_lut (.I0(n63_adj_3), .I1(n23947), .I2(r_SM_Main_2__N_3585[0]), 
            .I3(tx_active), .O(n24918));
    defparam i20197_3_lut_4_lut.LUT_INIT = 16'haaa8;
    SB_LUT4 i13325_3_lut_4_lut (.I0(n8_adj_4399), .I1(n35006), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n18064));
    defparam i13325_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13326_3_lut_4_lut (.I0(n8_adj_4399), .I1(n35006), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n18065));
    defparam i13326_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13380_3_lut_4_lut (.I0(n24712), .I1(n35006), .I2(rx_data[1]), 
            .I3(\data_in_frame[23] [1]), .O(n18119));
    defparam i13380_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13379_3_lut_4_lut (.I0(n24712), .I1(n35006), .I2(rx_data[0]), 
            .I3(\data_in_frame[23] [0]), .O(n18118));
    defparam i13379_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13386_3_lut_4_lut (.I0(n24712), .I1(n35006), .I2(rx_data[7]), 
            .I3(\data_in_frame[23] [7]), .O(n18125));
    defparam i13386_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13385_3_lut_4_lut (.I0(n24712), .I1(n35006), .I2(rx_data[6]), 
            .I3(\data_in_frame[23] [6]), .O(n18124));
    defparam i13385_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13327_3_lut_4_lut (.I0(n8_adj_4399), .I1(n35006), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n18066));
    defparam i13327_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13384_3_lut_4_lut (.I0(n24712), .I1(n35006), .I2(rx_data[5]), 
            .I3(\data_in_frame[23] [5]), .O(n18123));
    defparam i13384_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut (.I0(\byte_transmit_counter[4] ), 
            .I1(\byte_transmit_counter[3] ), .I2(n38651), .I3(n38650), 
            .O(tx_data[7]));   // verilog/coms.v(105[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i31_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i13328_3_lut_4_lut (.I0(n8_adj_4399), .I1(n35006), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n18067));
    defparam i13328_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13383_3_lut_4_lut (.I0(n24712), .I1(n35006), .I2(rx_data[4]), 
            .I3(\data_in_frame[23] [4]), .O(n18122));
    defparam i13383_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i13358_3_lut_4_lut (.I0(n8), .I1(n35006), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n18097));
    defparam i13358_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13357_3_lut_4_lut (.I0(n8), .I1(n35006), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n18096));
    defparam i13357_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i13356_3_lut_4_lut (.I0(n8), .I1(n35006), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n18095));
    defparam i13356_3_lut_4_lut.LUT_INIT = 16'hfe10;
    uart_tx tx (.n17500(n17500), .r_Clock_Count({\r_Clock_Count[8] , \r_Clock_Count[7] , 
            \r_Clock_Count[6] , \r_Clock_Count[5] , \r_Clock_Count[4] , 
            \r_Clock_Count[3] , \r_Clock_Count[2] , \r_Clock_Count[1] , 
            Open_0}), .clk32MHz(clk32MHz), .n17497(n17497), .n17494(n17494), 
            .n17491(n17491), .n17488(n17488), .n17485(n17485), .n17513(n17513), 
            .r_Bit_Index({r_Bit_Index}), .n17510(n17510), .n17506(n17506), 
            .n17503(n17503), .r_SM_Main({r_SM_Main}), .n17637(n17637), 
            .tx_data({tx_data}), .n313(n313), .GND_net(GND_net), .n314(n314), 
            .n315(n315), .n316(n316), .n317(n317), .n318(n318), .n319(n319), 
            .n320(n320), .VCC_net(VCC_net), .n17505(n17505), .tx_o(tx_o), 
            .tx_enable(tx_enable), .n17607(n17607), .n17606(n17606), .tx_active(tx_active), 
            .n17605(n17605), .n19670(n19670), .n4(n4), .n4720(n4720), 
            .n17256(n17256), .n17385(n17385), .n3(n3_adj_5), .\r_SM_Main_2__N_3585[0] (r_SM_Main_2__N_3585[0]), 
            .n8950(n8950), .n29(n29)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(106[10:70])
    uart_rx rx (.clk32MHz(clk32MHz), .n17537(n17537), .r_Bit_Index({r_Bit_Index_adj_14}), 
            .n17540(n17540), .n24794(n24794), .r_SM_Main({\r_SM_Main[2]_adj_10 , 
            \r_SM_Main[1]_adj_9 , Open_1}), .rx_data_ready(rx_data_ready), 
            .r_Rx_Data(r_Rx_Data), .PIN_13_N_105(PIN_13_N_105), .GND_net(GND_net), 
            .VCC_net(VCC_net), .n15851(n15851), .n15740(n15740), .n17250(n17250), 
            .n40690(n40690), .n40689(n40689), .n17656(n17656), .rx_data({rx_data}), 
            .n17623(n17623), .n17622(n17622), .n17621(n17621), .n17620(n17620), 
            .n17619(n17619), .n17618(n17618), .n17598(n17598), .n17541(n17541), 
            .n43694(n43694), .n17376(n17376), .n4698(n4698), .n23989(n23989), 
            .n4(n4_adj_11), .n4_adj_1(n4_adj_12), .n4_adj_2(n4_adj_13)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;   // verilog/coms.v(92[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (n17500, r_Clock_Count, clk32MHz, n17497, n17494, n17491, 
            n17488, n17485, n17513, r_Bit_Index, n17510, n17506, 
            n17503, r_SM_Main, n17637, tx_data, n313, GND_net, n314, 
            n315, n316, n317, n318, n319, n320, VCC_net, n17505, 
            tx_o, tx_enable, n17607, n17606, tx_active, n17605, 
            n19670, n4, n4720, n17256, n17385, n3, \r_SM_Main_2__N_3585[0] , 
            n8950, n29) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n17500;
    output [8:0]r_Clock_Count;
    input clk32MHz;
    input n17497;
    input n17494;
    input n17491;
    input n17488;
    input n17485;
    input n17513;
    output [2:0]r_Bit_Index;
    input n17510;
    input n17506;
    input n17503;
    output [2:0]r_SM_Main;
    input n17637;
    input [7:0]tx_data;
    output n313;
    input GND_net;
    output n314;
    output n315;
    output n316;
    output n317;
    output n318;
    output n319;
    output n320;
    input VCC_net;
    output n17505;
    output tx_o;
    output tx_enable;
    input n17607;
    input n17606;
    output tx_active;
    input n17605;
    output n19670;
    output n4;
    output n4720;
    output n17256;
    output n17385;
    output n3;
    input \r_SM_Main_2__N_3585[0] ;
    output n8950;
    output n29;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n18228, n34691;
    wire [8:0]r_Clock_Count_c;   // verilog/uart_tx.v(32[16:29])
    
    wire n13289;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n27941, n27940, n27939, n27938, n27937, n27936, n27935, 
        n27934, n40752, n10, n88, n8, n43811, n43814, n36424, 
        n24402, n43658, o_Tx_Serial_N_3613, n43655;
    
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n17500));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n17497));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n17494));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .D(n17491));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .D(n17488));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i8 (.Q(r_Clock_Count[8]), .C(clk32MHz), .D(n17485));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n17513));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n17510));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n17506));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n17503));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n18228));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n17637));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count_c[0]), .C(clk32MHz), .D(n34691));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(clk32MHz), .E(n13289), 
            .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 add_59_10_lut (.I0(GND_net), .I1(r_Clock_Count[8]), .I2(GND_net), 
            .I3(n27941), .O(n313)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_59_9_lut (.I0(GND_net), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n27940), .O(n314)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_9 (.CI(n27940), .I0(r_Clock_Count[7]), .I1(GND_net), 
            .CO(n27941));
    SB_LUT4 add_59_8_lut (.I0(GND_net), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n27939), .O(n315)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_8 (.CI(n27939), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n27940));
    SB_LUT4 add_59_7_lut (.I0(GND_net), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n27938), .O(n316)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_7 (.CI(n27938), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n27939));
    SB_LUT4 add_59_6_lut (.I0(GND_net), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n27937), .O(n317)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_6 (.CI(n27937), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n27938));
    SB_LUT4 add_59_5_lut (.I0(GND_net), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n27936), .O(n318)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_5 (.CI(n27936), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n27937));
    SB_LUT4 add_59_4_lut (.I0(GND_net), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n27935), .O(n319)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_4 (.CI(n27935), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n27936));
    SB_LUT4 add_59_3_lut (.I0(GND_net), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n27934), .O(n320)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_59_3 (.CI(n27934), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n27935));
    SB_LUT4 add_59_2_lut (.I0(n17505), .I1(r_Clock_Count_c[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n40752)) /* synthesis syn_instantiated=1 */ ;
    defparam add_59_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_59_2 (.CI(VCC_net), .I0(r_Clock_Count_c[0]), .I1(GND_net), 
            .CO(n27934));
    SB_LUT4 i20_3_lut (.I0(r_Clock_Count_c[0]), .I1(n40752), .I2(r_SM_Main[2]), 
            .I3(GND_net), .O(n34691));
    defparam i20_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count_c[0]), 
            .I3(r_Clock_Count[4]), .O(n10));   // verilog/uart_tx.v(32[16:29])
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(r_Clock_Count[5]), .I1(n10), .I2(r_Clock_Count[1]), 
            .I3(GND_net), .O(n88));   // verilog/uart_tx.v(32[16:29])
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i19330_4_lut (.I0(r_SM_Main[2]), .I1(n88), .I2(n8), .I3(r_Clock_Count[7]), 
            .O(n17505));
    defparam i19330_4_lut.LUT_INIT = 16'haaba;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[2]), 
            .I2(r_Tx_Data[3]), .I3(r_Bit_Index[1]), .O(n43811));
    defparam r_Bit_Index_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n43811_bdd_4_lut (.I0(n43811), .I1(r_Tx_Data[1]), .I2(r_Tx_Data[0]), 
            .I3(r_Bit_Index[1]), .O(n43814));
    defparam n43811_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(clk32MHz), .E(n13289), 
            .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(clk32MHz), .E(n13289), 
            .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(clk32MHz), .E(n13289), 
            .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(clk32MHz), .E(n13289), 
            .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(clk32MHz), .E(n13289), 
            .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(clk32MHz), .E(n13289), 
            .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(clk32MHz), .E(n13289), 
            .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(clk32MHz), .D(n17607));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(clk32MHz), .D(n17606));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFF o_Tx_Serial_45 (.Q(tx_o), .C(clk32MHz), .D(n17605));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i3_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(n19670), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main[2]), .O(n36424));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h0080;
    SB_LUT4 i13489_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(n19670), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main[2]), .O(n18228));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i13489_3_lut_4_lut.LUT_INIT = 16'h0078;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[0]), .I1(n19670), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main[2]), .O(n4));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h008f;
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(n36424));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1337_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4720));   // verilog/uart_tx.v(98[36:51])
    defparam i1337_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n24402));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[8]), .I1(r_Clock_Count[6]), .I2(r_Clock_Count[7]), 
            .I3(n88), .O(n19670));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i3_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main[2]), .I2(r_SM_Main[1]), 
            .I3(n19670), .O(n17256));
    defparam i2_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i12646_3_lut (.I0(n17256), .I1(r_SM_Main[1]), .I2(n24402), 
            .I3(GND_net), .O(n17385));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i12646_3_lut.LUT_INIT = 16'ha2a2;
    SB_LUT4 i2031336_i1_3_lut (.I0(n43814), .I1(n43658), .I2(r_Bit_Index[2]), 
            .I3(GND_net), .O(o_Tx_Serial_N_3613));
    defparam i2031336_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 r_SM_Main_2__I_0_56_i3_3_lut (.I0(r_SM_Main[0]), .I1(o_Tx_Serial_N_3613), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3));   // verilog/uart_tx.v(43[7] 142[14])
    defparam r_SM_Main_2__I_0_56_i3_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_3585[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n8950));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i27_4_lut (.I0(\r_SM_Main_2__N_3585[0] ), .I1(n24402), .I2(r_SM_Main[1]), 
            .I3(n19670), .O(n29));   // verilog/uart_tx.v(31[16:25])
    defparam i27_4_lut.LUT_INIT = 16'hca0a;
    SB_LUT4 r_Bit_Index_0__bdd_4_lut_36939 (.I0(r_Bit_Index[0]), .I1(r_Tx_Data[6]), 
            .I2(r_Tx_Data[7]), .I3(r_Bit_Index[1]), .O(n43655));
    defparam r_Bit_Index_0__bdd_4_lut_36939.LUT_INIT = 16'he4aa;
    SB_LUT4 n43655_bdd_4_lut (.I0(n43655), .I1(r_Tx_Data[5]), .I2(r_Tx_Data[4]), 
            .I3(r_Bit_Index[1]), .O(n43658));
    defparam n43655_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_3_lut_4_lut_adj_995 (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[2]), .I3(\r_SM_Main_2__N_3585[0] ), .O(n13289));   // verilog/uart_tx.v(31[16:25])
    defparam i3_3_lut_4_lut_adj_995.LUT_INIT = 16'h0100;
    SB_LUT4 i3_3_lut_4_lut_adj_996 (.I0(r_SM_Main[1]), .I1(r_SM_Main[0]), 
            .I2(r_Clock_Count[8]), .I3(r_Clock_Count[6]), .O(n8));   // verilog/uart_tx.v(31[16:25])
    defparam i3_3_lut_4_lut_adj_996.LUT_INIT = 16'h000e;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (clk32MHz, n17537, r_Bit_Index, n17540, n24794, r_SM_Main, 
            rx_data_ready, r_Rx_Data, PIN_13_N_105, GND_net, VCC_net, 
            n15851, n15740, n17250, n40690, n40689, n17656, rx_data, 
            n17623, n17622, n17621, n17620, n17619, n17618, n17598, 
            n17541, n43694, n17376, n4698, n23989, n4, n4_adj_1, 
            n4_adj_2) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input clk32MHz;
    input n17537;
    output [2:0]r_Bit_Index;
    input n17540;
    input n24794;
    output [2:0]r_SM_Main;
    output rx_data_ready;
    output r_Rx_Data;
    input PIN_13_N_105;
    input GND_net;
    input VCC_net;
    output n15851;
    output n15740;
    output n17250;
    output n40690;
    output n40689;
    input n17656;
    output [7:0]rx_data;
    input n17623;
    input n17622;
    input n17621;
    input n17620;
    input n17619;
    input n17618;
    input n17598;
    input n17541;
    output n43694;
    output n17376;
    output n4698;
    output n23989;
    output n4;
    output n4_adj_1;
    output n4_adj_2;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n17467;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n17464, n17482, n17479, n17476, n17473, n45, n35697, 
        n34519, n34537, r_Rx_Data_R;
    wire [2:0]r_SM_Main_2__N_3511;
    
    wire n34968;
    wire [31:0]n194;
    
    wire n27933, n27932, n27931, n27930, n27929, n27928, n27927, 
        n35014;
    wire [2:0]r_SM_Main_c;   // verilog/uart_rx.v(36[17:26])
    
    wire n19568, n2586, n34944, n40623, n43691, n24830, n24732, 
        n34993, n37703, n19549, n37488, n6, n6_adj_4256, n17175;
    
    SB_DFF r_Clock_Count__i6 (.Q(r_Clock_Count[6]), .C(clk32MHz), .D(n17467));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i7 (.Q(r_Clock_Count[7]), .C(clk32MHz), .D(n17464));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i1 (.Q(r_Clock_Count[1]), .C(clk32MHz), .D(n17482));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i2 (.Q(r_Clock_Count[2]), .C(clk32MHz), .D(n17479));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i3 (.Q(r_Clock_Count[3]), .C(clk32MHz), .D(n17476));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i4 (.Q(r_Clock_Count[4]), .C(clk32MHz), .D(n17473));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i5 (.Q(r_Clock_Count[5]), .C(clk32MHz), .D(n45));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(clk32MHz), .D(n17537));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(clk32MHz), .D(n17540));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Clock_Count__i0 (.Q(r_Clock_Count[0]), .C(clk32MHz), .D(n35697));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(clk32MHz), .D(n24794));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(clk32MHz), .D(n34519));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(clk32MHz), .D(n34537));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(clk32MHz), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(clk32MHz), .D(PIN_13_N_105));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFFSR r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(clk32MHz), .D(r_SM_Main_2__N_3511[2]), 
            .R(n34968));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 add_62_9_lut (.I0(GND_net), .I1(r_Clock_Count[7]), .I2(GND_net), 
            .I3(n27933), .O(n194[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_62_8_lut (.I0(GND_net), .I1(r_Clock_Count[6]), .I2(GND_net), 
            .I3(n27932), .O(n194[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_8 (.CI(n27932), .I0(r_Clock_Count[6]), .I1(GND_net), 
            .CO(n27933));
    SB_LUT4 add_62_7_lut (.I0(GND_net), .I1(r_Clock_Count[5]), .I2(GND_net), 
            .I3(n27931), .O(n194[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_7 (.CI(n27931), .I0(r_Clock_Count[5]), .I1(GND_net), 
            .CO(n27932));
    SB_LUT4 add_62_6_lut (.I0(GND_net), .I1(r_Clock_Count[4]), .I2(GND_net), 
            .I3(n27930), .O(n194[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_6 (.CI(n27930), .I0(r_Clock_Count[4]), .I1(GND_net), 
            .CO(n27931));
    SB_LUT4 add_62_5_lut (.I0(GND_net), .I1(r_Clock_Count[3]), .I2(GND_net), 
            .I3(n27929), .O(n194[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_5 (.CI(n27929), .I0(r_Clock_Count[3]), .I1(GND_net), 
            .CO(n27930));
    SB_LUT4 add_62_4_lut (.I0(GND_net), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(n27928), .O(n194[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_4 (.CI(n27928), .I0(r_Clock_Count[2]), .I1(GND_net), 
            .CO(n27929));
    SB_LUT4 add_62_3_lut (.I0(GND_net), .I1(r_Clock_Count[1]), .I2(GND_net), 
            .I3(n27927), .O(n194[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_3 (.CI(n27927), .I0(r_Clock_Count[1]), .I1(GND_net), 
            .CO(n27928));
    SB_LUT4 add_62_2_lut (.I0(GND_net), .I1(r_Clock_Count[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n194[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_62_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_62_2 (.CI(VCC_net), .I0(r_Clock_Count[0]), .I1(GND_net), 
            .CO(n27927));
    SB_LUT4 i1_2_lut_4_lut (.I0(r_SM_Main_2__N_3511[2]), .I1(n35014), .I2(r_SM_Main_c[0]), 
            .I3(r_Bit_Index[0]), .O(n15851));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut_4_lut_adj_990 (.I0(r_SM_Main_2__N_3511[2]), .I1(n35014), 
            .I2(r_SM_Main_c[0]), .I3(r_Bit_Index[0]), .O(n15740));
    defparam i1_2_lut_4_lut_adj_990.LUT_INIT = 16'hfffd;
    SB_LUT4 i12_3_lut (.I0(n17250), .I1(r_Bit_Index[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n34537));   // verilog/uart_rx.v(36[17:26])
    defparam i12_3_lut.LUT_INIT = 16'h6464;
    SB_LUT4 i34229_2_lut (.I0(r_SM_Main_2__N_3511[2]), .I1(r_SM_Main_c[0]), 
            .I2(GND_net), .I3(GND_net), .O(n40690));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i34229_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34269_3_lut (.I0(r_SM_Main_c[0]), .I1(n19568), .I2(r_Rx_Data), 
            .I3(GND_net), .O(n40689));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i34269_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i28946_4_lut (.I0(r_Clock_Count[0]), .I1(n194[0]), .I2(n2586), 
            .I3(n34944), .O(n35697));
    defparam i28946_4_lut.LUT_INIT = 16'ha0ac;
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(clk32MHz), .D(n17656));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(clk32MHz), .D(n17623));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i12740_4_lut_4_lut (.I0(n2586), .I1(n34944), .I2(n194[2]), 
            .I3(r_Clock_Count[2]), .O(n17479));
    defparam i12740_4_lut_4_lut.LUT_INIT = 16'hba10;
    SB_LUT4 i12725_4_lut_4_lut (.I0(n2586), .I1(n34944), .I2(n194[7]), 
            .I3(r_Clock_Count[7]), .O(n17464));
    defparam i12725_4_lut_4_lut.LUT_INIT = 16'hba10;
    SB_LUT4 i12728_4_lut_4_lut (.I0(n2586), .I1(n34944), .I2(n194[6]), 
            .I3(r_Clock_Count[6]), .O(n17467));
    defparam i12728_4_lut_4_lut.LUT_INIT = 16'hba10;
    SB_LUT4 i12743_4_lut_4_lut (.I0(n2586), .I1(n34944), .I2(n194[1]), 
            .I3(r_Clock_Count[1]), .O(n17482));
    defparam i12743_4_lut_4_lut.LUT_INIT = 16'hba10;
    SB_LUT4 i12737_4_lut_4_lut (.I0(n2586), .I1(n34944), .I2(n194[3]), 
            .I3(r_Clock_Count[3]), .O(n17476));
    defparam i12737_4_lut_4_lut.LUT_INIT = 16'hba10;
    SB_LUT4 i12734_4_lut_4_lut (.I0(n2586), .I1(n34944), .I2(n194[4]), 
            .I3(r_Clock_Count[4]), .O(n17473));
    defparam i12734_4_lut_4_lut.LUT_INIT = 16'hba10;
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(clk32MHz), .D(n17622));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(clk32MHz), .D(n17621));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1_4_lut_4_lut (.I0(n2586), .I1(n34944), .I2(n194[5]), .I3(r_Clock_Count[5]), 
            .O(n45));
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hba10;
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(clk32MHz), .D(n17620));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(clk32MHz), .D(n17619));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(clk32MHz), .D(n17618));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i0 (.Q(r_SM_Main_c[0]), .C(clk32MHz), .D(n17598));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(clk32MHz), .D(n17541));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_SM_Main_0__bdd_4_lut_4_lut (.I0(r_SM_Main_2__N_3511[2]), .I1(r_SM_Main[1]), 
            .I2(n40623), .I3(r_SM_Main_c[0]), .O(n43691));
    defparam r_SM_Main_0__bdd_4_lut_4_lut.LUT_INIT = 16'h77c0;
    SB_LUT4 n43691_bdd_4_lut_4_lut (.I0(r_Rx_Data), .I1(r_SM_Main[1]), .I2(n19568), 
            .I3(n43691), .O(n43694));   // verilog/uart_rx.v(30[17:26])
    defparam n43691_bdd_4_lut_4_lut.LUT_INIT = 16'hfc11;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n24830));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_3_lut (.I0(r_SM_Main[1]), .I1(n17250), .I2(n24830), .I3(GND_net), 
            .O(n17376));   // verilog/uart_rx.v(36[17:26])
    defparam i1_3_lut.LUT_INIT = 16'hc4c4;
    SB_LUT4 i1315_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n4698));   // verilog/uart_rx.v(102[36:51])
    defparam i1315_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_Clock_Count[5]), .I1(n24732), .I2(r_Clock_Count[7]), 
            .I3(r_Clock_Count[6]), .O(n19568));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main_c[0]), .I2(GND_net), 
            .I3(GND_net), .O(n34993));
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_991 (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(GND_net), 
            .I3(GND_net), .O(n35014));
    defparam i1_2_lut_adj_991.LUT_INIT = 16'hbbbb;
    SB_LUT4 i3_4_lut (.I0(n24732), .I1(r_Clock_Count[6]), .I2(r_Clock_Count[7]), 
            .I3(r_Clock_Count[5]), .O(n37703));
    defparam i3_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i2_4_lut (.I0(n19549), .I1(n35014), .I2(r_Clock_Count[5]), 
            .I3(n24732), .O(n37488));
    defparam i2_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_4_lut (.I0(n37488), .I1(n37703), .I2(n34993), .I3(r_SM_Main[2]), 
            .O(n34944));
    defparam i1_4_lut.LUT_INIT = 16'haaa8;
    SB_LUT4 i1_2_lut_adj_992 (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[6]), 
            .I2(GND_net), .I3(GND_net), .O(n19549));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_adj_992.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_993 (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[3]), 
            .I2(GND_net), .I3(GND_net), .O(n6));
    defparam i1_2_lut_adj_993.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[1]), .I2(r_Clock_Count[2]), 
            .I3(n6), .O(n24732));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i2_2_lut (.I0(n19568), .I1(r_SM_Main_c[0]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4256));
    defparam i2_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i2_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main_c[0]), .I2(r_SM_Main[2]), 
            .I3(r_SM_Main_2__N_3511[2]), .O(n17250));
    defparam i2_4_lut_4_lut.LUT_INIT = 16'h0301;
    SB_LUT4 i1_3_lut_4_lut (.I0(r_Clock_Count[7]), .I1(r_Clock_Count[6]), 
            .I2(r_Clock_Count[5]), .I3(n24732), .O(r_SM_Main_2__N_3511[2]));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_4_lut_adj_994 (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6_adj_4256), 
            .I3(r_Rx_Data), .O(n2586));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_4_lut_adj_994.LUT_INIT = 16'hbaaa;
    SB_LUT4 i19273_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), .I2(GND_net), 
            .I3(GND_net), .O(n23989));
    defparam i19273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 equal_132_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_132_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_134_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_1));   // verilog/uart_rx.v(97[17:39])
    defparam equal_134_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i34131_2_lut_4_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(r_Bit_Index[0]), .I3(r_SM_Main_2__N_3511[2]), .O(n40623));   // verilog/uart_rx.v(36[17:26])
    defparam i34131_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 equal_136_i4_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_2));   // verilog/uart_rx.v(97[17:39])
    defparam equal_136_i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i36746_2_lut_3_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_c[0]), 
            .I3(GND_net), .O(n34968));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i36746_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i13_4_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main_2__N_3511[2]), 
            .I3(r_SM_Main_c[0]), .O(n17175));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i13_4_lut_4_lut.LUT_INIT = 16'h2055;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(n17175), 
            .I3(rx_data_ready), .O(n34519));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h2f20;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100) 
//

module \quad(DEBOUNCE_TICKS=100)  (encoder1_position, GND_net, n18184, 
            clk32MHz, n18185, n18186, n18187, n18188, n18189, n18190, 
            n18181, n18202, n18203, n18200, n18201, n18198, n18199, 
            n18196, n18197, n18194, n18195, n18191, n18192, n18193, 
            n18182, n18183, data_o, n17596, n2942, count_enable, 
            n18229, reg_B, n36342, PIN_6_c_1, PIN_7_c_0, n17608) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    output [23:0]encoder1_position;
    input GND_net;
    input n18184;
    input clk32MHz;
    input n18185;
    input n18186;
    input n18187;
    input n18188;
    input n18189;
    input n18190;
    input n18181;
    input n18202;
    input n18203;
    input n18200;
    input n18201;
    input n18198;
    input n18199;
    input n18196;
    input n18197;
    input n18194;
    input n18195;
    input n18191;
    input n18192;
    input n18193;
    input n18182;
    input n18183;
    output [1:0]data_o;
    input n17596;
    output [23:0]n2942;
    output count_enable;
    input n18229;
    output [1:0]reg_B;
    output n36342;
    input PIN_6_c_1;
    input PIN_7_c_0;
    input n17608;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire n28046, count_direction, n28047, n2929, B_delayed, A_delayed, 
        n28069, n28068, n28067, n28066, n28065, n28064, n28063, 
        n28062, n28061, n28060, n28059, n28058, n28057, n28056, 
        n28055, n28054, n28053, n28052, n28051, n28050, n28049, 
        n28048;
    
    SB_CARRY add_605_2 (.CI(n28046), .I0(encoder1_position[0]), .I1(count_direction), 
            .CO(n28047));
    SB_CARRY add_605_1 (.CI(GND_net), .I0(n2929), .I1(n2929), .CO(n28046));
    SB_DFF count_i0_i4 (.Q(encoder1_position[4]), .C(clk32MHz), .D(n18184));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder1_position[5]), .C(clk32MHz), .D(n18185));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder1_position[6]), .C(clk32MHz), .D(n18186));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder1_position[7]), .C(clk32MHz), .D(n18187));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder1_position[8]), .C(clk32MHz), .D(n18188));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder1_position[9]), .C(clk32MHz), .D(n18189));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder1_position[10]), .C(clk32MHz), .D(n18190));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder1_position[1]), .C(clk32MHz), .D(n18181));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder1_position[22]), .C(clk32MHz), .D(n18202));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder1_position[23]), .C(clk32MHz), .D(n18203));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i20 (.Q(encoder1_position[20]), .C(clk32MHz), .D(n18200));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder1_position[21]), .C(clk32MHz), .D(n18201));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder1_position[18]), .C(clk32MHz), .D(n18198));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder1_position[19]), .C(clk32MHz), .D(n18199));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder1_position[16]), .C(clk32MHz), .D(n18196));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder1_position[17]), .C(clk32MHz), .D(n18197));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder1_position[14]), .C(clk32MHz), .D(n18194));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder1_position[15]), .C(clk32MHz), .D(n18195));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder1_position[11]), .C(clk32MHz), .D(n18191));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder1_position[12]), .C(clk32MHz), .D(n18192));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder1_position[13]), .C(clk32MHz), .D(n18193));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder1_position[2]), .C(clk32MHz), .D(n18182));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder1_position[3]), .C(clk32MHz), .D(n18183));   // quad.v(35[10] 41[6])
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_DFF count_i0_i0 (.Q(encoder1_position[0]), .C(clk32MHz), .D(n17596));   // quad.v(35[10] 41[6])
    SB_LUT4 add_605_25_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(n2929), 
            .I3(n28069), .O(n2942[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_605_24_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(n2929), 
            .I3(n28068), .O(n2942[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_24 (.CI(n28068), .I0(encoder1_position[22]), .I1(n2929), 
            .CO(n28069));
    SB_LUT4 add_605_23_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(n2929), 
            .I3(n28067), .O(n2942[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_23 (.CI(n28067), .I0(encoder1_position[21]), .I1(n2929), 
            .CO(n28068));
    SB_LUT4 add_605_22_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(n2929), 
            .I3(n28066), .O(n2942[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_22 (.CI(n28066), .I0(encoder1_position[20]), .I1(n2929), 
            .CO(n28067));
    SB_LUT4 add_605_21_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(n2929), 
            .I3(n28065), .O(n2942[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_21 (.CI(n28065), .I0(encoder1_position[19]), .I1(n2929), 
            .CO(n28066));
    SB_LUT4 add_605_20_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(n2929), 
            .I3(n28064), .O(n2942[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_20 (.CI(n28064), .I0(encoder1_position[18]), .I1(n2929), 
            .CO(n28065));
    SB_LUT4 add_605_19_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(n2929), 
            .I3(n28063), .O(n2942[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_19 (.CI(n28063), .I0(encoder1_position[17]), .I1(n2929), 
            .CO(n28064));
    SB_LUT4 add_605_18_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(n2929), 
            .I3(n28062), .O(n2942[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_18 (.CI(n28062), .I0(encoder1_position[16]), .I1(n2929), 
            .CO(n28063));
    SB_LUT4 add_605_17_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(n2929), 
            .I3(n28061), .O(n2942[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_17 (.CI(n28061), .I0(encoder1_position[15]), .I1(n2929), 
            .CO(n28062));
    SB_LUT4 add_605_16_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(n2929), 
            .I3(n28060), .O(n2942[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_16 (.CI(n28060), .I0(encoder1_position[14]), .I1(n2929), 
            .CO(n28061));
    SB_LUT4 add_605_15_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(n2929), 
            .I3(n28059), .O(n2942[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_15 (.CI(n28059), .I0(encoder1_position[13]), .I1(n2929), 
            .CO(n28060));
    SB_LUT4 add_605_14_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(n2929), 
            .I3(n28058), .O(n2942[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_14 (.CI(n28058), .I0(encoder1_position[12]), .I1(n2929), 
            .CO(n28059));
    SB_LUT4 add_605_13_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(n2929), 
            .I3(n28057), .O(n2942[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_13 (.CI(n28057), .I0(encoder1_position[11]), .I1(n2929), 
            .CO(n28058));
    SB_LUT4 add_605_12_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(n2929), 
            .I3(n28056), .O(n2942[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_12 (.CI(n28056), .I0(encoder1_position[10]), .I1(n2929), 
            .CO(n28057));
    SB_LUT4 add_605_11_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(n2929), 
            .I3(n28055), .O(n2942[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_11 (.CI(n28055), .I0(encoder1_position[9]), .I1(n2929), 
            .CO(n28056));
    SB_LUT4 add_605_10_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(n2929), 
            .I3(n28054), .O(n2942[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_10 (.CI(n28054), .I0(encoder1_position[8]), .I1(n2929), 
            .CO(n28055));
    SB_LUT4 add_605_9_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(n2929), 
            .I3(n28053), .O(n2942[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_9 (.CI(n28053), .I0(encoder1_position[7]), .I1(n2929), 
            .CO(n28054));
    SB_LUT4 add_605_8_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(n2929), 
            .I3(n28052), .O(n2942[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_8 (.CI(n28052), .I0(encoder1_position[6]), .I1(n2929), 
            .CO(n28053));
    SB_LUT4 add_605_7_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(n2929), 
            .I3(n28051), .O(n2942[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_7 (.CI(n28051), .I0(encoder1_position[5]), .I1(n2929), 
            .CO(n28052));
    SB_LUT4 add_605_6_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(n2929), 
            .I3(n28050), .O(n2942[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_6 (.CI(n28050), .I0(encoder1_position[4]), .I1(n2929), 
            .CO(n28051));
    SB_LUT4 add_605_5_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(n2929), 
            .I3(n28049), .O(n2942[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_5 (.CI(n28049), .I0(encoder1_position[3]), .I1(n2929), 
            .CO(n28050));
    SB_LUT4 add_605_4_lut (.I0(GND_net), .I1(encoder1_position[2]), .I2(n2929), 
            .I3(n28048), .O(n2942[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_4 (.CI(n28048), .I0(encoder1_position[2]), .I1(n2929), 
            .CO(n28049));
    SB_LUT4 add_605_3_lut (.I0(GND_net), .I1(encoder1_position[1]), .I2(n2929), 
            .I3(n28047), .O(n2942[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_605_3 (.CI(n28047), .I0(encoder1_position[1]), .I1(n2929), 
            .CO(n28048));
    SB_LUT4 add_605_2_lut (.I0(GND_net), .I1(encoder1_position[0]), .I2(count_direction), 
            .I3(n28046), .O(n2942[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_605_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i944_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2929));   // quad.v(37[5] 40[8])
    defparam i944_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)  debounce (.n18229(n18229), .data_o({data_o}), .clk32MHz(clk32MHz), 
            .reg_B({reg_B}), .GND_net(GND_net), .n36342(n36342), .PIN_6_c_1(PIN_6_c_1), 
            .PIN_7_c_0(PIN_7_c_0), .n17608(n17608)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5) 
//

module \grp_debouncer(2,5)  (n18229, data_o, clk32MHz, reg_B, GND_net, 
            n36342, PIN_6_c_1, PIN_7_c_0, n17608) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n18229;
    output [1:0]data_o;
    input clk32MHz;
    output [1:0]reg_B;
    input GND_net;
    output n36342;
    input PIN_6_c_1;
    input PIN_7_c_0;
    input n17608;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_2__N_3821;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    wire [2:0]n17;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n18229));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n36342), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3821));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i22834_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22834_1_lut.LUT_INIT = 16'h5555;
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_6_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1227__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3821));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n36342));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_7_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n17608));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1227__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3821));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1227__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3821));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i22843_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22843_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i22836_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22836_2_lut.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (GND_net, \Kp[2] , \Kp[3] , duty, IntegralLimit, 
            \Kp[1] , \Kp[0] , \Kp[4] , \Kp[5] , \Kp[6] , \Kp[7] , 
            \Kp[8] , PWMLimit, \Kp[9] , \Kp[10] , \Kp[11] , \Kp[12] , 
            \Kp[13] , \Kp[14] , \Kp[15] , clk32MHz, VCC_net, n25, 
            \Ki[0] , \Ki[3] , \Ki[2] , \Ki[1] , motor_state, \Ki[4] , 
            \Ki[5] , \Ki[6] , \Ki[7] , \Ki[8] , \Ki[9] , \Ki[10] , 
            \Ki[11] , \Ki[12] , \Ki[13] , \Ki[14] , \Ki[15] , n43653, 
            setpoint) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input GND_net;
    input \Kp[2] ;
    input \Kp[3] ;
    output [23:0]duty;
    input [23:0]IntegralLimit;
    input \Kp[1] ;
    input \Kp[0] ;
    input \Kp[4] ;
    input \Kp[5] ;
    input \Kp[6] ;
    input \Kp[7] ;
    input \Kp[8] ;
    input [23:0]PWMLimit;
    input \Kp[9] ;
    input \Kp[10] ;
    input \Kp[11] ;
    input \Kp[12] ;
    input \Kp[13] ;
    input \Kp[14] ;
    input \Kp[15] ;
    input clk32MHz;
    input VCC_net;
    input n25;
    input \Ki[0] ;
    input \Ki[3] ;
    input \Ki[2] ;
    input \Ki[1] ;
    input [23:0]motor_state;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Ki[6] ;
    input \Ki[7] ;
    input \Ki[8] ;
    input \Ki[9] ;
    input \Ki[10] ;
    input \Ki[11] ;
    input \Ki[12] ;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[15] ;
    output n43653;
    input [23:0]setpoint;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [20:0]n7879;
    wire [19:0]n7902;
    
    wire n29438;
    wire [23:0]duty_23__N_3740;
    wire [23:0]n3048;
    wire [23:0]n3073;
    
    wire n27954;
    wire [23:0]\PID_CONTROLLER.err ;   // verilog/motorControl.v(29[23:26])
    
    wire n180, n28629;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(31[23:31])
    
    wire n28630;
    wire [23:0]n1;
    
    wire n28628, n27955, n253, n47;
    wire [23:0]n1_adj_4253;
    
    wire n28045, n27953, n29437;
    wire [23:0]n1_adj_4254;
    wire [8:0]n8089;
    
    wire n47_adj_3826, n116, n29593, n28627, n29436, n74, n5;
    wire [9:0]n8077;
    
    wire n770, n29592, n29435, n28626;
    wire [23:0]n257;
    
    wire n28044, n697, n29591, n29434, n28625, n28624, n29433, 
        n624, n29590, n1102, n29432, n28623, n28622, n28621, n1029, 
        n29431, n28620, n551, n29589, n956, n29430, n28619, n28043, 
        n28618, n28042, n883, n29429, n478, n29588, n810, n29428, 
        n28041, n28617, n28040, n326, n399, n147, n223, n220, 
        n396, n293, n296, n28039, n28616, n369, n469, n366, 
        n442, n472, n515, n588, n28038, n737, n29427, n542, 
        n545, n618, n664, n29426, n439, n691, n28037, n764, 
        n512, n530, n837, n661, n615, n910, n585, n28615, n734, 
        n110_adj_3833, n41, n688, n183, n603, n676, n749, n256, 
        n822, n658, n731, n804, n895, n968, n1041, n1114, n591, 
        n29425, n877, n950, n405, n29587, n329, n1023, n807, 
        n28036, n28614, n28613, n761, n518, n29424, n332, n29586, 
        n880, n445, n29423, n259_adj_3836, n29585, n372, n29422, 
        n1096, n186, n29584, n299, n29421, n953, n44, n113_adj_3837, 
        n402, n1026, n28035, n28034, n17, n9_adj_3838, n11_adj_3839, 
        n226, n29420, n40877, n40822, n28033, n44557, n42071, 
        n41464, n834, n44539, n153, n29419, n42051, n42045, n44533, 
        n27, n15, n13_adj_3841, n11_adj_3842, n41308, n21_adj_3843, 
        n19, n17_adj_3844, n9_adj_3845, n41333, n43, n16, n1099, 
        n41266, n8_adj_3846, n45, n24_adj_3847, n907, n28032;
    wire [10:0]n8064;
    
    wire n840, n29583, n28031, n475, n7_adj_3850, n5_adj_3851, n41382, 
        n767, n29582, n11_adj_3852, n80, n41997, n41987, n980, 
        n25_adj_3853, n23_adj_3854, n42683, n31, n29, n42257, n41_adj_3855, 
        n39, n45_adj_3856, n107, n37, n35, n33, n42769, n43_adj_3857, 
        n694, n29581, n29_adj_3858, n31_adj_3859, n38, n41483, n44526;
    wire [0:0]n6308;
    wire [21:0]n7855;
    
    wire n29418, n29417, n24250, n28030, n621, n29580, n28612, 
        n29416, n28029, n548, n29579, n29415, n37_adj_3861, n42031, 
        n44521, n23_adj_3862, n25_adj_3863, n12_adj_3864, n41406, 
        n44544, n28028, n10_adj_3866, n30, n35_adj_3867, n42301, 
        n29414, n28027, n33_adj_3868;
    wire [23:0]duty_23__N_3617;
    wire [23:0]\PID_CONTROLLER.err_23__N_3641 ;
    
    wire n11_adj_3869, n13_adj_3870, n15_adj_3871, n27_adj_3872, n29413, 
        n29578, n41423, n29412, n9_adj_3873, n44524, n17_adj_3874, 
        n42291, n44550, n19_adj_3875, n42691, n44515, n21_adj_3876, 
        n41232, n42837, n41184, n44512, n16_adj_3877, n41387, n24_adj_3878, 
        n29577, n29411, n6_adj_3879, n42470, n12_adj_3880, n30_adj_3881, 
        n29410, n42471, n41392, n8_adj_3882, n44510, n42361, n41262, 
        n41901, n41628;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3716 ;
    
    wire n3_adj_3883, n4_adj_3884, n42432, n41893, n42433, n12_adj_3885, 
        n42663, n41298, n42203, n10_adj_3886, n42765, n30_adj_3887, 
        n29409, n29576, n41302, n29408, n6_adj_3888, n42405, n42406, 
        n42709, n41640, n29407, n42843, n42844, n16_adj_3889, n24_adj_3890, 
        n39_adj_3891, n42819, n41124, n6_adj_3892, n42436, n8_adj_3893, 
        n41120, n42365, n41648, n4_adj_3894, n42437, n29406, n42401, 
        n41278, n29405, n29404, n42402, n41150, n42363, n29575, 
        n41638, n41_adj_3895, n41282, n29574, n10_adj_3896, n41145, 
        n42717, n41650, n28026, n42739, n42847, n41646, n42741, 
        n28025, n42848, n4_adj_3897, n42468, n42469, n42815, n41411, 
        n41126, n42699, n42582, n41630, n42833, n42834, n42826, 
        n41394, n42735, n41636, n41656, \PID_CONTROLLER.integral_23__N_3715 , 
        n42743, n42737, \PID_CONTROLLER.integral_23__N_3713 , duty_23__N_3764, 
        n29403;
    wire [11:0]n8050;
    
    wire n29573, n29572, n28024, n29402, n29571, n28023, n29570, 
        n29401, n29569, n29568, n40615, n29567, n28631, n29400, 
        n29399, n29398, n256_adj_3900, n29397, n29566, n29565, n28022, 
        n29396, n29395, n28021, n29564, n29394, n29393, n29563, 
        n28020, n29392, n28019, n29391, n29390;
    wire [12:0]n8035;
    
    wire n29562, n29561, n29389, n29560, n28018, n29388, n29387, 
        n29386, n29559, n29385, n28632, n28017, n29558, n29384, 
        n29557, n29383, n28016, n29556, n29382, n29381, n95, n26, 
        n168, n29380, n29555, n29379, n29378, n28015, n29554, 
        n29377, n241, n314, n150, n29376, n323, n29553, n8_adj_3904, 
        n77, n250, n29552, n28014, n387, n177, n29551, n28013, 
        n460, n35_adj_3907, n104, n533;
    wire [13:0]n8019;
    
    wire n1050, n29550, n977, n29549, n904, n29548, n606, n831, 
        n29547, n758, n29546, n685, n29545, n612, n29544, n28012, 
        n539, n29543, n28011, n28010, n466, n29542, n28009, n28008, 
        n28007, n393, n29541, n28006, n320, n29540, n28005, n247, 
        n29539, n28004, n174, n29538, n32, n101;
    wire [14:0]n8002;
    
    wire n1120, n29537, n1047, n29536, n974, n29535, n901, n29534, 
        n828, n29533, n755, n29532, n682, n29531, n28003, n609, 
        n29530, n536, n29529, n463, n29528, n390, n29527, n317, 
        n29526, n244, n29525, n171, n29524, n29_adj_3919, n98;
    wire [15:0]n7984;
    
    wire n29523, n1117, n29522, n1044, n29521, n971, n29520, n898, 
        n29519, n28002, n825, n29518, n752, n29517, n679, n29516, 
        n28001, n29515, n29514, n29513, n29512, n29511, n29510, 
        n29509;
    wire [16:0]n7965;
    
    wire n29508, n29507, n28000, n29506, n29505, n29504, n29503, 
        n29502, n29501, n29500, n29499, n29498;
    wire [47:0]n155;
    
    wire n457, n29497, n384, n29496, n311, n29495, n238, n29494, 
        n165, n29493, n23_adj_3921, n92;
    wire [17:0]n7945;
    
    wire n29492, n29491, n45_adj_3922, n29490, n1111, n29489, n21_adj_3923, 
        n19_adj_3924, n17_adj_3925, n9_adj_3926, n41069, n27_adj_3927, 
        n15_adj_3928, n13_adj_3929, n11_adj_3930, n41051, n33_adj_3931, 
        n12_adj_3932, n1038, n29488, n965, n29487, n10_adj_3933, 
        n35_adj_3934, n30_adj_3935, n892, n29486, n819, n29485, 
        n4_adj_3936;
    wire [3:0]n8431;
    
    wire n6_adj_3937;
    wire [4:0]n8424;
    
    wire n27690, n746, n29484, n673, n29483, n600, n29482, n527, 
        n29481, n454, n29480, n381, n29479, n308, n29478, n235, 
        n29477, n162, n29476, n27767;
    wire [1:0]n8442;
    
    wire n4_adj_3938;
    wire [2:0]n8437;
    
    wire n62, n131, n204, n4_adj_3939, n20_adj_3940, n89, n41111, 
        n41799, n41791, n25_adj_3941, n23_adj_3942, n42647, n31_adj_3943, 
        n29_adj_3944, n42173, n37_adj_3945, n42749, n43_adj_3946, 
        n16_adj_3947, n6_adj_3948, n42381, n42382, n8_adj_3949, n24_adj_3950, 
        n40965, n40955, n42367, n41658, n4_adj_3951, n42379, n42380, 
        n41024, n41016, n42383, n41660, n42810, n42811, n39_adj_3952, 
        n42748, n41_adj_3953, n40969, n42584, n41666, n42745;
    wire [18:0]n7924;
    
    wire n29475, n29474, n29473, n29472, n1108, n29471, n1035, 
        n29470, n962, n29469, n889, n29468, n816, n29467, n27975, 
        n743, n29466, n27974, n670, n29465, n27973, n597, n29464, 
        n524, n29463, n27972, n451, n29462, n27971, n378, n29461, 
        n305, n29460, n27970, n232, n29459;
    wire [5:0]n8416;
    
    wire n36379, n490, n29861, n417, n29860, n344, n29859, n271_adj_3955, 
        n29858, n198, n29857, n28634, n56, n125_adj_3956, n28633;
    wire [6:0]n8407;
    
    wire n560, n29856, n487, n29855, n414, n29854, n341, n29853, 
        n268_adj_3957, n29852, n195, n29851, n159, n29458, n53, 
        n122_adj_3958;
    wire [7:0]n8397;
    
    wire n630, n29850, n557, n29849, n484, n29848, n411, n29847, 
        n338, n29846, n27969, n265_adj_3959, n29845, n17_adj_3960, 
        n86, n192, n29844, n50, n119_adj_3961, n29457;
    wire [8:0]n8386;
    
    wire n700, n29843, n627, n29842, n554, n29841, n481, n29840, 
        n408, n29839, n335, n29838, n262_adj_3962, n29837, n189, 
        n29836, n47_adj_3963, n116_adj_3964, n27968;
    wire [9:0]n8374;
    
    wire n770_adj_3965, n29835, n697_adj_3966, n29834, n624_adj_3967, 
        n29833, n551_adj_3968, n29832, n478_adj_3969, n29831, n29456, 
        n405_adj_3970, n29830;
    wire [23:0]n1_adj_4255;
    
    wire n28165, n28164, n332_adj_3973, n29829, n259_adj_3974, n29828, 
        n186_adj_3975, n29827, n44_adj_3976, n113_adj_3977;
    wire [10:0]n8361;
    
    wire n840_adj_3978, n29826, n767_adj_3979, n29825, n694_adj_3980, 
        n29824, n28163, n28162, n28161, n621_adj_3984, n29823, n548_adj_3985, 
        n29822, n475_adj_3986, n29821, n402_adj_3987, n29820, n29455, 
        n28160, n329_adj_3989, n29819, n29454, n256_adj_3990, n29818, 
        n183_adj_3991, n29817, n41_adj_3992, n110_adj_3993, n28159, 
        n28158;
    wire [11:0]n8347;
    
    wire n910_adj_3996, n29816, n28157, n837_adj_3998, n29815, n764_adj_3999, 
        n29814, n28156, n691_adj_4001, n29813, n618_adj_4002, n29812, 
        n545_adj_4003, n29811, n472_adj_4004, n29810, n399_adj_4005, 
        n29809, n326_adj_4006, n29808, n253_adj_4007, n29807, n180_adj_4008, 
        n29806, n38_adj_4009, n107_adj_4010;
    wire [12:0]n8332;
    
    wire n980_adj_4011, n29805, n907_adj_4012, n29804, n27967, n834_adj_4013, 
        n29803, n28155, n761_adj_4015, n29802, n688_adj_4016, n29801, 
        n28154, n615_adj_4018, n29800, n542_adj_4019, n29799, n28153, 
        n469_adj_4021, n29798, n28152, n396_adj_4023, n29797, n28151, 
        n323_adj_4025, n29796, n250_adj_4026, n29795, n28150, n177_adj_4028, 
        n29794, n28149, n35_adj_4030, n104_adj_4031, n28148, n28147;
    wire [13:0]n8316;
    
    wire n1050_adj_4034, n29793, n977_adj_4035, n29792, n28146, n904_adj_4037, 
        n29791, n831_adj_4038, n29790, n28145, n758_adj_4040, n29789, 
        n685_adj_4041, n29788, n612_adj_4042, n29787, n28144, n28143, 
        n539_adj_4045, n29786, n466_adj_4046, n29785, n393_adj_4048, 
        n29784, n320_adj_4049, n29783, n247_adj_4050, n29782, n174_adj_4051, 
        n29781, n32_adj_4052, n101_adj_4053;
    wire [14:0]n8299;
    
    wire n1120_adj_4054, n29780, n1047_adj_4055, n29779, n974_adj_4056, 
        n29778, n901_adj_4057, n29777, n828_adj_4058, n29776, n755_adj_4059, 
        n29775, n27966, n682_adj_4060, n29774, n609_adj_4061, n29773, 
        n29453, n536_adj_4062, n29772, n463_adj_4063, n29771, n390_adj_4064, 
        n29770, n317_adj_4065, n29769, n244_adj_4066, n29768, n171_adj_4067, 
        n29767, n27965, n29_adj_4068, n98_adj_4069;
    wire [15:0]n8281;
    
    wire n29766, n1117_adj_4070, n29765, n1044_adj_4071, n29764, n27964, 
        n971_adj_4072, n29763, n898_adj_4073, n29762, n825_adj_4074, 
        n29761, n752_adj_4075, n29760, n679_adj_4076, n29759, n27963, 
        n606_adj_4077, n29758, n533_adj_4078, n29757, n460_adj_4079, 
        n29756, n387_adj_4080, n29755, n314_adj_4081, n29754, n241_adj_4082, 
        n29753, n168_adj_4083, n29752, n1105, n29452, n26_adj_4084, 
        n95_adj_4085;
    wire [16:0]n8262;
    
    wire n29751, n29750, n27962, n1114_adj_4086, n29749, n1041_adj_4087, 
        n29748, n968_adj_4088, n29747, n895_adj_4089, n29746, n822_adj_4090, 
        n29745, n749_adj_4091, n29744, n676_adj_4092, n29743, n603_adj_4093, 
        n29742, n530_adj_4094, n29741, n457_adj_4095, n29740, n384_adj_4096, 
        n29739, n311_adj_4097, n29738, n27961, n238_adj_4098, n29737, 
        n165_adj_4099, n29736, n23_adj_4100, n92_adj_4101;
    wire [17:0]n8242;
    
    wire n29735, n29734, n29733, n1111_adj_4102, n29732, n1038_adj_4103, 
        n29731, n27960, n965_adj_4104, n29730, n892_adj_4105, n29729, 
        n819_adj_4106, n29728, n1032, n29451, n746_adj_4107, n29727, 
        n673_adj_4108, n29726, n600_adj_4109, n29725, n527_adj_4110, 
        n29724, n454_adj_4111, n29723, n381_adj_4112, n29722, n308_adj_4113, 
        n29721, n235_adj_4114, n29720, n162_adj_4115, n29719, n20_adj_4116, 
        n89_adj_4117;
    wire [18:0]n8221;
    
    wire n29718, n29717, n29716, n29715, n27959, n1108_adj_4118, 
        n29714, n1035_adj_4119, n29713, n962_adj_4120, n29712, n889_adj_4121, 
        n29711, n816_adj_4122, n29710, n743_adj_4123, n29709, n670_adj_4124, 
        n29708, n597_adj_4125, n29707, n27958, n27563;
    wire [2:0]n8140;
    
    wire n4_adj_4126;
    wire [3:0]n8134;
    
    wire n959, n29450, n886, n29449, n524_adj_4127, n29706, n451_adj_4128, 
        n29705, n378_adj_4129, n29704, n305_adj_4130, n29703, n232_adj_4131, 
        n29702, n159_adj_4132, n29701, n17_adj_4133, n86_adj_4134;
    wire [19:0]n8199;
    
    wire n29700, n29699, n27957, n29698, n29697, n29696, n27597;
    wire [1:0]n8145;
    
    wire n4_adj_4135, n1105_adj_4136, n29695, n1032_adj_4137, n29694, 
        n959_adj_4138, n29693, n886_adj_4139, n29692, n813, n29691, 
        n740, n29690, n667, n29689, n594, n29688, n521, n29687, 
        n448, n29686, n375, n29685, n813_adj_4140, n29448, n302, 
        n29684, n229, n29683, n156, n29682, n14_adj_4141, n83;
    wire [20:0]n8176;
    
    wire n29681, n29680, n29679, n29678, n29677, n29676, n1102_adj_4142, 
        n29675, n1029_adj_4143, n29674, n956_adj_4144, n29673, n883_adj_4145, 
        n29672, n740_adj_4146, n29447, n810_adj_4147, n29671, n737_adj_4148, 
        n29670, n664_adj_4149, n29669, n591_adj_4150, n29668, n518_adj_4151, 
        n29667, n445_adj_4152, n29666, n372_adj_4153, n29665, n299_adj_4154, 
        n29664, n226_adj_4155, n29663, n153_adj_4156, n29662, n11_adj_4157, 
        n80_adj_4158, n40677;
    wire [21:0]n8152;
    
    wire n29661, n667_adj_4159, n29446, n29660, n29659, n29658, 
        n29657, n594_adj_4161, n29445, n29656, n29655, n29654, n1096_adj_4163, 
        n29653, n1023_adj_4165, n29652, n950_adj_4166, n29651, n877_adj_4167, 
        n29650, n804_adj_4169, n29649, n731_adj_4170, n29648, n658_adj_4171, 
        n29647, n585_adj_4173, n29646, n521_adj_4174, n29444, n512_adj_4175, 
        n29645, n439_adj_4176, n29644, n366_adj_4178, n29643, n293_adj_4179, 
        n29642, n220_adj_4180, n29641, n147_adj_4181, n29640, n5_adj_4182, 
        n74_adj_4183, n29639, n29638, n29637, n29636, n29635, n29634, 
        n29633, n1099_adj_4184, n29632, n1026_adj_4185, n29631, n953_adj_4186, 
        n29630, n448_adj_4187, n29443, n880_adj_4188, n29629, n27956, 
        n807_adj_4189, n29628, n375_adj_4190, n29442, n734_adj_4191, 
        n29627, n661_adj_4192, n29626, n588_adj_4193, n29625, n515_adj_4194, 
        n29624, n442_adj_4195, n29623, n302_adj_4196, n29441, n229_adj_4197, 
        n29440, n369_adj_4198, n29622, n296_adj_4199, n29621, n223_adj_4200, 
        n29620, n150_adj_4201, n29619, n8_adj_4202, n77_adj_4203;
    wire [5:0]n8119;
    
    wire n37305, n490_adj_4204, n29618;
    wire [4:0]n8127;
    
    wire n417_adj_4205, n29617, n344_adj_4206, n29616, n271_adj_4207, 
        n29615, n198_adj_4208, n29614, n56_adj_4209, n125_adj_4210;
    wire [6:0]n8110;
    
    wire n560_adj_4211, n29613, n487_adj_4212, n29612, n414_adj_4213, 
        n29611, n156_adj_4214, n29439, n341_adj_4215, n29610, n268_adj_4216, 
        n29609, n14_adj_4217, n83_adj_4218, n195_adj_4219, n29608, 
        n53_adj_4220, n122_adj_4221;
    wire [7:0]n8100;
    
    wire n630_adj_4222, n29607, n557_adj_4223, n29606, n484_adj_4224, 
        n29605, n411_adj_4225, n29604, n338_adj_4226, n29603, n265_adj_4227, 
        n29602, n192_adj_4228, n29601, n50_adj_4229, n119_adj_4230, 
        n700_adj_4231, n29600, n627_adj_4232, n29599, n554_adj_4233, 
        n29598, n481_adj_4234, n29597, n408_adj_4235, n29596, n335_adj_4236, 
        n29595, n262_adj_4237, n29594, n189_adj_4238, n4_adj_4239, 
        n6_adj_4240, n12_adj_4241, n6_adj_4242, n11_adj_4243, n8_adj_4244, 
        n27622, n18_adj_4245, n13_adj_4246, n27520, n12_adj_4247, 
        n8_adj_4248, n11_adj_4249, n6_adj_4250, n27792, n18_adj_4251, 
        n13_adj_4252;
    
    SB_LUT4 add_3771_22_lut (.I0(GND_net), .I1(n7902[19]), .I2(GND_net), 
            .I3(n29438), .O(n7879[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_639_4_lut (.I0(GND_net), .I1(n3048[2]), .I2(n3073[2]), 
            .I3(n27954), .O(duty_23__N_3740[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_20  (.CI(n28629), .I0(\PID_CONTROLLER.err [18]), 
            .I1(\PID_CONTROLLER.integral [18]), .CO(n28630));
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_19_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(n28628), .O(n1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_19_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_639_4 (.CI(n27954), .I0(n3048[2]), .I1(n3073[2]), .CO(n27955));
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_19  (.CI(n28628), .I0(\PID_CONTROLLER.err [17]), 
            .I1(\PID_CONTROLLER.integral [17]), .CO(n28629));
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(duty[23]), .I1(GND_net), .I2(n1_adj_4253[23]), 
            .I3(n28045), .O(n47)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_639_3_lut (.I0(GND_net), .I1(n3048[1]), .I2(n3073[1]), 
            .I3(n27953), .O(duty_23__N_3740[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3771_21_lut (.I0(GND_net), .I1(n7902[18]), .I2(GND_net), 
            .I3(n29437), .O(n7879[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[22]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3783_2_lut (.I0(GND_net), .I1(n47_adj_3826), .I2(n116), 
            .I3(GND_net), .O(n8089[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3783_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_639_3 (.CI(n27953), .I0(n3048[1]), .I1(n3073[1]), .CO(n27954));
    SB_CARRY add_3783_2 (.CI(GND_net), .I0(n47_adj_3826), .I1(n116), .CO(n29593));
    SB_CARRY add_3771_21 (.CI(n29437), .I0(n7902[18]), .I1(GND_net), .CO(n29438));
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_18_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(n28627), .O(n1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_18_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3771_20_lut (.I0(GND_net), .I1(n7902[17]), .I2(GND_net), 
            .I3(n29436), .O(n7879[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_639_2_lut (.I0(GND_net), .I1(n3048[0]), .I2(n3073[0]), 
            .I3(GND_net), .O(duty_23__N_3740[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_639_2 (.CI(GND_net), .I0(n3048[0]), .I1(n3073[0]), .CO(n27953));
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3782_11_lut (.I0(GND_net), .I1(n8089[8]), .I2(n770), .I3(n29592), 
            .O(n8077[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3782_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3771_20 (.CI(n29436), .I0(n7902[17]), .I1(GND_net), .CO(n29437));
    SB_LUT4 add_3771_19_lut (.I0(GND_net), .I1(n7902[16]), .I2(GND_net), 
            .I3(n29435), .O(n7879[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_18  (.CI(n28627), .I0(\PID_CONTROLLER.err [16]), 
            .I1(\PID_CONTROLLER.integral [16]), .CO(n28628));
    SB_CARRY add_3771_19 (.CI(n29435), .I0(n7902[16]), .I1(GND_net), .CO(n29436));
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_17_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [15]), 
            .I2(\PID_CONTROLLER.integral [15]), .I3(n28626), .O(n1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_17_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[22]), 
            .I3(n28044), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_17  (.CI(n28626), .I0(\PID_CONTROLLER.err [15]), 
            .I1(\PID_CONTROLLER.integral [15]), .CO(n28627));
    SB_LUT4 add_3782_10_lut (.I0(GND_net), .I1(n8089[7]), .I2(n697), .I3(n29591), 
            .O(n8077[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3782_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3771_18_lut (.I0(GND_net), .I1(n7902[15]), .I2(GND_net), 
            .I3(n29434), .O(n7879[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_16_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [14]), 
            .I2(\PID_CONTROLLER.integral [14]), .I3(n28625), .O(n1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_16_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3771_18 (.CI(n29434), .I0(n7902[15]), .I1(GND_net), .CO(n29435));
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_16  (.CI(n28625), .I0(\PID_CONTROLLER.err [14]), 
            .I1(\PID_CONTROLLER.integral [14]), .CO(n28626));
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_15_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [13]), 
            .I2(\PID_CONTROLLER.integral [13]), .I3(n28624), .O(n1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_15_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3782_10 (.CI(n29591), .I0(n8089[7]), .I1(n697), .CO(n29592));
    SB_LUT4 add_3771_17_lut (.I0(GND_net), .I1(n7902[14]), .I2(GND_net), 
            .I3(n29433), .O(n7879[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3771_17 (.CI(n29433), .I0(n7902[14]), .I1(GND_net), .CO(n29434));
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_15  (.CI(n28624), .I0(\PID_CONTROLLER.err [13]), 
            .I1(\PID_CONTROLLER.integral [13]), .CO(n28625));
    SB_LUT4 add_3782_9_lut (.I0(GND_net), .I1(n8089[6]), .I2(n624), .I3(n29590), 
            .O(n8077[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3782_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3771_16_lut (.I0(GND_net), .I1(n7902[13]), .I2(n1102), 
            .I3(n29432), .O(n7879[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_14_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [12]), 
            .I2(\PID_CONTROLLER.integral [12]), .I3(n28623), .O(n1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_14_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3771_16 (.CI(n29432), .I0(n7902[13]), .I1(n1102), .CO(n29433));
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_14  (.CI(n28623), .I0(\PID_CONTROLLER.err [12]), 
            .I1(\PID_CONTROLLER.integral [12]), .CO(n28624));
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_13_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [11]), 
            .I2(\PID_CONTROLLER.integral [11]), .I3(n28622), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_13_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_13  (.CI(n28622), .I0(\PID_CONTROLLER.err [11]), 
            .I1(\PID_CONTROLLER.integral [11]), .CO(n28623));
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_12_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [10]), 
            .I2(\PID_CONTROLLER.integral [10]), .I3(n28621), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_12_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3782_9 (.CI(n29590), .I0(n8089[6]), .I1(n624), .CO(n29591));
    SB_LUT4 add_3771_15_lut (.I0(GND_net), .I1(n7902[12]), .I2(n1029), 
            .I3(n29431), .O(n7879[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_12  (.CI(n28621), .I0(\PID_CONTROLLER.err [10]), 
            .I1(\PID_CONTROLLER.integral [10]), .CO(n28622));
    SB_CARRY add_3771_15 (.CI(n29431), .I0(n7902[12]), .I1(n1029), .CO(n29432));
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_11_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [9]), 
            .I2(\PID_CONTROLLER.integral [9]), .I3(n28620), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_11_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_11  (.CI(n28620), .I0(\PID_CONTROLLER.err [9]), 
            .I1(\PID_CONTROLLER.integral [9]), .CO(n28621));
    SB_CARRY unary_minus_16_add_3_24 (.CI(n28044), .I0(GND_net), .I1(n1_adj_4253[22]), 
            .CO(n28045));
    SB_LUT4 add_3782_8_lut (.I0(GND_net), .I1(n8089[5]), .I2(n551), .I3(n29589), 
            .O(n8077[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3782_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3771_14_lut (.I0(GND_net), .I1(n7902[11]), .I2(n956), 
            .I3(n29430), .O(n7879[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_10_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(n28619), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_10_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3771_14 (.CI(n29430), .I0(n7902[11]), .I1(n956), .CO(n29431));
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[21]), 
            .I3(n28043), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_10  (.CI(n28619), .I0(\PID_CONTROLLER.err [8]), 
            .I1(\PID_CONTROLLER.integral [8]), .CO(n28620));
    SB_CARRY unary_minus_16_add_3_23 (.CI(n28043), .I0(GND_net), .I1(n1_adj_4253[21]), 
            .CO(n28044));
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_9_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [7]), 
            .I2(\PID_CONTROLLER.integral [7]), .I3(n28618), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_9_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[20]), 
            .I3(n28042), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3782_8 (.CI(n29589), .I0(n8089[5]), .I1(n551), .CO(n29590));
    SB_LUT4 add_3771_13_lut (.I0(GND_net), .I1(n7902[10]), .I2(n883), 
            .I3(n29429), .O(n7879[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3771_13 (.CI(n29429), .I0(n7902[10]), .I1(n883), .CO(n29430));
    SB_CARRY unary_minus_16_add_3_22 (.CI(n28042), .I0(GND_net), .I1(n1_adj_4253[20]), 
            .CO(n28043));
    SB_LUT4 add_3782_7_lut (.I0(GND_net), .I1(n8089[4]), .I2(n478), .I3(n29588), 
            .O(n8077[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3782_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3771_12_lut (.I0(GND_net), .I1(n7902[9]), .I2(n810), .I3(n29428), 
            .O(n7879[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[19]), 
            .I3(n28041), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_9  (.CI(n28618), .I0(\PID_CONTROLLER.err [7]), 
            .I1(\PID_CONTROLLER.integral [7]), .CO(n28619));
    SB_CARRY add_3771_12 (.CI(n29428), .I0(n7902[9]), .I1(n810), .CO(n29429));
    SB_CARRY unary_minus_16_add_3_21 (.CI(n28041), .I0(GND_net), .I1(n1_adj_4253[19]), 
            .CO(n28042));
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_8_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(n28617), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_8_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[18]), 
            .I3(n28040), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_8  (.CI(n28617), .I0(\PID_CONTROLLER.err [6]), 
            .I1(\PID_CONTROLLER.integral [6]), .CO(n28618));
    SB_CARRY unary_minus_16_add_3_20 (.CI(n28040), .I0(GND_net), .I1(n1_adj_4253[18]), 
            .CO(n28041));
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[23]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[16]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[17]), 
            .I3(n28039), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_7_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [5]), 
            .I2(\PID_CONTROLLER.integral [5]), .I3(n28616), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_7_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_19 (.CI(n28039), .I0(GND_net), .I1(n1_adj_4253[17]), 
            .CO(n28040));
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_7  (.CI(n28616), .I0(\PID_CONTROLLER.err [5]), 
            .I1(\PID_CONTROLLER.integral [5]), .CO(n28617));
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[16]), 
            .I3(n28038), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3771_11_lut (.I0(GND_net), .I1(n7902[8]), .I2(n737), .I3(n29427), 
            .O(n7879[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[0]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3771_11 (.CI(n29427), .I0(n7902[8]), .I1(n737), .CO(n29428));
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3771_10_lut (.I0(GND_net), .I1(n7902[7]), .I2(n664), .I3(n29426), 
            .O(n7879[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_18 (.CI(n28038), .I0(GND_net), .I1(n1_adj_4253[16]), 
            .CO(n28039));
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[15]), 
            .I3(n28037), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[1]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[17]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[2]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_6_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [4]), 
            .I2(\PID_CONTROLLER.integral [4]), .I3(n28615), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_6_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_6  (.CI(n28615), .I0(\PID_CONTROLLER.err [4]), 
            .I1(\PID_CONTROLLER.integral [4]), .CO(n28616));
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[3]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_3833));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[4]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[18]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3771_10 (.CI(n29426), .I0(n7902[7]), .I1(n664), .CO(n29427));
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3782_7 (.CI(n29588), .I0(n8089[4]), .I1(n478), .CO(n29589));
    SB_LUT4 add_3771_9_lut (.I0(GND_net), .I1(n7902[6]), .I2(n591), .I3(n29425), 
            .O(n7879[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[0]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3782_6_lut (.I0(GND_net), .I1(n8089[3]), .I2(n405), .I3(n29587), 
            .O(n8077[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3782_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_17 (.CI(n28037), .I0(GND_net), .I1(n1_adj_4253[15]), 
            .CO(n28038));
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[14]), 
            .I3(n28036), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_16 (.CI(n28036), .I0(GND_net), .I1(n1_adj_4253[14]), 
            .CO(n28037));
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_5_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(n28614), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_5_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_5  (.CI(n28614), .I0(\PID_CONTROLLER.err [3]), 
            .I1(\PID_CONTROLLER.integral [3]), .CO(n28615));
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_4_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [2]), 
            .I2(\PID_CONTROLLER.integral [2]), .I3(n28613), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_4_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3782_6 (.CI(n29587), .I0(n8089[3]), .I1(n405), .CO(n29588));
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3771_9 (.CI(n29425), .I0(n7902[6]), .I1(n591), .CO(n29426));
    SB_LUT4 add_3771_8_lut (.I0(GND_net), .I1(n7902[5]), .I2(n518), .I3(n29424), 
            .O(n7879[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3782_5_lut (.I0(GND_net), .I1(n8089[2]), .I2(n332), .I3(n29586), 
            .O(n8077[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3782_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3782_5 (.CI(n29586), .I0(n8089[2]), .I1(n332), .CO(n29587));
    SB_CARRY add_3771_8 (.CI(n29424), .I0(n7902[5]), .I1(n518), .CO(n29425));
    SB_LUT4 add_3771_7_lut (.I0(GND_net), .I1(n7902[4]), .I2(n445), .I3(n29423), 
            .O(n7879[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3782_4_lut (.I0(GND_net), .I1(n8089[1]), .I2(n259_adj_3836), 
            .I3(n29585), .O(n8077[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3782_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3771_7 (.CI(n29423), .I0(n7902[4]), .I1(n445), .CO(n29424));
    SB_LUT4 add_3771_6_lut (.I0(GND_net), .I1(n7902[3]), .I2(n372), .I3(n29422), 
            .O(n7879[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3782_4 (.CI(n29585), .I0(n8089[1]), .I1(n259_adj_3836), 
            .CO(n29586));
    SB_LUT4 add_3782_3_lut (.I0(GND_net), .I1(n8089[0]), .I2(n186), .I3(n29584), 
            .O(n8077[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3782_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3771_6 (.CI(n29422), .I0(n7902[3]), .I1(n372), .CO(n29423));
    SB_LUT4 add_3771_5_lut (.I0(GND_net), .I1(n7902[2]), .I2(n299), .I3(n29421), 
            .O(n7879[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3782_3 (.CI(n29584), .I0(n8089[0]), .I1(n186), .CO(n29585));
    SB_CARRY add_3771_5 (.CI(n29421), .I0(n7902[2]), .I1(n299), .CO(n29422));
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3782_2_lut (.I0(GND_net), .I1(n44), .I2(n113_adj_3837), 
            .I3(GND_net), .O(n8077[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3782_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[13]), 
            .I3(n28035), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n28035), .I0(GND_net), .I1(n1_adj_4253[13]), 
            .CO(n28036));
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[12]), 
            .I3(n28034), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_3838));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_3839));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n28034), .I0(GND_net), .I1(n1_adj_4253[12]), 
            .CO(n28035));
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[19]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3782_2 (.CI(GND_net), .I0(n44), .I1(n113_adj_3837), .CO(n29584));
    SB_LUT4 add_3771_4_lut (.I0(GND_net), .I1(n7902[1]), .I2(n226), .I3(n29420), 
            .O(n7879[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34031_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n40877));
    defparam i34031_4_lut.LUT_INIT = 16'h7bde;
    SB_CARRY add_3771_4 (.CI(n29420), .I0(n7902[1]), .I1(n226), .CO(n29421));
    SB_LUT4 i33976_3_lut (.I0(n11_adj_3839), .I1(n9_adj_3838), .I2(n40877), 
            .I3(GND_net), .O(n40822));
    defparam i33976_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[11]), 
            .I3(n28033), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_443_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n44557));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_443_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35224_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n44557), 
            .I2(IntegralLimit[7]), .I3(n40822), .O(n42071));
    defparam i35224_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i34617_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17), .I2(IntegralLimit[9]), 
            .I3(n42071), .O(n41464));
    defparam i34617_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_425_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n44539));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_425_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3771_3_lut (.I0(GND_net), .I1(n7902[0]), .I2(n153), .I3(n29419), 
            .O(n7879[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35204_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17), .I2(IntegralLimit[9]), 
            .I3(n9_adj_3838), .O(n42051));
    defparam i35204_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i35198_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n44539), 
            .I2(IntegralLimit[11]), .I3(n42051), .O(n42045));
    defparam i35198_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_419_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n44533));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_419_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34461_4_lut (.I0(n27), .I1(n15), .I2(n13_adj_3841), .I3(n11_adj_3842), 
            .O(n41308));
    defparam i34461_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34486_4_lut (.I0(n21_adj_3843), .I1(n19), .I2(n17_adj_3844), 
            .I3(n9_adj_3845), .O(n41333));
    defparam i34486_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43), .I3(GND_net), 
            .O(n16));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34419_2_lut (.I0(n43), .I1(n19), .I2(GND_net), .I3(GND_net), 
            .O(n41266));
    defparam i34419_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_3844), .I3(GND_net), 
            .O(n8_adj_3846));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n45), .I3(GND_net), .O(n24_adj_3847));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n28033), .I0(GND_net), .I1(n1_adj_4253[11]), 
            .CO(n28034));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[10]), 
            .I3(n28032), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n28032), .I0(GND_net), .I1(n1_adj_4253[10]), 
            .CO(n28033));
    SB_LUT4 add_3781_12_lut (.I0(GND_net), .I1(n8077[9]), .I2(n840), .I3(n29583), 
            .O(n8064[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3781_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[9]), 
            .I3(n28031), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34535_2_lut (.I0(n7_adj_3850), .I1(n5_adj_3851), .I2(GND_net), 
            .I3(GND_net), .O(n41382));
    defparam i34535_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 add_3781_11_lut (.I0(GND_net), .I1(n8077[8]), .I2(n767), .I3(n29582), 
            .O(n8064[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3781_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3781_11 (.CI(n29582), .I0(n8077[8]), .I1(n767), .CO(n29583));
    SB_CARRY add_3771_3 (.CI(n29419), .I0(n7902[0]), .I1(n153), .CO(n29420));
    SB_LUT4 add_3771_2_lut (.I0(GND_net), .I1(n11_adj_3852), .I2(n80), 
            .I3(GND_net), .O(n7879[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3771_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35150_4_lut (.I0(n13_adj_3841), .I1(n11_adj_3842), .I2(n9_adj_3845), 
            .I3(n41382), .O(n41997));
    defparam i35150_4_lut.LUT_INIT = 16'heeef;
    SB_CARRY add_3771_2 (.CI(GND_net), .I0(n11_adj_3852), .I1(n80), .CO(n29419));
    SB_LUT4 i35140_4_lut (.I0(n19), .I1(n17_adj_3844), .I2(n15), .I3(n41997), 
            .O(n41987));
    defparam i35140_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35836_4_lut (.I0(n25_adj_3853), .I1(n23_adj_3854), .I2(n21_adj_3843), 
            .I3(n41987), .O(n42683));
    defparam i35836_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35410_4_lut (.I0(n31), .I1(n29), .I2(n27), .I3(n42683), 
            .O(n42257));
    defparam i35410_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 duty_23__I_0_i41_2_lut (.I0(PWMLimit[20]), .I1(duty[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_3855));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i39_2_lut (.I0(PWMLimit[19]), .I1(duty[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i45_2_lut (.I0(PWMLimit[22]), .I1(duty[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_3856));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35922_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n42257), 
            .O(n42769));
    defparam i35922_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n28031), .I0(GND_net), .I1(n1_adj_4253[9]), 
            .CO(n28032));
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_4  (.CI(n28613), .I0(\PID_CONTROLLER.err [2]), 
            .I1(\PID_CONTROLLER.integral [2]), .CO(n28614));
    SB_LUT4 duty_23__I_0_i43_2_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_3857));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 add_3781_10_lut (.I0(GND_net), .I1(n8077[7]), .I2(n694), .I3(n29581), 
            .O(n8064[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3781_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i29_2_lut (.I0(PWMLimit[14]), .I1(duty[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_3858));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i31_2_lut (.I0(PWMLimit[15]), .I1(duty[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_3859));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i34636_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n44557), 
            .I2(IntegralLimit[7]), .I3(n11_adj_3839), .O(n41483));
    defparam i34636_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_412_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n44526));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_412_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3781_10 (.CI(n29581), .I0(n8077[7]), .I1(n694), .CO(n29582));
    SB_LUT4 mult_10_add_1225_24_lut (.I0(\PID_CONTROLLER.err [23]), .I1(n7855[21]), 
            .I2(GND_net), .I3(n29418), .O(n6308[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(n24250), .I1(n7855[20]), .I2(GND_net), 
            .I3(n29417), .O(n3048[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[8]), 
            .I3(n28030), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3781_9_lut (.I0(GND_net), .I1(n8077[6]), .I2(n621), .I3(n29580), 
            .O(n8064[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3781_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_23 (.CI(n29417), .I0(n7855[20]), .I1(GND_net), 
            .CO(n29418));
    SB_CARRY unary_minus_16_add_3_10 (.CI(n28030), .I0(GND_net), .I1(n1_adj_4253[8]), 
            .CO(n28031));
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_3_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [1]), 
            .I2(\PID_CONTROLLER.integral [1]), .I3(n28612), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_3_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_22_lut (.I0(n24250), .I1(n7855[19]), .I2(GND_net), 
            .I3(n29416), .O(n3048[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[7]), 
            .I3(n28029), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3781_9 (.CI(n29580), .I0(n8077[6]), .I1(n621), .CO(n29581));
    SB_CARRY mult_10_add_1225_22 (.CI(n29416), .I0(n7855[19]), .I1(GND_net), 
            .CO(n29417));
    SB_LUT4 add_3781_8_lut (.I0(GND_net), .I1(n8077[5]), .I2(n548), .I3(n29579), 
            .O(n8064[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3781_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n28029), .I0(GND_net), .I1(n1_adj_4253[7]), 
            .CO(n28030));
    SB_LUT4 mult_10_add_1225_21_lut (.I0(n24250), .I1(n7855[18]), .I2(GND_net), 
            .I3(n29415), .O(n3048[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 duty_23__I_0_i37_2_lut (.I0(PWMLimit[18]), .I1(duty[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_3861));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i37_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_3781_8 (.CI(n29579), .I0(n8077[5]), .I1(n548), .CO(n29580));
    SB_LUT4 i35184_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n44526), 
            .I2(IntegralLimit[14]), .I3(n41483), .O(n42031));
    defparam i35184_4_lut.LUT_INIT = 16'hdeff;
    SB_CARRY mult_10_add_1225_21 (.CI(n29415), .I0(n7855[18]), .I1(GND_net), 
            .CO(n29416));
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_407_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n44521));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_407_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i23_2_lut (.I0(PWMLimit[11]), .I1(duty[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_3862));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i25_2_lut (.I0(PWMLimit[12]), .I1(duty[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_3863));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_3864));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34559_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n41406));
    defparam i34559_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_430_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n44544));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_430_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[6]), 
            .I3(n28028), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_3866));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_3864), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i35_2_lut (.I0(PWMLimit[17]), .I1(duty[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_3867));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35454_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n44539), 
            .I2(IntegralLimit[11]), .I3(n41464), .O(n42301));
    defparam i35454_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_10_add_1225_20_lut (.I0(n24250), .I1(n7855[17]), .I2(GND_net), 
            .I3(n29414), .O(n3048[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n28028), .I0(GND_net), .I1(n1_adj_4253[6]), 
            .CO(n28029));
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[5]), 
            .I3(n28027), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_3  (.CI(n28612), .I0(\PID_CONTROLLER.err [1]), 
            .I1(\PID_CONTROLLER.integral [1]), .CO(n28613));
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_2_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [0]), 
            .I2(\PID_CONTROLLER.integral [0]), .I3(GND_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_2_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_2  (.CI(GND_net), .I0(\PID_CONTROLLER.err [0]), 
            .I1(\PID_CONTROLLER.integral [0]), .CO(n28612));
    SB_CARRY mult_10_add_1225_20 (.CI(n29414), .I0(n7855[17]), .I1(GND_net), 
            .CO(n29415));
    SB_LUT4 duty_23__I_0_i33_2_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_3868));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i33_2_lut.LUT_INIT = 16'h6666;
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3617[0]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i0  (.Q(\PID_CONTROLLER.err [0]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [0]));   // verilog/motorControl.v(37[14] 56[8])
    SB_LUT4 duty_23__I_0_i11_2_lut (.I0(PWMLimit[5]), .I1(duty[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_3869));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i13_2_lut (.I0(PWMLimit[6]), .I1(duty[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_3870));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i15_2_lut (.I0(PWMLimit[7]), .I1(duty[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_3871));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i27_2_lut (.I0(PWMLimit[13]), .I1(duty[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_3872));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_add_1225_19_lut (.I0(n24250), .I1(n7855[16]), .I2(GND_net), 
            .I3(n29413), .O(n3048[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_19 (.CI(n29413), .I0(n7855[16]), .I1(GND_net), 
            .CO(n29414));
    SB_LUT4 add_3781_7_lut (.I0(GND_net), .I1(n8077[4]), .I2(n475), .I3(n29578), 
            .O(n8064[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3781_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34576_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n44533), 
            .I2(IntegralLimit[13]), .I3(n42301), .O(n41423));
    defparam i34576_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_10_add_1225_18_lut (.I0(n24250), .I1(n7855[15]), .I2(GND_net), 
            .I3(n29412), .O(n3048[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3781_7 (.CI(n29578), .I0(n8077[4]), .I1(n475), .CO(n29579));
    SB_CARRY mult_10_add_1225_18 (.CI(n29412), .I0(n7855[15]), .I1(GND_net), 
            .CO(n29413));
    SB_LUT4 duty_23__I_0_i9_2_lut (.I0(PWMLimit[4]), .I1(duty[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_3873));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_410_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n44524));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_410_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i17_2_lut (.I0(PWMLimit[8]), .I1(duty[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_3874));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35444_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n44524), 
            .I2(IntegralLimit[15]), .I3(n41423), .O(n42291));
    defparam i35444_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_436_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n44550));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_436_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i19_2_lut (.I0(PWMLimit[9]), .I1(duty[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_3875));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35844_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n44550), 
            .I2(IntegralLimit[17]), .I3(n42291), .O(n42691));
    defparam i35844_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_401_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n44515));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_401_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_0_i21_2_lut (.I0(PWMLimit[10]), .I1(duty[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_3876));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34385_4_lut (.I0(n21_adj_3876), .I1(n19_adj_3875), .I2(n17_adj_3874), 
            .I3(n9_adj_3873), .O(n41232));
    defparam i34385_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35990_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n44515), 
            .I2(IntegralLimit[19]), .I3(n42691), .O(n42837));
    defparam i35990_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i34337_4_lut (.I0(n27_adj_3872), .I1(n15_adj_3871), .I2(n13_adj_3870), 
            .I3(n11_adj_3869), .O(n41184));
    defparam i34337_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_398_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n44512));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_398_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_3877));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34540_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n41387));
    defparam i34540_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_3877), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_3878));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_3781_6_lut (.I0(GND_net), .I1(n8077[3]), .I2(n402), .I3(n29577), 
            .O(n8064[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3781_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_17_lut (.I0(n24250), .I1(n7855[14]), .I2(GND_net), 
            .I3(n29411), .O(n3048[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_3879));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35623_3_lut (.I0(n6_adj_3879), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n42470));   // verilog/motorControl.v(39[10:34])
    defparam i35623_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY add_3781_6 (.CI(n29577), .I0(n8077[3]), .I1(n402), .CO(n29578));
    SB_LUT4 duty_23__I_0_i30_3_lut (.I0(n12_adj_3880), .I1(duty[17]), .I2(n35_adj_3867), 
            .I3(GND_net), .O(n30_adj_3881));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_10_add_1225_17 (.CI(n29411), .I0(n7855[14]), .I1(GND_net), 
            .CO(n29412));
    SB_LUT4 mult_10_add_1225_16_lut (.I0(n24250), .I1(n7855[13]), .I2(n1096), 
            .I3(n29410), .O(n3048[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i35624_3_lut (.I0(n42470), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n42471));   // verilog/motorControl.v(39[10:34])
    defparam i35624_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34545_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n44533), 
            .I2(IntegralLimit[21]), .I3(n42045), .O(n41392));
    defparam i34545_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i35514_4_lut (.I0(n24_adj_3878), .I1(n8_adj_3882), .I2(n44510), 
            .I3(n41387), .O(n42361));   // verilog/motorControl.v(39[10:34])
    defparam i35514_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35054_4_lut (.I0(n13_adj_3870), .I1(n11_adj_3869), .I2(n9_adj_3873), 
            .I3(n41262), .O(n41901));
    defparam i35054_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34781_3_lut (.I0(n42471), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n41628));   // verilog/motorControl.v(39[10:34])
    defparam i34781_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3716 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3_adj_3883), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_3884));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_LUT4 i35585_3_lut (.I0(n4_adj_3884), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27), .I3(GND_net), .O(n42432));   // verilog/motorControl.v(39[38:63])
    defparam i35585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35046_4_lut (.I0(n19_adj_3875), .I1(n17_adj_3874), .I2(n15_adj_3871), 
            .I3(n41901), .O(n41893));
    defparam i35046_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35586_3_lut (.I0(n42432), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29), .I3(GND_net), .O(n42433));   // verilog/motorControl.v(39[38:63])
    defparam i35586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33), .I3(GND_net), 
            .O(n12_adj_3885));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i35816_4_lut (.I0(n25_adj_3863), .I1(n23_adj_3862), .I2(n21_adj_3876), 
            .I3(n41893), .O(n42663));
    defparam i35816_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34451_2_lut (.I0(n33), .I1(n15), .I2(GND_net), .I3(GND_net), 
            .O(n41298));
    defparam i34451_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i35356_4_lut (.I0(n31_adj_3859), .I1(n29_adj_3858), .I2(n27_adj_3872), 
            .I3(n42663), .O(n42203));
    defparam i35356_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_3841), .I3(GND_net), 
            .O(n10_adj_3886));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i35918_4_lut (.I0(n37_adj_3861), .I1(n35_adj_3867), .I2(n33_adj_3868), 
            .I3(n42203), .O(n42765));
    defparam i35918_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_3885), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35), .I3(GND_net), 
            .O(n30_adj_3887));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_CARRY mult_10_add_1225_16 (.CI(n29410), .I0(n7855[13]), .I1(n1096), 
            .CO(n29411));
    SB_LUT4 mult_10_add_1225_15_lut (.I0(n24250), .I1(n7855[12]), .I2(n1023), 
            .I3(n29409), .O(n3048[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3781_5_lut (.I0(GND_net), .I1(n8077[2]), .I2(n329), .I3(n29576), 
            .O(n8064[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3781_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34455_4_lut (.I0(n33), .I1(n31), .I2(n29), .I3(n41308), 
            .O(n41302));
    defparam i34455_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY mult_10_add_1225_15 (.CI(n29409), .I0(n7855[12]), .I1(n1023), 
            .CO(n29410));
    SB_LUT4 mult_10_add_1225_14_lut (.I0(n24250), .I1(n7855[11]), .I2(n950), 
            .I3(n29408), .O(n3048[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i35558_3_lut (.I0(n6_adj_3888), .I1(duty[10]), .I2(n21_adj_3876), 
            .I3(GND_net), .O(n42405));   // verilog/motorControl.v(44[10:25])
    defparam i35558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35559_3_lut (.I0(n42405), .I1(duty[11]), .I2(n23_adj_3862), 
            .I3(GND_net), .O(n42406));   // verilog/motorControl.v(44[10:25])
    defparam i35559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35862_4_lut (.I0(n30_adj_3887), .I1(n10_adj_3886), .I2(n35), 
            .I3(n41298), .O(n42709));   // verilog/motorControl.v(39[38:63])
    defparam i35862_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34793_3_lut (.I0(n42433), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31), .I3(GND_net), .O(n41640));   // verilog/motorControl.v(39[38:63])
    defparam i34793_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mult_10_add_1225_14 (.CI(n29408), .I0(n7855[11]), .I1(n950), 
            .CO(n29409));
    SB_LUT4 mult_10_add_1225_13_lut (.I0(n24250), .I1(n7855[10]), .I2(n877), 
            .I3(n29407), .O(n3048[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_13 (.CI(n29407), .I0(n7855[10]), .I1(n877), 
            .CO(n29408));
    SB_LUT4 i35996_4_lut (.I0(n41640), .I1(n42709), .I2(n35), .I3(n41302), 
            .O(n42843));   // verilog/motorControl.v(39[38:63])
    defparam i35996_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35997_3_lut (.I0(n42843), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37), .I3(GND_net), .O(n42844));   // verilog/motorControl.v(39[38:63])
    defparam i35997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(n16_adj_3889), .I1(duty[22]), .I2(n45_adj_3856), 
            .I3(GND_net), .O(n24_adj_3890));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35972_3_lut (.I0(n42844), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39_adj_3891), .I3(GND_net), .O(n42819));   // verilog/motorControl.v(39[38:63])
    defparam i35972_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34277_4_lut (.I0(n43_adj_3857), .I1(n25_adj_3863), .I2(n23_adj_3862), 
            .I3(n41232), .O(n41124));
    defparam i34277_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_3850), .I3(GND_net), 
            .O(n6_adj_3892));   // verilog/motorControl.v(39[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i35589_3_lut (.I0(n6_adj_3892), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_3843), .I3(GND_net), .O(n42436));   // verilog/motorControl.v(39[38:63])
    defparam i35589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35518_4_lut (.I0(n24_adj_3890), .I1(n8_adj_3893), .I2(n45_adj_3856), 
            .I3(n41120), .O(n42365));   // verilog/motorControl.v(44[10:25])
    defparam i35518_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34801_3_lut (.I0(n42406), .I1(duty[12]), .I2(n25_adj_3863), 
            .I3(GND_net), .O(n41648));   // verilog/motorControl.v(44[10:25])
    defparam i34801_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i4_4_lut (.I0(duty[0]), .I1(duty[1]), .I2(PWMLimit[1]), 
            .I3(PWMLimit[0]), .O(n4_adj_3894));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i35590_3_lut (.I0(n42436), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_3854), .I3(GND_net), .O(n42437));   // verilog/motorControl.v(39[38:63])
    defparam i35590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_add_1225_12_lut (.I0(n24250), .I1(n7855[9]), .I2(n804), 
            .I3(n29406), .O(n3048[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_12 (.CI(n29406), .I0(n7855[9]), .I1(n804), 
            .CO(n29407));
    SB_LUT4 i35554_3_lut (.I0(n4_adj_3894), .I1(duty[13]), .I2(n27_adj_3872), 
            .I3(GND_net), .O(n42401));   // verilog/motorControl.v(44[10:25])
    defparam i35554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34431_4_lut (.I0(n43), .I1(n25_adj_3853), .I2(n23_adj_3854), 
            .I3(n41333), .O(n41278));
    defparam i34431_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 mult_10_add_1225_11_lut (.I0(n24250), .I1(n7855[8]), .I2(n731), 
            .I3(n29405), .O(n3048[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_11 (.CI(n29405), .I0(n7855[8]), .I1(n731), 
            .CO(n29406));
    SB_CARRY add_3781_5 (.CI(n29576), .I0(n8077[2]), .I1(n329), .CO(n29577));
    SB_LUT4 mult_10_add_1225_10_lut (.I0(n24250), .I1(n7855[7]), .I2(n658), 
            .I3(n29404), .O(n3048[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i35555_3_lut (.I0(n42401), .I1(duty[14]), .I2(n29_adj_3858), 
            .I3(GND_net), .O(n42402));   // verilog/motorControl.v(44[10:25])
    defparam i35555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34303_4_lut (.I0(n33_adj_3868), .I1(n31_adj_3859), .I2(n29_adj_3858), 
            .I3(n41184), .O(n41150));
    defparam i34303_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35516_4_lut (.I0(n24_adj_3847), .I1(n8_adj_3846), .I2(n45), 
            .I3(n41266), .O(n42363));   // verilog/motorControl.v(39[38:63])
    defparam i35516_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 add_3781_4_lut (.I0(GND_net), .I1(n8077[1]), .I2(n256), .I3(n29575), 
            .O(n8064[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3781_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3781_4 (.CI(n29575), .I0(n8077[1]), .I1(n256), .CO(n29576));
    SB_LUT4 i34791_3_lut (.I0(n42437), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_3853), .I3(GND_net), .O(n41638));   // verilog/motorControl.v(39[38:63])
    defparam i34791_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n28027), .I0(GND_net), .I1(n1_adj_4253[5]), 
            .CO(n28028));
    SB_LUT4 i34435_4_lut (.I0(n43), .I1(n41_adj_3895), .I2(n39_adj_3891), 
            .I3(n42769), .O(n41282));
    defparam i34435_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_3781_3_lut (.I0(GND_net), .I1(n8077[0]), .I2(n183), .I3(n29574), 
            .O(n8064[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3781_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35870_4_lut (.I0(n30_adj_3881), .I1(n10_adj_3896), .I2(n35_adj_3867), 
            .I3(n41145), .O(n42717));   // verilog/motorControl.v(44[10:25])
    defparam i35870_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34803_3_lut (.I0(n42402), .I1(duty[15]), .I2(n31_adj_3859), 
            .I3(GND_net), .O(n41650));   // verilog/motorControl.v(44[10:25])
    defparam i34803_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[4]), 
            .I3(n28026), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35892_4_lut (.I0(n41638), .I1(n42363), .I2(n45), .I3(n41278), 
            .O(n42739));   // verilog/motorControl.v(39[38:63])
    defparam i35892_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i36000_4_lut (.I0(n41650), .I1(n42717), .I2(n35_adj_3867), 
            .I3(n41150), .O(n42847));   // verilog/motorControl.v(44[10:25])
    defparam i36000_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n28026), .I0(GND_net), .I1(n1_adj_4253[4]), 
            .CO(n28027));
    SB_LUT4 i34799_3_lut (.I0(n42819), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41_adj_3895), .I3(GND_net), .O(n41646));   // verilog/motorControl.v(39[38:63])
    defparam i34799_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3781_3 (.CI(n29574), .I0(n8077[0]), .I1(n183), .CO(n29575));
    SB_LUT4 add_3781_2_lut (.I0(GND_net), .I1(n41), .I2(n110_adj_3833), 
            .I3(GND_net), .O(n8064[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3781_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35894_4_lut (.I0(n41646), .I1(n42739), .I2(n45), .I3(n41282), 
            .O(n42741));   // verilog/motorControl.v(39[38:63])
    defparam i35894_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[3]), 
            .I3(n28025), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n28025), .I0(GND_net), .I1(n1_adj_4253[3]), 
            .CO(n28026));
    SB_LUT4 i36001_3_lut (.I0(n42847), .I1(duty[18]), .I2(n37_adj_3861), 
            .I3(GND_net), .O(n42848));   // verilog/motorControl.v(44[10:25])
    defparam i36001_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_3897));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_CARRY add_3781_2 (.CI(GND_net), .I0(n41), .I1(n110_adj_3833), .CO(n29574));
    SB_CARRY mult_10_add_1225_10 (.CI(n29404), .I0(n7855[7]), .I1(n658), 
            .CO(n29405));
    SB_LUT4 i35621_3_lut (.I0(n4_adj_3897), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n42468));   // verilog/motorControl.v(39[10:34])
    defparam i35621_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35622_3_lut (.I0(n42468), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n42469));   // verilog/motorControl.v(39[10:34])
    defparam i35622_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35968_3_lut (.I0(n42848), .I1(duty[19]), .I2(n39), .I3(GND_net), 
            .O(n42815));   // verilog/motorControl.v(44[10:25])
    defparam i35968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34564_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n44521), 
            .I2(IntegralLimit[16]), .I3(n42031), .O(n41411));
    defparam i34564_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i34279_4_lut (.I0(n43_adj_3857), .I1(n41_adj_3855), .I2(n39), 
            .I3(n42765), .O(n41126));
    defparam i34279_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35852_4_lut (.I0(n30), .I1(n10_adj_3866), .I2(n44544), .I3(n41406), 
            .O(n42699));   // verilog/motorControl.v(39[10:34])
    defparam i35852_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35735_4_lut (.I0(n41648), .I1(n42365), .I2(n45_adj_3856), 
            .I3(n41124), .O(n42582));   // verilog/motorControl.v(44[10:25])
    defparam i35735_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34783_3_lut (.I0(n42469), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n41630));   // verilog/motorControl.v(39[10:34])
    defparam i34783_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35986_4_lut (.I0(n41630), .I1(n42699), .I2(n44544), .I3(n41411), 
            .O(n42833));   // verilog/motorControl.v(39[10:34])
    defparam i35986_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35987_3_lut (.I0(n42833), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n42834));   // verilog/motorControl.v(39[10:34])
    defparam i35987_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35979_3_lut (.I0(n42834), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n42826));   // verilog/motorControl.v(39[10:34])
    defparam i35979_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34547_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n44512), 
            .I2(IntegralLimit[21]), .I3(n42837), .O(n41394));
    defparam i34547_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_396_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n44510));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_396_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35888_4_lut (.I0(n41628), .I1(n42361), .I2(n44510), .I3(n41392), 
            .O(n42735));   // verilog/motorControl.v(39[10:34])
    defparam i35888_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34789_3_lut (.I0(n42826), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n41636));   // verilog/motorControl.v(39[10:34])
    defparam i34789_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34809_3_lut (.I0(n42815), .I1(duty[20]), .I2(n41_adj_3855), 
            .I3(GND_net), .O(n41656));   // verilog/motorControl.v(44[10:25])
    defparam i34809_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35895_3_lut (.I0(n42741), .I1(\PID_CONTROLLER.integral_23__N_3716 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3715 ));   // verilog/motorControl.v(39[38:63])
    defparam i35895_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35896_4_lut (.I0(n41656), .I1(n42582), .I2(n45_adj_3856), 
            .I3(n41126), .O(n42743));   // verilog/motorControl.v(44[10:25])
    defparam i35896_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35890_4_lut (.I0(n41636), .I1(n42735), .I2(n44510), .I3(n41394), 
            .O(n42737));   // verilog/motorControl.v(39[10:34])
    defparam i35890_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_967_4_lut  (.I0(n42737), .I1(\PID_CONTROLLER.integral_23__N_3715 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3713 ));   // verilog/motorControl.v(39[10:63])
    defparam \PID_CONTROLLER.integral_23__I_967_4_lut .LUT_INIT = 16'h80c8;
    SB_LUT4 i35897_3_lut (.I0(n42743), .I1(PWMLimit[23]), .I2(duty[23]), 
            .I3(GND_net), .O(duty_23__N_3764));   // verilog/motorControl.v(44[10:25])
    defparam i35897_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_29_i1_3_lut (.I0(duty_23__N_3740[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[0]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_add_1225_9_lut (.I0(n24250), .I1(n7855[6]), .I2(n585), 
            .I3(n29403), .O(n3048[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3780_13_lut (.I0(GND_net), .I1(n8064[10]), .I2(n910), 
            .I3(n29573), .O(n8050[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3780_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_9 (.CI(n29403), .I0(n7855[6]), .I1(n585), 
            .CO(n29404));
    SB_LUT4 add_3780_12_lut (.I0(GND_net), .I1(n8064[9]), .I2(n837), .I3(n29572), 
            .O(n8050[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3780_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3780_12 (.CI(n29572), .I0(n8064[9]), .I1(n837), .CO(n29573));
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[2]), 
            .I3(n28024), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n28024), .I0(GND_net), .I1(n1_adj_4253[2]), 
            .CO(n28025));
    SB_LUT4 mult_10_add_1225_8_lut (.I0(n24250), .I1(n7855[5]), .I2(n512), 
            .I3(n29402), .O(n3048[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'h8228;
    SB_CARRY mult_10_add_1225_8 (.CI(n29402), .I0(n7855[5]), .I1(n512), 
            .CO(n29403));
    SB_LUT4 add_3780_11_lut (.I0(GND_net), .I1(n8064[8]), .I2(n764), .I3(n29571), 
            .O(n8050[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3780_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4253[1]), 
            .I3(n28023), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n28023), .I0(GND_net), .I1(n1_adj_4253[1]), 
            .CO(n28024));
    SB_CARRY add_3780_11 (.CI(n29571), .I0(n8064[8]), .I1(n764), .CO(n29572));
    SB_LUT4 add_3780_10_lut (.I0(GND_net), .I1(n8064[7]), .I2(n691), .I3(n29570), 
            .O(n8050[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3780_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_7_lut (.I0(n24250), .I1(n7855[4]), .I2(n439), 
            .I3(n29401), .O(n3048[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3780_10 (.CI(n29570), .I0(n8064[7]), .I1(n691), .CO(n29571));
    SB_LUT4 add_3780_9_lut (.I0(GND_net), .I1(n8064[6]), .I2(n618), .I3(n29569), 
            .O(n8050[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3780_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3780_9 (.CI(n29569), .I0(n8064[6]), .I1(n618), .CO(n29570));
    SB_LUT4 add_3780_8_lut (.I0(GND_net), .I1(n8064[5]), .I2(n545), .I3(n29568), 
            .O(n8050[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3780_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3780_8 (.CI(n29568), .I0(n8064[5]), .I1(n545), .CO(n29569));
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[5]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_20_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [18]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(n28629), .O(n1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_20_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(n25), .I1(GND_net), .I2(n1_adj_4253[0]), 
            .I3(VCC_net), .O(n40615)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3780_7_lut (.I0(GND_net), .I1(n8064[4]), .I2(n472), .I3(n29567), 
            .O(n8050[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3780_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_7 (.CI(n29401), .I0(n7855[4]), .I1(n439), 
            .CO(n29402));
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_21  (.CI(n28630), .I0(\PID_CONTROLLER.err [19]), 
            .I1(\PID_CONTROLLER.integral [19]), .CO(n28631));
    SB_LUT4 mult_10_add_1225_6_lut (.I0(n24250), .I1(n7855[3]), .I2(n366), 
            .I3(n29400), .O(n3048[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[6]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_21_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.integral [19]), .I3(n28630), .O(n1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_21_lut .LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_6 (.CI(n29400), .I0(n7855[3]), .I1(n366), 
            .CO(n29401));
    SB_LUT4 mult_10_add_1225_5_lut (.I0(n24250), .I1(n7855[2]), .I2(n293), 
            .I3(n29399), .O(n3048[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3780_7 (.CI(n29567), .I0(n8064[4]), .I1(n472), .CO(n29568));
    SB_CARRY mult_10_add_1225_5 (.CI(n29399), .I0(n7855[2]), .I1(n293), 
            .CO(n29400));
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4253[0]), 
            .CO(n28023));
    SB_LUT4 mult_10_add_1225_4_lut (.I0(n24250), .I1(n7855[1]), .I2(n220), 
            .I3(n29398), .O(n3048[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[7]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY mult_10_add_1225_4 (.CI(n29398), .I0(n7855[1]), .I1(n220), 
            .CO(n29399));
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[8]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i19532_1_lut (.I0(n256_adj_3900), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24250));   // verilog/motorControl.v(46[19:35])
    defparam i19532_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_add_1225_3_lut (.I0(n24250), .I1(n7855[0]), .I2(n147), 
            .I3(n29397), .O(n3048[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_3780_6_lut (.I0(GND_net), .I1(n8064[3]), .I2(n399), .I3(n29566), 
            .O(n8050[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3780_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3780_6 (.CI(n29566), .I0(n8064[3]), .I1(n399), .CO(n29567));
    SB_LUT4 add_3780_5_lut (.I0(GND_net), .I1(n8064[2]), .I2(n326), .I3(n29565), 
            .O(n8050[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3780_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_3 (.CI(n29397), .I0(n7855[0]), .I1(n147), 
            .CO(n29398));
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4254[23]), 
            .I3(n28022), .O(\PID_CONTROLLER.integral_23__N_3716 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_2_lut (.I0(n24250), .I1(n5), .I2(n74), .I3(GND_net), 
            .O(n3048[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_3780_5 (.CI(n29565), .I0(n8064[2]), .I1(n326), .CO(n29566));
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5), .I1(n74), .CO(n29397));
    SB_LUT4 add_3770_23_lut (.I0(GND_net), .I1(n7879[20]), .I2(GND_net), 
            .I3(n29396), .O(n7855[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3770_22_lut (.I0(GND_net), .I1(n7879[19]), .I2(GND_net), 
            .I3(n29395), .O(n7855[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1_adj_4254[22]), .I3(n28021), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n28021), .I0(GND_net), .I1(n1_adj_4254[22]), 
            .CO(n28022));
    SB_LUT4 add_3780_4_lut (.I0(GND_net), .I1(n8064[1]), .I2(n253), .I3(n29564), 
            .O(n8050[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3780_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3770_22 (.CI(n29395), .I0(n7879[19]), .I1(GND_net), .CO(n29396));
    SB_CARRY add_3780_4 (.CI(n29564), .I0(n8064[1]), .I1(n253), .CO(n29565));
    SB_LUT4 add_3770_21_lut (.I0(GND_net), .I1(n7879[18]), .I2(GND_net), 
            .I3(n29394), .O(n7855[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3770_21 (.CI(n29394), .I0(n7879[18]), .I1(GND_net), .CO(n29395));
    SB_LUT4 add_3770_20_lut (.I0(GND_net), .I1(n7879[17]), .I2(GND_net), 
            .I3(n29393), .O(n7855[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3780_3_lut (.I0(GND_net), .I1(n8064[0]), .I2(n180), .I3(n29563), 
            .O(n8050[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3780_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1_adj_4254[21]), .I3(n28020), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3770_20 (.CI(n29393), .I0(n7879[17]), .I1(GND_net), .CO(n29394));
    SB_CARRY add_3780_3 (.CI(n29563), .I0(n8064[0]), .I1(n180), .CO(n29564));
    SB_LUT4 add_3770_19_lut (.I0(GND_net), .I1(n7879[16]), .I2(GND_net), 
            .I3(n29392), .O(n7855[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_23 (.CI(n28020), .I0(GND_net), .I1(n1_adj_4254[21]), 
            .CO(n28021));
    SB_CARRY add_3770_19 (.CI(n29392), .I0(n7879[16]), .I1(GND_net), .CO(n29393));
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1_adj_4254[20]), .I3(n28019), .O(n41_adj_3895)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_22 (.CI(n28019), .I0(GND_net), .I1(n1_adj_4254[20]), 
            .CO(n28020));
    SB_LUT4 add_3780_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n8050[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3780_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3770_18_lut (.I0(GND_net), .I1(n7879[15]), .I2(GND_net), 
            .I3(n29391), .O(n7855[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3780_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n29563));
    SB_CARRY add_3770_18 (.CI(n29391), .I0(n7879[15]), .I1(GND_net), .CO(n29392));
    SB_LUT4 add_3770_17_lut (.I0(GND_net), .I1(n7879[14]), .I2(GND_net), 
            .I3(n29390), .O(n7855[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3779_14_lut (.I0(GND_net), .I1(n8050[11]), .I2(n980), 
            .I3(n29562), .O(n8035[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3779_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3779_13_lut (.I0(GND_net), .I1(n8050[10]), .I2(n907), 
            .I3(n29561), .O(n8035[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3779_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3770_17 (.CI(n29390), .I0(n7879[14]), .I1(GND_net), .CO(n29391));
    SB_CARRY add_3779_13 (.CI(n29561), .I0(n8050[10]), .I1(n907), .CO(n29562));
    SB_LUT4 add_3770_16_lut (.I0(GND_net), .I1(n7879[13]), .I2(n1099), 
            .I3(n29389), .O(n7855[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3779_12_lut (.I0(GND_net), .I1(n8050[9]), .I2(n834), .I3(n29560), 
            .O(n8035[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3779_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3779_12 (.CI(n29560), .I0(n8050[9]), .I1(n834), .CO(n29561));
    SB_CARRY add_3770_16 (.CI(n29389), .I0(n7879[13]), .I1(n1099), .CO(n29390));
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1_adj_4254[19]), .I3(n28018), .O(n39_adj_3891)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3770_15_lut (.I0(GND_net), .I1(n7879[12]), .I2(n1026), 
            .I3(n29388), .O(n7855[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3770_15 (.CI(n29388), .I0(n7879[12]), .I1(n1026), .CO(n29389));
    SB_LUT4 add_3770_14_lut (.I0(GND_net), .I1(n7879[11]), .I2(n953), 
            .I3(n29387), .O(n7855[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3770_14 (.CI(n29387), .I0(n7879[11]), .I1(n953), .CO(n29388));
    SB_LUT4 add_3770_13_lut (.I0(GND_net), .I1(n7879[10]), .I2(n880), 
            .I3(n29386), .O(n7855[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3779_11_lut (.I0(GND_net), .I1(n8050[8]), .I2(n761), .I3(n29559), 
            .O(n8035[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3779_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3770_13 (.CI(n29386), .I0(n7879[10]), .I1(n880), .CO(n29387));
    SB_CARRY unary_minus_5_add_3_21 (.CI(n28018), .I0(GND_net), .I1(n1_adj_4254[19]), 
            .CO(n28019));
    SB_CARRY add_3779_11 (.CI(n29559), .I0(n8050[8]), .I1(n761), .CO(n29560));
    SB_LUT4 add_3770_12_lut (.I0(GND_net), .I1(n7879[9]), .I2(n807), .I3(n29385), 
            .O(n7855[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[1]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3770_12 (.CI(n29385), .I0(n7879[9]), .I1(n807), .CO(n29386));
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_22_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(n28631), .O(n1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_22_lut .LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_22  (.CI(n28631), .I0(\PID_CONTROLLER.err [20]), 
            .I1(\PID_CONTROLLER.integral [20]), .CO(n28632));
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1_adj_4254[18]), .I3(n28017), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3779_10_lut (.I0(GND_net), .I1(n8050[7]), .I2(n688), .I3(n29558), 
            .O(n8035[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3779_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3770_11_lut (.I0(GND_net), .I1(n7879[8]), .I2(n734), .I3(n29384), 
            .O(n7855[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3779_10 (.CI(n29558), .I0(n8050[7]), .I1(n688), .CO(n29559));
    SB_LUT4 add_3779_9_lut (.I0(GND_net), .I1(n8050[6]), .I2(n615), .I3(n29557), 
            .O(n8035[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3779_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3770_11 (.CI(n29384), .I0(n7879[8]), .I1(n734), .CO(n29385));
    SB_LUT4 add_3770_10_lut (.I0(GND_net), .I1(n7879[7]), .I2(n661), .I3(n29383), 
            .O(n7855[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_20 (.CI(n28017), .I0(GND_net), .I1(n1_adj_4254[18]), 
            .CO(n28018));
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1_adj_4254[17]), .I3(n28016), .O(n35)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3770_10 (.CI(n29383), .I0(n7879[7]), .I1(n661), .CO(n29384));
    SB_CARRY add_3779_9 (.CI(n29557), .I0(n8050[6]), .I1(n615), .CO(n29558));
    SB_LUT4 add_3779_8_lut (.I0(GND_net), .I1(n8050[5]), .I2(n542), .I3(n29556), 
            .O(n8035[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3779_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3770_9_lut (.I0(GND_net), .I1(n7879[6]), .I2(n588), .I3(n29382), 
            .O(n7855[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3779_8 (.CI(n29556), .I0(n8050[5]), .I1(n542), .CO(n29557));
    SB_CARRY add_3770_9 (.CI(n29382), .I0(n7879[6]), .I1(n588), .CO(n29383));
    SB_LUT4 add_3770_8_lut (.I0(GND_net), .I1(n7879[5]), .I2(n515), .I3(n29381), 
            .O(n7855[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3770_8 (.CI(n29381), .I0(n7879[5]), .I1(n515), .CO(n29382));
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_3852));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3770_7_lut (.I0(GND_net), .I1(n7879[4]), .I2(n442), .I3(n29380), 
            .O(n7855[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[9]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3770_7 (.CI(n29380), .I0(n7879[4]), .I1(n442), .CO(n29381));
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[10]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3779_7_lut (.I0(GND_net), .I1(n8050[4]), .I2(n469), .I3(n29555), 
            .O(n8035[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3779_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3770_6_lut (.I0(GND_net), .I1(n7879[3]), .I2(n369), .I3(n29379), 
            .O(n7855[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3770_6 (.CI(n29379), .I0(n7879[3]), .I1(n369), .CO(n29380));
    SB_LUT4 add_3770_5_lut (.I0(GND_net), .I1(n7879[2]), .I2(n296), .I3(n29378), 
            .O(n7855[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n28016), .I0(GND_net), .I1(n1_adj_4254[17]), 
            .CO(n28017));
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1_adj_4254[16]), .I3(n28015), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3779_7 (.CI(n29555), .I0(n8050[4]), .I1(n469), .CO(n29556));
    SB_CARRY add_3770_5 (.CI(n29378), .I0(n7879[2]), .I1(n296), .CO(n29379));
    SB_LUT4 add_3779_6_lut (.I0(GND_net), .I1(n8050[3]), .I2(n396), .I3(n29554), 
            .O(n8035[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3779_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3770_4_lut (.I0(GND_net), .I1(n7879[1]), .I2(n223), .I3(n29377), 
            .O(n7855[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3770_4 (.CI(n29377), .I0(n7879[1]), .I1(n223), .CO(n29378));
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[11]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3779_6 (.CI(n29554), .I0(n8050[3]), .I1(n396), .CO(n29555));
    SB_LUT4 add_3770_3_lut (.I0(GND_net), .I1(n7879[0]), .I2(n150), .I3(n29376), 
            .O(n7855[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[12]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n28015), .I0(GND_net), .I1(n1_adj_4254[16]), 
            .CO(n28016));
    SB_LUT4 add_3779_5_lut (.I0(GND_net), .I1(n8050[2]), .I2(n323), .I3(n29553), 
            .O(n8035[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3779_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3770_3 (.CI(n29376), .I0(n7879[0]), .I1(n150), .CO(n29377));
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[13]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_3779_5 (.CI(n29553), .I0(n8050[2]), .I1(n323), .CO(n29554));
    SB_LUT4 add_3770_2_lut (.I0(GND_net), .I1(n8_adj_3904), .I2(n77), 
            .I3(GND_net), .O(n7855[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3770_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3770_2 (.CI(GND_net), .I0(n8_adj_3904), .I1(n77), .CO(n29376));
    SB_LUT4 add_3779_4_lut (.I0(GND_net), .I1(n8050[1]), .I2(n250), .I3(n29552), 
            .O(n8035[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3779_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1_adj_4254[15]), .I3(n28014), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_17 (.CI(n28014), .I0(GND_net), .I1(n1_adj_4254[15]), 
            .CO(n28015));
    SB_CARRY add_3779_4 (.CI(n29552), .I0(n8050[1]), .I1(n250), .CO(n29553));
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3779_3_lut (.I0(GND_net), .I1(n8050[0]), .I2(n177), .I3(n29551), 
            .O(n8035[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3779_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1_adj_4254[14]), .I3(n28013), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3779_3 (.CI(n29551), .I0(n8050[0]), .I1(n177), .CO(n29552));
    SB_LUT4 add_3779_2_lut (.I0(GND_net), .I1(n35_adj_3907), .I2(n104), 
            .I3(GND_net), .O(n8035[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3779_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3779_2 (.CI(GND_net), .I0(n35_adj_3907), .I1(n104), .CO(n29551));
    SB_LUT4 add_3778_15_lut (.I0(GND_net), .I1(n8035[12]), .I2(n1050), 
            .I3(n29550), .O(n8019[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3778_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3778_14_lut (.I0(GND_net), .I1(n8035[11]), .I2(n977), 
            .I3(n29549), .O(n8019[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3778_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3778_14 (.CI(n29549), .I0(n8035[11]), .I1(n977), .CO(n29550));
    SB_LUT4 add_3778_13_lut (.I0(GND_net), .I1(n8035[10]), .I2(n904), 
            .I3(n29548), .O(n8019[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3778_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3778_13 (.CI(n29548), .I0(n8035[10]), .I1(n904), .CO(n29549));
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n28013), .I0(GND_net), .I1(n1_adj_4254[14]), 
            .CO(n28014));
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[2]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3778_12_lut (.I0(GND_net), .I1(n8035[9]), .I2(n831), .I3(n29547), 
            .O(n8019[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3778_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3778_12 (.CI(n29547), .I0(n8035[9]), .I1(n831), .CO(n29548));
    SB_LUT4 add_3778_11_lut (.I0(GND_net), .I1(n8035[8]), .I2(n758), .I3(n29546), 
            .O(n8019[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3778_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3778_11 (.CI(n29546), .I0(n8035[8]), .I1(n758), .CO(n29547));
    SB_LUT4 add_3778_10_lut (.I0(GND_net), .I1(n8035[7]), .I2(n685), .I3(n29545), 
            .O(n8019[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3778_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3778_10 (.CI(n29545), .I0(n8035[7]), .I1(n685), .CO(n29546));
    SB_LUT4 add_3778_9_lut (.I0(GND_net), .I1(n8035[6]), .I2(n612), .I3(n29544), 
            .O(n8019[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3778_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1_adj_4254[13]), .I3(n28012), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n28012), .I0(GND_net), .I1(n1_adj_4254[13]), 
            .CO(n28013));
    SB_CARRY add_3778_9 (.CI(n29544), .I0(n8035[6]), .I1(n612), .CO(n29545));
    SB_LUT4 add_3778_8_lut (.I0(GND_net), .I1(n8035[5]), .I2(n539), .I3(n29543), 
            .O(n8019[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3778_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1_adj_4254[12]), .I3(n28011), .O(n25_adj_3853)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n28011), .I0(GND_net), .I1(n1_adj_4254[12]), 
            .CO(n28012));
    SB_CARRY add_3778_8 (.CI(n29543), .I0(n8035[5]), .I1(n539), .CO(n29544));
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_3837));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1_adj_4254[11]), .I3(n28010), .O(n23_adj_3854)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3778_7_lut (.I0(GND_net), .I1(n8035[4]), .I2(n466), .I3(n29542), 
            .O(n8019[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3778_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n28010), .I0(GND_net), .I1(n1_adj_4254[11]), 
            .CO(n28011));
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1_adj_4254[10]), .I3(n28009), .O(n21_adj_3843)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_12 (.CI(n28009), .I0(GND_net), .I1(n1_adj_4254[10]), 
            .CO(n28010));
    SB_CARRY add_3778_7 (.CI(n29542), .I0(n8035[4]), .I1(n466), .CO(n29543));
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1_adj_4254[9]), .I3(n28008), .O(n19)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_11 (.CI(n28008), .I0(GND_net), .I1(n1_adj_4254[9]), 
            .CO(n28009));
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1_adj_4254[8]), .I3(n28007), .O(n17_adj_3844)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n28007), .I0(GND_net), .I1(n1_adj_4254[8]), 
            .CO(n28008));
    SB_LUT4 add_3778_6_lut (.I0(GND_net), .I1(n8035[3]), .I2(n393), .I3(n29541), 
            .O(n8019[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3778_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3778_6 (.CI(n29541), .I0(n8035[3]), .I1(n393), .CO(n29542));
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1_adj_4254[7]), .I3(n28006), .O(n15)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n28006), .I0(GND_net), .I1(n1_adj_4254[7]), 
            .CO(n28007));
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_3836));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3778_5_lut (.I0(GND_net), .I1(n8035[2]), .I2(n320), .I3(n29540), 
            .O(n8019[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3778_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[14]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1_adj_4254[6]), .I3(n28005), .O(n13_adj_3841)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3778_5 (.CI(n29540), .I0(n8035[2]), .I1(n320), .CO(n29541));
    SB_CARRY unary_minus_5_add_3_8 (.CI(n28005), .I0(GND_net), .I1(n1_adj_4254[6]), 
            .CO(n28006));
    SB_LUT4 add_3778_4_lut (.I0(GND_net), .I1(n8035[1]), .I2(n247), .I3(n29539), 
            .O(n8019[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3778_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1_adj_4254[5]), .I3(n28004), .O(n11_adj_3842)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[15]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n28004), .I0(GND_net), .I1(n1_adj_4254[5]), 
            .CO(n28005));
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3778_4 (.CI(n29539), .I0(n8035[1]), .I1(n247), .CO(n29540));
    SB_LUT4 add_3778_3_lut (.I0(GND_net), .I1(n8035[0]), .I2(n174), .I3(n29538), 
            .O(n8019[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3778_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3778_3 (.CI(n29538), .I0(n8035[0]), .I1(n174), .CO(n29539));
    SB_LUT4 add_3778_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n8019[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3778_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3778_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n29538));
    SB_LUT4 add_3777_16_lut (.I0(GND_net), .I1(n8019[13]), .I2(n1120), 
            .I3(n29537), .O(n8002[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3777_15_lut (.I0(GND_net), .I1(n8019[12]), .I2(n1047), 
            .I3(n29536), .O(n8002[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3777_15 (.CI(n29536), .I0(n8019[12]), .I1(n1047), .CO(n29537));
    SB_LUT4 add_3777_14_lut (.I0(GND_net), .I1(n8019[11]), .I2(n974), 
            .I3(n29535), .O(n8002[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3777_14 (.CI(n29535), .I0(n8019[11]), .I1(n974), .CO(n29536));
    SB_LUT4 add_3777_13_lut (.I0(GND_net), .I1(n8019[10]), .I2(n901), 
            .I3(n29534), .O(n8002[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3777_13 (.CI(n29534), .I0(n8019[10]), .I1(n901), .CO(n29535));
    SB_LUT4 add_3777_12_lut (.I0(GND_net), .I1(n8019[9]), .I2(n828), .I3(n29533), 
            .O(n8002[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3777_12 (.CI(n29533), .I0(n8019[9]), .I1(n828), .CO(n29534));
    SB_LUT4 add_3777_11_lut (.I0(GND_net), .I1(n8019[8]), .I2(n755), .I3(n29532), 
            .O(n8002[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3777_11 (.CI(n29532), .I0(n8019[8]), .I1(n755), .CO(n29533));
    SB_LUT4 add_3777_10_lut (.I0(GND_net), .I1(n8019[7]), .I2(n682), .I3(n29531), 
            .O(n8002[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3777_10 (.CI(n29531), .I0(n8019[7]), .I1(n682), .CO(n29532));
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1_adj_4254[4]), .I3(n28003), .O(n9_adj_3845)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3777_9_lut (.I0(GND_net), .I1(n8019[6]), .I2(n609), .I3(n29530), 
            .O(n8002[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3777_9 (.CI(n29530), .I0(n8019[6]), .I1(n609), .CO(n29531));
    SB_LUT4 add_3777_8_lut (.I0(GND_net), .I1(n8019[5]), .I2(n536), .I3(n29529), 
            .O(n8002[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3777_8 (.CI(n29529), .I0(n8019[5]), .I1(n536), .CO(n29530));
    SB_LUT4 add_3777_7_lut (.I0(GND_net), .I1(n8019[4]), .I2(n463), .I3(n29528), 
            .O(n8002[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3777_7 (.CI(n29528), .I0(n8019[4]), .I1(n463), .CO(n29529));
    SB_CARRY unary_minus_5_add_3_6 (.CI(n28003), .I0(GND_net), .I1(n1_adj_4254[4]), 
            .CO(n28004));
    SB_LUT4 add_3777_6_lut (.I0(GND_net), .I1(n8019[3]), .I2(n390), .I3(n29527), 
            .O(n8002[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3777_6 (.CI(n29527), .I0(n8019[3]), .I1(n390), .CO(n29528));
    SB_LUT4 add_3777_5_lut (.I0(GND_net), .I1(n8019[2]), .I2(n317), .I3(n29526), 
            .O(n8002[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3777_5 (.CI(n29526), .I0(n8019[2]), .I1(n317), .CO(n29527));
    SB_LUT4 add_3777_4_lut (.I0(GND_net), .I1(n8019[1]), .I2(n244), .I3(n29525), 
            .O(n8002[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3777_4 (.CI(n29525), .I0(n8019[1]), .I1(n244), .CO(n29526));
    SB_LUT4 add_3777_3_lut (.I0(GND_net), .I1(n8019[0]), .I2(n171), .I3(n29524), 
            .O(n8002[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3777_3 (.CI(n29524), .I0(n8019[0]), .I1(n171), .CO(n29525));
    SB_LUT4 add_3777_2_lut (.I0(GND_net), .I1(n29_adj_3919), .I2(n98), 
            .I3(GND_net), .O(n8002[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3777_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3777_2 (.CI(GND_net), .I0(n29_adj_3919), .I1(n98), .CO(n29524));
    SB_LUT4 add_3776_17_lut (.I0(GND_net), .I1(n8002[14]), .I2(GND_net), 
            .I3(n29523), .O(n7984[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3776_16_lut (.I0(GND_net), .I1(n8002[13]), .I2(n1117), 
            .I3(n29522), .O(n7984[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3776_16 (.CI(n29522), .I0(n8002[13]), .I1(n1117), .CO(n29523));
    SB_LUT4 add_3776_15_lut (.I0(GND_net), .I1(n8002[12]), .I2(n1044), 
            .I3(n29521), .O(n7984[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3776_15 (.CI(n29521), .I0(n8002[12]), .I1(n1044), .CO(n29522));
    SB_LUT4 add_3776_14_lut (.I0(GND_net), .I1(n8002[11]), .I2(n971), 
            .I3(n29520), .O(n7984[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3776_14 (.CI(n29520), .I0(n8002[11]), .I1(n971), .CO(n29521));
    SB_LUT4 add_3776_13_lut (.I0(GND_net), .I1(n8002[10]), .I2(n898), 
            .I3(n29519), .O(n7984[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1_adj_4254[3]), .I3(n28002), .O(n7_adj_3850)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_3776_13 (.CI(n29519), .I0(n8002[10]), .I1(n898), .CO(n29520));
    SB_LUT4 add_3776_12_lut (.I0(GND_net), .I1(n8002[9]), .I2(n825), .I3(n29518), 
            .O(n7984[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3776_12 (.CI(n29518), .I0(n8002[9]), .I1(n825), .CO(n29519));
    SB_LUT4 add_3776_11_lut (.I0(GND_net), .I1(n8002[8]), .I2(n752), .I3(n29517), 
            .O(n7984[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3776_11 (.CI(n29517), .I0(n8002[8]), .I1(n752), .CO(n29518));
    SB_LUT4 add_3776_10_lut (.I0(GND_net), .I1(n8002[7]), .I2(n679), .I3(n29516), 
            .O(n7984[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3776_10 (.CI(n29516), .I0(n8002[7]), .I1(n679), .CO(n29517));
    SB_CARRY unary_minus_5_add_3_5 (.CI(n28002), .I0(GND_net), .I1(n1_adj_4254[3]), 
            .CO(n28003));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1_adj_4254[2]), .I3(n28001), .O(n5_adj_3851)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_4 (.CI(n28001), .I0(GND_net), .I1(n1_adj_4254[2]), 
            .CO(n28002));
    SB_LUT4 add_3776_9_lut (.I0(GND_net), .I1(n8002[6]), .I2(n606), .I3(n29515), 
            .O(n7984[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3776_9 (.CI(n29515), .I0(n8002[6]), .I1(n606), .CO(n29516));
    SB_LUT4 add_3776_8_lut (.I0(GND_net), .I1(n8002[5]), .I2(n533), .I3(n29514), 
            .O(n7984[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3776_8 (.CI(n29514), .I0(n8002[5]), .I1(n533), .CO(n29515));
    SB_LUT4 add_3776_7_lut (.I0(GND_net), .I1(n8002[4]), .I2(n460), .I3(n29513), 
            .O(n7984[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3776_7 (.CI(n29513), .I0(n8002[4]), .I1(n460), .CO(n29514));
    SB_LUT4 add_3776_6_lut (.I0(GND_net), .I1(n8002[3]), .I2(n387), .I3(n29512), 
            .O(n7984[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3776_6 (.CI(n29512), .I0(n8002[3]), .I1(n387), .CO(n29513));
    SB_LUT4 add_3776_5_lut (.I0(GND_net), .I1(n8002[2]), .I2(n314), .I3(n29511), 
            .O(n7984[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3776_5 (.CI(n29511), .I0(n8002[2]), .I1(n314), .CO(n29512));
    SB_LUT4 add_3776_4_lut (.I0(GND_net), .I1(n8002[1]), .I2(n241), .I3(n29510), 
            .O(n7984[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3776_4 (.CI(n29510), .I0(n8002[1]), .I1(n241), .CO(n29511));
    SB_LUT4 add_3776_3_lut (.I0(GND_net), .I1(n8002[0]), .I2(n168), .I3(n29509), 
            .O(n7984[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3776_3 (.CI(n29509), .I0(n8002[0]), .I1(n168), .CO(n29510));
    SB_LUT4 add_3776_2_lut (.I0(GND_net), .I1(n26), .I2(n95), .I3(GND_net), 
            .O(n7984[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3776_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3776_2 (.CI(GND_net), .I0(n26), .I1(n95), .CO(n29509));
    SB_LUT4 add_3775_18_lut (.I0(GND_net), .I1(n7984[15]), .I2(GND_net), 
            .I3(n29508), .O(n7965[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3775_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3775_17_lut (.I0(GND_net), .I1(n7984[14]), .I2(GND_net), 
            .I3(n29507), .O(n7965[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3775_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[16]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3775_17 (.CI(n29507), .I0(n7984[14]), .I1(GND_net), .CO(n29508));
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1_adj_4254[1]), .I3(n28000), .O(n3_adj_3883)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_DFFE \PID_CONTROLLER.integral_1225__i0  (.Q(\PID_CONTROLLER.integral [0]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[0]));   // verilog/motorControl.v(40[21:33])
    SB_CARRY unary_minus_5_add_3_3 (.CI(n28000), .I0(GND_net), .I1(n1_adj_4254[1]), 
            .CO(n28001));
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4254[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3716 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4254[0]), 
            .CO(n28000));
    SB_LUT4 add_3775_16_lut (.I0(GND_net), .I1(n7984[13]), .I2(n1114), 
            .I3(n29506), .O(n7965[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3775_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3775_16 (.CI(n29506), .I0(n7984[13]), .I1(n1114), .CO(n29507));
    SB_LUT4 add_3775_15_lut (.I0(GND_net), .I1(n7984[12]), .I2(n1041), 
            .I3(n29505), .O(n7965[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3775_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3775_15 (.CI(n29505), .I0(n7984[12]), .I1(n1041), .CO(n29506));
    SB_LUT4 add_3775_14_lut (.I0(GND_net), .I1(n7984[11]), .I2(n968), 
            .I3(n29504), .O(n7965[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3775_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3775_14 (.CI(n29504), .I0(n7984[11]), .I1(n968), .CO(n29505));
    SB_LUT4 add_3775_13_lut (.I0(GND_net), .I1(n7984[10]), .I2(n895), 
            .I3(n29503), .O(n7965[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3775_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3775_13 (.CI(n29503), .I0(n7984[10]), .I1(n895), .CO(n29504));
    SB_LUT4 add_3775_12_lut (.I0(GND_net), .I1(n7984[9]), .I2(n822), .I3(n29502), 
            .O(n7965[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3775_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3775_12 (.CI(n29502), .I0(n7984[9]), .I1(n822), .CO(n29503));
    SB_LUT4 add_3775_11_lut (.I0(GND_net), .I1(n7984[8]), .I2(n749), .I3(n29501), 
            .O(n7965[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3775_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3775_11 (.CI(n29501), .I0(n7984[8]), .I1(n749), .CO(n29502));
    SB_LUT4 add_3775_10_lut (.I0(GND_net), .I1(n7984[7]), .I2(n676), .I3(n29500), 
            .O(n7965[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3775_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3775_10 (.CI(n29500), .I0(n7984[7]), .I1(n676), .CO(n29501));
    SB_LUT4 add_3775_9_lut (.I0(GND_net), .I1(n7984[6]), .I2(n603), .I3(n29499), 
            .O(n7965[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3775_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3775_9 (.CI(n29499), .I0(n7984[6]), .I1(n603), .CO(n29500));
    SB_LUT4 add_3775_8_lut (.I0(GND_net), .I1(n7984[5]), .I2(n530), .I3(n29498), 
            .O(n7965[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3775_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3775_8 (.CI(n29498), .I0(n7984[5]), .I1(n530), .CO(n29499));
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[3]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[17]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[18]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[19]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[20]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[21]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[22]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i1_4_lut (.I0(\PID_CONTROLLER.integral [0]), .I1(PWMLimit[0]), 
            .I2(n256_adj_3900), .I3(\Ki[0] ), .O(n3073[0]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i1_4_lut.LUT_INIT = 16'h3a30;
    SB_LUT4 i19229_3_lut (.I0(\Kp[0] ), .I1(n256_adj_3900), .I2(\PID_CONTROLLER.err [0]), 
            .I3(GND_net), .O(n3048[0]));   // verilog/motorControl.v(46[16] 48[10])
    defparam i19229_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_3826));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i2_3_lut (.I0(n155[1]), .I1(PWMLimit[1]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[1]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i2_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4253[23]));   // verilog/motorControl.v(47[19:28])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3775_7_lut (.I0(GND_net), .I1(n7984[4]), .I2(n457), .I3(n29497), 
            .O(n7965[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3775_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3775_7 (.CI(n29497), .I0(n7984[4]), .I1(n457), .CO(n29498));
    SB_LUT4 add_3775_6_lut (.I0(GND_net), .I1(n7984[3]), .I2(n384), .I3(n29496), 
            .O(n7965[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3775_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_3919));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3775_6 (.CI(n29496), .I0(n7984[3]), .I1(n384), .CO(n29497));
    SB_LUT4 add_3775_5_lut (.I0(GND_net), .I1(n7984[2]), .I2(n311), .I3(n29495), 
            .O(n7965[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3775_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3775_5 (.CI(n29495), .I0(n7984[2]), .I1(n311), .CO(n29496));
    SB_LUT4 add_3775_4_lut (.I0(GND_net), .I1(n7984[1]), .I2(n238), .I3(n29494), 
            .O(n7965[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3775_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3775_4 (.CI(n29494), .I0(n7984[1]), .I1(n238), .CO(n29495));
    SB_LUT4 add_3775_3_lut (.I0(GND_net), .I1(n7984[0]), .I2(n165), .I3(n29493), 
            .O(n7965[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3775_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3775_3 (.CI(n29493), .I0(n7984[0]), .I1(n165), .CO(n29494));
    SB_LUT4 add_3775_2_lut (.I0(GND_net), .I1(n23_adj_3921), .I2(n92), 
            .I3(GND_net), .O(n7965[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3775_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3775_2 (.CI(GND_net), .I0(n23_adj_3921), .I1(n92), .CO(n29493));
    SB_LUT4 add_3774_19_lut (.I0(GND_net), .I1(n7965[16]), .I2(GND_net), 
            .I3(n29492), .O(n7945[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3774_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3774_18_lut (.I0(GND_net), .I1(n7965[15]), .I2(GND_net), 
            .I3(n29491), .O(n7945[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3774_18_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3617[1]));   // verilog/motorControl.v(37[14] 56[8])
    SB_CARRY add_3774_18 (.CI(n29491), .I0(n7965[15]), .I1(GND_net), .CO(n29492));
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty[22]), .I1(n257[22]), .I2(GND_net), 
            .I3(GND_net), .O(n45_adj_3922));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[4]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_3774_17_lut (.I0(GND_net), .I1(n7965[14]), .I2(GND_net), 
            .I3(n29490), .O(n7945[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3774_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3774_17 (.CI(n29490), .I0(n7965[14]), .I1(GND_net), .CO(n29491));
    SB_LUT4 add_3774_16_lut (.I0(GND_net), .I1(n7965[13]), .I2(n1111), 
            .I3(n29489), .O(n7945[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3774_16_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3617[2]));   // verilog/motorControl.v(37[14] 56[8])
    SB_CARRY add_3774_16 (.CI(n29489), .I0(n7965[13]), .I1(n1111), .CO(n29490));
    SB_LUT4 i34223_4_lut (.I0(n21_adj_3923), .I1(n19_adj_3924), .I2(n17_adj_3925), 
            .I3(n9_adj_3926), .O(n41069));
    defparam i34223_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34205_4_lut (.I0(n27_adj_3927), .I1(n15_adj_3928), .I2(n13_adj_3929), 
            .I3(n11_adj_3930), .O(n41051));
    defparam i34205_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_3931), 
            .I3(GND_net), .O(n12_adj_3932));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3617[3]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3617[4]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3617[5]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3617[6]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3617[7]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3617[8]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3617[9]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3617[10]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3617[11]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3617[12]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3617[13]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3617[14]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3617[15]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3617[16]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3617[17]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3617[18]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3617[19]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3617[20]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3617[21]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3617[22]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3617[23]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i1  (.Q(\PID_CONTROLLER.err [1]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [1]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i2  (.Q(\PID_CONTROLLER.err [2]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [2]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i3  (.Q(\PID_CONTROLLER.err [3]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [3]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i4  (.Q(\PID_CONTROLLER.err [4]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [4]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i5  (.Q(\PID_CONTROLLER.err [5]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [5]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i6  (.Q(\PID_CONTROLLER.err [6]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [6]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i7  (.Q(\PID_CONTROLLER.err [7]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [7]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i8  (.Q(\PID_CONTROLLER.err [8]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [8]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i9  (.Q(\PID_CONTROLLER.err [9]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [9]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i10  (.Q(\PID_CONTROLLER.err [10]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [10]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i11  (.Q(\PID_CONTROLLER.err [11]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [11]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i12  (.Q(\PID_CONTROLLER.err [12]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [12]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i13  (.Q(\PID_CONTROLLER.err [13]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [13]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i14  (.Q(\PID_CONTROLLER.err [14]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [14]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i15  (.Q(\PID_CONTROLLER.err [15]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [15]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i16  (.Q(\PID_CONTROLLER.err [16]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [16]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i17  (.Q(\PID_CONTROLLER.err [17]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [17]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i18  (.Q(\PID_CONTROLLER.err [18]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [18]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i19  (.Q(\PID_CONTROLLER.err [19]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [19]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i20  (.Q(\PID_CONTROLLER.err [20]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [20]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i21  (.Q(\PID_CONTROLLER.err [21]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [21]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i22  (.Q(\PID_CONTROLLER.err [22]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [22]));   // verilog/motorControl.v(37[14] 56[8])
    SB_DFF \PID_CONTROLLER.err_i23  (.Q(\PID_CONTROLLER.err [23]), .C(clk32MHz), 
           .D(\PID_CONTROLLER.err_23__N_3641 [23]));   // verilog/motorControl.v(37[14] 56[8])
    SB_LUT4 add_3774_15_lut (.I0(GND_net), .I1(n7965[12]), .I2(n1038), 
            .I3(n29488), .O(n7945[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3774_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3774_15 (.CI(n29488), .I0(n7965[12]), .I1(n1038), .CO(n29489));
    SB_LUT4 add_3774_14_lut (.I0(GND_net), .I1(n7965[11]), .I2(n965), 
            .I3(n29487), .O(n7945[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3774_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3774_14 (.CI(n29487), .I0(n7965[11]), .I1(n965), .CO(n29488));
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_3929), 
            .I3(GND_net), .O(n10_adj_3933));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_3932), .I1(n257[17]), .I2(n35_adj_3934), 
            .I3(GND_net), .O(n30_adj_3935));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_3774_13_lut (.I0(GND_net), .I1(n7965[10]), .I2(n892), 
            .I3(n29486), .O(n7945[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3774_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3774_13 (.CI(n29486), .I0(n7965[10]), .I1(n892), .CO(n29487));
    SB_LUT4 add_3774_12_lut (.I0(GND_net), .I1(n7965[9]), .I2(n819), .I3(n29485), 
            .O(n7945[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3774_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23045_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n4_adj_3936), .I3(n8431[1]), .O(n6_adj_3937));   // verilog/motorControl.v(42[26:37])
    defparam i23045_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n8431[1]), .I3(n4_adj_3936), .O(n8424[2]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_974 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n8431[0]), .I3(n27690), .O(n8424[1]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut_adj_974.LUT_INIT = 16'h8778;
    SB_CARRY add_3774_12 (.CI(n29485), .I0(n7965[9]), .I1(n819), .CO(n29486));
    SB_LUT4 add_3774_11_lut (.I0(GND_net), .I1(n7965[8]), .I2(n746), .I3(n29484), 
            .O(n7945[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3774_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3774_11 (.CI(n29484), .I0(n7965[8]), .I1(n746), .CO(n29485));
    SB_LUT4 add_3774_10_lut (.I0(GND_net), .I1(n7965[7]), .I2(n673), .I3(n29483), 
            .O(n7945[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3774_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3774_10 (.CI(n29483), .I0(n7965[7]), .I1(n673), .CO(n29484));
    SB_LUT4 add_3774_9_lut (.I0(GND_net), .I1(n7965[6]), .I2(n600), .I3(n29482), 
            .O(n7945[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3774_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3774_9 (.CI(n29482), .I0(n7965[6]), .I1(n600), .CO(n29483));
    SB_LUT4 i23037_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n27690), .I3(n8431[0]), .O(n4_adj_3936));   // verilog/motorControl.v(42[26:37])
    defparam i23037_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 add_3774_8_lut (.I0(GND_net), .I1(n7965[5]), .I2(n527), .I3(n29481), 
            .O(n7945[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3774_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3774_8 (.CI(n29481), .I0(n7965[5]), .I1(n527), .CO(n29482));
    SB_LUT4 add_3774_7_lut (.I0(GND_net), .I1(n7965[4]), .I2(n454), .I3(n29480), 
            .O(n7945[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3774_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3774_7 (.CI(n29480), .I0(n7965[4]), .I1(n454), .CO(n29481));
    SB_LUT4 add_3774_6_lut (.I0(GND_net), .I1(n7965[3]), .I2(n381), .I3(n29479), 
            .O(n7945[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3774_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i23024_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(\Ki[1] ), .O(n8424[0]));   // verilog/motorControl.v(42[26:37])
    defparam i23024_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i23026_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(\PID_CONTROLLER.integral [18]), .I3(\Ki[1] ), .O(n27690));   // verilog/motorControl.v(42[26:37])
    defparam i23026_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_3774_6 (.CI(n29479), .I0(n7965[3]), .I1(n381), .CO(n29480));
    SB_LUT4 add_3774_5_lut (.I0(GND_net), .I1(n7965[2]), .I2(n308), .I3(n29478), 
            .O(n7945[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3774_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3774_5 (.CI(n29478), .I0(n7965[2]), .I1(n308), .CO(n29479));
    SB_LUT4 add_3774_4_lut (.I0(GND_net), .I1(n7965[1]), .I2(n235), .I3(n29477), 
            .O(n7945[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3774_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3774_4 (.CI(n29477), .I0(n7965[1]), .I1(n235), .CO(n29478));
    SB_LUT4 add_3774_3_lut (.I0(GND_net), .I1(n7965[0]), .I2(n162), .I3(n29476), 
            .O(n7945[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3774_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3774_3 (.CI(n29476), .I0(n7965[0]), .I1(n162), .CO(n29477));
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23107_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n27767), .I3(n8442[0]), .O(n4_adj_3938));   // verilog/motorControl.v(42[26:37])
    defparam i23107_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_975 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n8442[0]), .I3(n27767), .O(n8437[1]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut_adj_975.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_976 (.I0(n62), .I1(n131), .I2(n8437[0]), 
            .I3(n204), .O(n8431[1]));   // verilog/motorControl.v(42[26:37])
    defparam i2_3_lut_4_lut_adj_976.LUT_INIT = 16'h8778;
    SB_LUT4 i23076_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n8437[0]), 
            .O(n4_adj_3939));   // verilog/motorControl.v(42[26:37])
    defparam i23076_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i23096_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(\Ki[1] ), .O(n27767));   // verilog/motorControl.v(42[26:37])
    defparam i23096_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23094_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(\PID_CONTROLLER.integral [20]), .I3(\Ki[1] ), .O(n8437[0]));   // verilog/motorControl.v(42[26:37])
    defparam i23094_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_3774_2_lut (.I0(GND_net), .I1(n20_adj_3940), .I2(n89), 
            .I3(GND_net), .O(n7945[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3774_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34952_4_lut (.I0(n13_adj_3929), .I1(n11_adj_3930), .I2(n9_adj_3926), 
            .I3(n41111), .O(n41799));
    defparam i34952_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i34944_4_lut (.I0(n19_adj_3924), .I1(n17_adj_3925), .I2(n15_adj_3928), 
            .I3(n41799), .O(n41791));
    defparam i34944_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35800_4_lut (.I0(n25_adj_3941), .I1(n23_adj_3942), .I2(n21_adj_3923), 
            .I3(n41791), .O(n42647));
    defparam i35800_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35326_4_lut (.I0(n31_adj_3943), .I1(n29_adj_3944), .I2(n27_adj_3927), 
            .I3(n42647), .O(n42173));
    defparam i35326_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35902_4_lut (.I0(n37_adj_3945), .I1(n35_adj_3934), .I2(n33_adj_3931), 
            .I3(n42173), .O(n42749));
    defparam i35902_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_3946), 
            .I3(GND_net), .O(n16_adj_3947));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35534_3_lut (.I0(n6_adj_3948), .I1(n257[10]), .I2(n21_adj_3923), 
            .I3(GND_net), .O(n42381));   // verilog/motorControl.v(46[19:35])
    defparam i35534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35535_3_lut (.I0(n42381), .I1(n257[11]), .I2(n23_adj_3942), 
            .I3(GND_net), .O(n42382));   // verilog/motorControl.v(46[19:35])
    defparam i35535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_3925), 
            .I3(GND_net), .O(n8_adj_3949));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_3947), .I1(n257[22]), .I2(n45_adj_3922), 
            .I3(GND_net), .O(n24_adj_3950));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34119_4_lut (.I0(n43_adj_3946), .I1(n25_adj_3941), .I2(n23_adj_3942), 
            .I3(n41069), .O(n40965));
    defparam i34119_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35520_4_lut (.I0(n24_adj_3950), .I1(n8_adj_3949), .I2(n45_adj_3922), 
            .I3(n40955), .O(n42367));   // verilog/motorControl.v(46[19:35])
    defparam i35520_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34811_3_lut (.I0(n42382), .I1(n257[12]), .I2(n25_adj_3941), 
            .I3(GND_net), .O(n41658));   // verilog/motorControl.v(46[19:35])
    defparam i34811_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_3_lut (.I0(n40615), .I1(n257[1]), .I2(duty[1]), 
            .I3(GND_net), .O(n4_adj_3951));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i4_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35532_3_lut (.I0(n4_adj_3951), .I1(n257[13]), .I2(n27_adj_3927), 
            .I3(GND_net), .O(n42379));   // verilog/motorControl.v(46[19:35])
    defparam i35532_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35533_3_lut (.I0(n42379), .I1(n257[14]), .I2(n29_adj_3944), 
            .I3(GND_net), .O(n42380));   // verilog/motorControl.v(46[19:35])
    defparam i35533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34178_4_lut (.I0(n33_adj_3931), .I1(n31_adj_3943), .I2(n29_adj_3944), 
            .I3(n41051), .O(n41024));
    defparam i34178_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35536_4_lut (.I0(n30_adj_3935), .I1(n10_adj_3933), .I2(n35_adj_3934), 
            .I3(n41016), .O(n42383));   // verilog/motorControl.v(46[19:35])
    defparam i35536_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i34813_3_lut (.I0(n42380), .I1(n257[15]), .I2(n31_adj_3943), 
            .I3(GND_net), .O(n41660));   // verilog/motorControl.v(46[19:35])
    defparam i34813_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35963_4_lut (.I0(n41660), .I1(n42383), .I2(n35_adj_3934), 
            .I3(n41024), .O(n42810));   // verilog/motorControl.v(46[19:35])
    defparam i35963_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35964_3_lut (.I0(n42810), .I1(n257[18]), .I2(n37_adj_3945), 
            .I3(GND_net), .O(n42811));   // verilog/motorControl.v(46[19:35])
    defparam i35964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35901_3_lut (.I0(n42811), .I1(n257[19]), .I2(n39_adj_3952), 
            .I3(GND_net), .O(n42748));   // verilog/motorControl.v(46[19:35])
    defparam i35901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34123_4_lut (.I0(n43_adj_3946), .I1(n41_adj_3953), .I2(n39_adj_3952), 
            .I3(n42749), .O(n40969));
    defparam i34123_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35737_4_lut (.I0(n41658), .I1(n42367), .I2(n45_adj_3922), 
            .I3(n40965), .O(n42584));   // verilog/motorControl.v(46[19:35])
    defparam i35737_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i34819_3_lut (.I0(n42748), .I1(n257[20]), .I2(n41_adj_3953), 
            .I3(GND_net), .O(n41666));   // verilog/motorControl.v(46[19:35])
    defparam i34819_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35898_4_lut (.I0(n41666), .I1(n42584), .I2(n45_adj_3922), 
            .I3(n40969), .O(n42745));   // verilog/motorControl.v(46[19:35])
    defparam i35898_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35899_3_lut (.I0(n42745), .I1(duty[23]), .I2(n47), .I3(GND_net), 
            .O(n256_adj_3900));   // verilog/motorControl.v(46[19:35])
    defparam i35899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_3774_2 (.CI(GND_net), .I0(n20_adj_3940), .I1(n89), .CO(n29476));
    SB_LUT4 add_3773_20_lut (.I0(GND_net), .I1(n7945[17]), .I2(GND_net), 
            .I3(n29475), .O(n7924[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3773_19_lut (.I0(GND_net), .I1(n7945[16]), .I2(GND_net), 
            .I3(n29474), .O(n7924[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3773_19 (.CI(n29474), .I0(n7945[16]), .I1(GND_net), .CO(n29475));
    SB_LUT4 add_3773_18_lut (.I0(GND_net), .I1(n7945[15]), .I2(GND_net), 
            .I3(n29473), .O(n7924[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3773_18 (.CI(n29473), .I0(n7945[15]), .I1(GND_net), .CO(n29474));
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_3773_17_lut (.I0(GND_net), .I1(n7945[14]), .I2(GND_net), 
            .I3(n29472), .O(n7924[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3773_17 (.CI(n29472), .I0(n7945[14]), .I1(GND_net), .CO(n29473));
    SB_LUT4 add_3773_16_lut (.I0(GND_net), .I1(n7945[13]), .I2(n1108), 
            .I3(n29471), .O(n7924[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3773_16 (.CI(n29471), .I0(n7945[13]), .I1(n1108), .CO(n29472));
    SB_LUT4 add_3773_15_lut (.I0(GND_net), .I1(n7945[12]), .I2(n1035), 
            .I3(n29470), .O(n7924[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3773_15 (.CI(n29470), .I0(n7945[12]), .I1(n1035), .CO(n29471));
    SB_DFFE \PID_CONTROLLER.integral_1225__i1  (.Q(\PID_CONTROLLER.integral [1]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[1]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i2  (.Q(\PID_CONTROLLER.integral [2]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[2]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i3  (.Q(\PID_CONTROLLER.integral [3]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[3]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i4  (.Q(\PID_CONTROLLER.integral [4]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[4]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i5  (.Q(\PID_CONTROLLER.integral [5]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[5]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i6  (.Q(\PID_CONTROLLER.integral [6]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[6]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i7  (.Q(\PID_CONTROLLER.integral [7]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[7]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i8  (.Q(\PID_CONTROLLER.integral [8]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[8]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i9  (.Q(\PID_CONTROLLER.integral [9]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[9]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i10  (.Q(\PID_CONTROLLER.integral [10]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[10]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i11  (.Q(\PID_CONTROLLER.integral [11]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[11]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i12  (.Q(\PID_CONTROLLER.integral [12]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[12]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i13  (.Q(\PID_CONTROLLER.integral [13]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[13]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i14  (.Q(\PID_CONTROLLER.integral [14]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[14]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i15  (.Q(\PID_CONTROLLER.integral [15]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[15]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i16  (.Q(\PID_CONTROLLER.integral [16]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[16]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i17  (.Q(\PID_CONTROLLER.integral [17]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[17]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i18  (.Q(\PID_CONTROLLER.integral [18]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[18]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i19  (.Q(\PID_CONTROLLER.integral [19]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[19]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i20  (.Q(\PID_CONTROLLER.integral [20]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[20]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i21  (.Q(\PID_CONTROLLER.integral [21]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[21]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i22  (.Q(\PID_CONTROLLER.integral [22]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[22]));   // verilog/motorControl.v(40[21:33])
    SB_DFFE \PID_CONTROLLER.integral_1225__i23  (.Q(\PID_CONTROLLER.integral [23]), 
            .C(clk32MHz), .E(\PID_CONTROLLER.integral_23__N_3713 ), .D(n1[23]));   // verilog/motorControl.v(40[21:33])
    SB_LUT4 add_3773_14_lut (.I0(GND_net), .I1(n7945[11]), .I2(n962), 
            .I3(n29469), .O(n7924[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3773_14 (.CI(n29469), .I0(n7945[11]), .I1(n962), .CO(n29470));
    SB_LUT4 add_3773_13_lut (.I0(GND_net), .I1(n7945[10]), .I2(n889), 
            .I3(n29468), .O(n7924[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3773_13 (.CI(n29468), .I0(n7945[10]), .I1(n889), .CO(n29469));
    SB_LUT4 add_3773_12_lut (.I0(GND_net), .I1(n7945[9]), .I2(n816), .I3(n29467), 
            .O(n7924[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_639_25_lut (.I0(GND_net), .I1(n3048[23]), .I2(n3073[23]), 
            .I3(n27975), .O(duty_23__N_3740[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3773_12 (.CI(n29467), .I0(n7945[9]), .I1(n816), .CO(n29468));
    SB_LUT4 add_3773_11_lut (.I0(GND_net), .I1(n7945[8]), .I2(n743), .I3(n29466), 
            .O(n7924[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_639_24_lut (.I0(GND_net), .I1(n3048[22]), .I2(n3073[22]), 
            .I3(n27974), .O(duty_23__N_3740[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3773_11 (.CI(n29466), .I0(n7945[8]), .I1(n743), .CO(n29467));
    SB_CARRY add_639_24 (.CI(n27974), .I0(n3048[22]), .I1(n3073[22]), 
            .CO(n27975));
    SB_LUT4 add_3773_10_lut (.I0(GND_net), .I1(n7945[7]), .I2(n670), .I3(n29465), 
            .O(n7924[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3773_10 (.CI(n29465), .I0(n7945[7]), .I1(n670), .CO(n29466));
    SB_LUT4 add_639_23_lut (.I0(GND_net), .I1(n3048[21]), .I2(n3073[21]), 
            .I3(n27973), .O(duty_23__N_3740[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3773_9_lut (.I0(GND_net), .I1(n7945[6]), .I2(n597), .I3(n29464), 
            .O(n7924[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3773_9 (.CI(n29464), .I0(n7945[6]), .I1(n597), .CO(n29465));
    SB_CARRY add_639_23 (.CI(n27973), .I0(n3048[21]), .I1(n3073[21]), 
            .CO(n27974));
    SB_LUT4 add_3773_8_lut (.I0(GND_net), .I1(n7945[5]), .I2(n524), .I3(n29463), 
            .O(n7924[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_639_22_lut (.I0(GND_net), .I1(n3048[20]), .I2(n3073[20]), 
            .I3(n27972), .O(duty_23__N_3740[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3773_8 (.CI(n29463), .I0(n7945[5]), .I1(n524), .CO(n29464));
    SB_CARRY add_639_22 (.CI(n27972), .I0(n3048[20]), .I1(n3073[20]), 
            .CO(n27973));
    SB_LUT4 add_3773_7_lut (.I0(GND_net), .I1(n7945[4]), .I2(n451), .I3(n29462), 
            .O(n7924[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_639_21_lut (.I0(GND_net), .I1(n3048[19]), .I2(n3073[19]), 
            .I3(n27971), .O(duty_23__N_3740[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3773_7 (.CI(n29462), .I0(n7945[4]), .I1(n451), .CO(n29463));
    SB_LUT4 add_3773_6_lut (.I0(GND_net), .I1(n7945[3]), .I2(n378), .I3(n29461), 
            .O(n7924[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3773_6 (.CI(n29461), .I0(n7945[3]), .I1(n378), .CO(n29462));
    SB_CARRY add_639_21 (.CI(n27971), .I0(n3048[19]), .I1(n3073[19]), 
            .CO(n27972));
    SB_LUT4 add_3773_5_lut (.I0(GND_net), .I1(n7945[2]), .I2(n305), .I3(n29460), 
            .O(n7924[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_639_20_lut (.I0(GND_net), .I1(n3048[18]), .I2(n3073[18]), 
            .I3(n27970), .O(duty_23__N_3740[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3773_5 (.CI(n29460), .I0(n7945[2]), .I1(n305), .CO(n29461));
    SB_CARRY add_639_20 (.CI(n27970), .I0(n3048[18]), .I1(n3073[18]), 
            .CO(n27971));
    SB_LUT4 add_3773_4_lut (.I0(GND_net), .I1(n7945[1]), .I2(n232), .I3(n29459), 
            .O(n7924[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3808_7_lut (.I0(GND_net), .I1(n36379), .I2(n490), .I3(n29861), 
            .O(n8416[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3808_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3808_6_lut (.I0(GND_net), .I1(n8424[3]), .I2(n417), .I3(n29860), 
            .O(n8416[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3808_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3808_6 (.CI(n29860), .I0(n8424[3]), .I1(n417), .CO(n29861));
    SB_LUT4 add_3808_5_lut (.I0(GND_net), .I1(n8424[2]), .I2(n344), .I3(n29859), 
            .O(n8416[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3808_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3808_5 (.CI(n29859), .I0(n8424[2]), .I1(n344), .CO(n29860));
    SB_LUT4 add_3808_4_lut (.I0(GND_net), .I1(n8424[1]), .I2(n271_adj_3955), 
            .I3(n29858), .O(n8416[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3808_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3808_4 (.CI(n29858), .I0(n8424[1]), .I1(n271_adj_3955), 
            .CO(n29859));
    SB_LUT4 add_3808_3_lut (.I0(GND_net), .I1(n8424[0]), .I2(n198), .I3(n29857), 
            .O(n8416[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3808_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_25_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(n28634), .O(n1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_25_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3808_3 (.CI(n29857), .I0(n8424[0]), .I1(n198), .CO(n29858));
    SB_LUT4 add_3808_2_lut (.I0(GND_net), .I1(n56), .I2(n125_adj_3956), 
            .I3(GND_net), .O(n8416[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3808_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3808_2 (.CI(GND_net), .I0(n56), .I1(n125_adj_3956), .CO(n29857));
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_24_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(n28633), .O(n1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_24_lut .LUT_INIT = 16'hC33C;
    SB_LUT4 add_3807_8_lut (.I0(GND_net), .I1(n8416[5]), .I2(n560), .I3(n29856), 
            .O(n8407[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3807_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3807_7_lut (.I0(GND_net), .I1(n8416[4]), .I2(n487), .I3(n29855), 
            .O(n8407[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3807_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3807_7 (.CI(n29855), .I0(n8416[4]), .I1(n487), .CO(n29856));
    SB_LUT4 add_3807_6_lut (.I0(GND_net), .I1(n8416[3]), .I2(n414), .I3(n29854), 
            .O(n8407[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3807_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3807_6 (.CI(n29854), .I0(n8416[3]), .I1(n414), .CO(n29855));
    SB_LUT4 add_3807_5_lut (.I0(GND_net), .I1(n8416[2]), .I2(n341), .I3(n29853), 
            .O(n8407[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3807_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_24  (.CI(n28633), .I0(\PID_CONTROLLER.err [22]), 
            .I1(\PID_CONTROLLER.integral [22]), .CO(n28634));
    SB_LUT4 \PID_CONTROLLER.integral_1225_add_4_23_lut  (.I0(GND_net), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(n28632), .O(n1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam \PID_CONTROLLER.integral_1225_add_4_23_lut .LUT_INIT = 16'hC33C;
    SB_CARRY add_3807_5 (.CI(n29853), .I0(n8416[2]), .I1(n341), .CO(n29854));
    SB_CARRY \PID_CONTROLLER.integral_1225_add_4_23  (.CI(n28632), .I0(\PID_CONTROLLER.err [21]), 
            .I1(\PID_CONTROLLER.integral [21]), .CO(n28633));
    SB_LUT4 add_3807_4_lut (.I0(GND_net), .I1(n8416[1]), .I2(n268_adj_3957), 
            .I3(n29852), .O(n8407[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3807_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3773_4 (.CI(n29459), .I0(n7945[1]), .I1(n232), .CO(n29460));
    SB_CARRY add_3807_4 (.CI(n29852), .I0(n8416[1]), .I1(n268_adj_3957), 
            .CO(n29853));
    SB_LUT4 add_3807_3_lut (.I0(GND_net), .I1(n8416[0]), .I2(n195), .I3(n29851), 
            .O(n8407[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3807_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3807_3 (.CI(n29851), .I0(n8416[0]), .I1(n195), .CO(n29852));
    SB_LUT4 add_3773_3_lut (.I0(GND_net), .I1(n7945[0]), .I2(n159), .I3(n29458), 
            .O(n7924[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3807_2_lut (.I0(GND_net), .I1(n53), .I2(n122_adj_3958), 
            .I3(GND_net), .O(n8407[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3807_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3807_2 (.CI(GND_net), .I0(n53), .I1(n122_adj_3958), .CO(n29851));
    SB_CARRY add_3773_3 (.CI(n29458), .I0(n7945[0]), .I1(n159), .CO(n29459));
    SB_LUT4 add_3806_9_lut (.I0(GND_net), .I1(n8407[6]), .I2(n630), .I3(n29850), 
            .O(n8397[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3806_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3806_8_lut (.I0(GND_net), .I1(n8407[5]), .I2(n557), .I3(n29849), 
            .O(n8397[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3806_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3806_8 (.CI(n29849), .I0(n8407[5]), .I1(n557), .CO(n29850));
    SB_LUT4 add_3806_7_lut (.I0(GND_net), .I1(n8407[4]), .I2(n484), .I3(n29848), 
            .O(n8397[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3806_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3806_7 (.CI(n29848), .I0(n8407[4]), .I1(n484), .CO(n29849));
    SB_LUT4 add_3806_6_lut (.I0(GND_net), .I1(n8407[3]), .I2(n411), .I3(n29847), 
            .O(n8397[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3806_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3806_6 (.CI(n29847), .I0(n8407[3]), .I1(n411), .CO(n29848));
    SB_LUT4 add_3806_5_lut (.I0(GND_net), .I1(n8407[2]), .I2(n338), .I3(n29846), 
            .O(n8397[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3806_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3806_5 (.CI(n29846), .I0(n8407[2]), .I1(n338), .CO(n29847));
    SB_LUT4 add_639_19_lut (.I0(GND_net), .I1(n3048[17]), .I2(n3073[17]), 
            .I3(n27969), .O(duty_23__N_3740[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3806_4_lut (.I0(GND_net), .I1(n8407[1]), .I2(n265_adj_3959), 
            .I3(n29845), .O(n8397[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3806_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3773_2_lut (.I0(GND_net), .I1(n17_adj_3960), .I2(n86), 
            .I3(GND_net), .O(n7924[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3773_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3806_4 (.CI(n29845), .I0(n8407[1]), .I1(n265_adj_3959), 
            .CO(n29846));
    SB_LUT4 add_3806_3_lut (.I0(GND_net), .I1(n8407[0]), .I2(n192), .I3(n29844), 
            .O(n8397[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3806_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3806_3 (.CI(n29844), .I0(n8407[0]), .I1(n192), .CO(n29845));
    SB_LUT4 add_3806_2_lut (.I0(GND_net), .I1(n50), .I2(n119_adj_3961), 
            .I3(GND_net), .O(n8397[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3806_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3773_2 (.CI(GND_net), .I0(n17_adj_3960), .I1(n86), .CO(n29458));
    SB_LUT4 add_3772_21_lut (.I0(GND_net), .I1(n7924[18]), .I2(GND_net), 
            .I3(n29457), .O(n7902[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3806_2 (.CI(GND_net), .I0(n50), .I1(n119_adj_3961), .CO(n29844));
    SB_LUT4 add_3805_10_lut (.I0(GND_net), .I1(n8397[7]), .I2(n700), .I3(n29843), 
            .O(n8386[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3805_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3805_9_lut (.I0(GND_net), .I1(n8397[6]), .I2(n627), .I3(n29842), 
            .O(n8386[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3805_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3805_9 (.CI(n29842), .I0(n8397[6]), .I1(n627), .CO(n29843));
    SB_LUT4 add_3805_8_lut (.I0(GND_net), .I1(n8397[5]), .I2(n554), .I3(n29841), 
            .O(n8386[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3805_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3805_8 (.CI(n29841), .I0(n8397[5]), .I1(n554), .CO(n29842));
    SB_LUT4 add_3805_7_lut (.I0(GND_net), .I1(n8397[4]), .I2(n481), .I3(n29840), 
            .O(n8386[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3805_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3805_7 (.CI(n29840), .I0(n8397[4]), .I1(n481), .CO(n29841));
    SB_LUT4 add_3805_6_lut (.I0(GND_net), .I1(n8397[3]), .I2(n408), .I3(n29839), 
            .O(n8386[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3805_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3805_6 (.CI(n29839), .I0(n8397[3]), .I1(n408), .CO(n29840));
    SB_LUT4 add_3805_5_lut (.I0(GND_net), .I1(n8397[2]), .I2(n335), .I3(n29838), 
            .O(n8386[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3805_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3805_5 (.CI(n29838), .I0(n8397[2]), .I1(n335), .CO(n29839));
    SB_CARRY add_639_19 (.CI(n27969), .I0(n3048[17]), .I1(n3073[17]), 
            .CO(n27970));
    SB_LUT4 add_3805_4_lut (.I0(GND_net), .I1(n8397[1]), .I2(n262_adj_3962), 
            .I3(n29837), .O(n8386[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3805_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3805_4 (.CI(n29837), .I0(n8397[1]), .I1(n262_adj_3962), 
            .CO(n29838));
    SB_LUT4 add_3805_3_lut (.I0(GND_net), .I1(n8397[0]), .I2(n189), .I3(n29836), 
            .O(n8386[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3805_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3805_3 (.CI(n29836), .I0(n8397[0]), .I1(n189), .CO(n29837));
    SB_LUT4 add_3805_2_lut (.I0(GND_net), .I1(n47_adj_3963), .I2(n116_adj_3964), 
            .I3(GND_net), .O(n8386[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3805_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3805_2 (.CI(GND_net), .I0(n47_adj_3963), .I1(n116_adj_3964), 
            .CO(n29836));
    SB_LUT4 add_639_18_lut (.I0(GND_net), .I1(n3048[16]), .I2(n3073[16]), 
            .I3(n27968), .O(duty_23__N_3740[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3804_11_lut (.I0(GND_net), .I1(n8386[8]), .I2(n770_adj_3965), 
            .I3(n29835), .O(n8374[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3804_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3804_10_lut (.I0(GND_net), .I1(n8386[7]), .I2(n697_adj_3966), 
            .I3(n29834), .O(n8374[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3804_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3804_10 (.CI(n29834), .I0(n8386[7]), .I1(n697_adj_3966), 
            .CO(n29835));
    SB_LUT4 add_3804_9_lut (.I0(GND_net), .I1(n8386[6]), .I2(n624_adj_3967), 
            .I3(n29833), .O(n8374[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3804_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3804_9 (.CI(n29833), .I0(n8386[6]), .I1(n624_adj_3967), 
            .CO(n29834));
    SB_LUT4 add_3804_8_lut (.I0(GND_net), .I1(n8386[5]), .I2(n551_adj_3968), 
            .I3(n29832), .O(n8374[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3804_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3804_8 (.CI(n29832), .I0(n8386[5]), .I1(n551_adj_3968), 
            .CO(n29833));
    SB_LUT4 add_3804_7_lut (.I0(GND_net), .I1(n8386[4]), .I2(n478_adj_3969), 
            .I3(n29831), .O(n8374[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3804_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3804_7 (.CI(n29831), .I0(n8386[4]), .I1(n478_adj_3969), 
            .CO(n29832));
    SB_LUT4 add_3772_20_lut (.I0(GND_net), .I1(n7924[17]), .I2(GND_net), 
            .I3(n29456), .O(n7902[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3804_6_lut (.I0(GND_net), .I1(n8386[3]), .I2(n405_adj_3970), 
            .I3(n29830), .O(n8374[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3804_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_25_lut (.I0(GND_net), .I1(motor_state[23]), 
            .I2(n1_adj_4255[23]), .I3(n28165), .O(\PID_CONTROLLER.err_23__N_3641 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3804_6 (.CI(n29830), .I0(n8386[3]), .I1(n405_adj_3970), 
            .CO(n29831));
    SB_LUT4 state_23__I_0_add_2_24_lut (.I0(GND_net), .I1(motor_state[22]), 
            .I2(n1_adj_4255[22]), .I3(n28164), .O(\PID_CONTROLLER.err_23__N_3641 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3804_5_lut (.I0(GND_net), .I1(n8386[2]), .I2(n332_adj_3973), 
            .I3(n29829), .O(n8374[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3804_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3804_5 (.CI(n29829), .I0(n8386[2]), .I1(n332_adj_3973), 
            .CO(n29830));
    SB_LUT4 add_3804_4_lut (.I0(GND_net), .I1(n8386[1]), .I2(n259_adj_3974), 
            .I3(n29828), .O(n8374[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3804_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3804_4 (.CI(n29828), .I0(n8386[1]), .I1(n259_adj_3974), 
            .CO(n29829));
    SB_LUT4 add_3804_3_lut (.I0(GND_net), .I1(n8386[0]), .I2(n186_adj_3975), 
            .I3(n29827), .O(n8374[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3804_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3772_20 (.CI(n29456), .I0(n7924[17]), .I1(GND_net), .CO(n29457));
    SB_CARRY add_3804_3 (.CI(n29827), .I0(n8386[0]), .I1(n186_adj_3975), 
            .CO(n29828));
    SB_LUT4 add_3804_2_lut (.I0(GND_net), .I1(n44_adj_3976), .I2(n113_adj_3977), 
            .I3(GND_net), .O(n8374[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3804_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3804_2 (.CI(GND_net), .I0(n44_adj_3976), .I1(n113_adj_3977), 
            .CO(n29827));
    SB_LUT4 add_3803_12_lut (.I0(GND_net), .I1(n8374[9]), .I2(n840_adj_3978), 
            .I3(n29826), .O(n8361[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3803_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_24 (.CI(n28164), .I0(motor_state[22]), 
            .I1(n1_adj_4255[22]), .CO(n28165));
    SB_LUT4 add_3803_11_lut (.I0(GND_net), .I1(n8374[8]), .I2(n767_adj_3979), 
            .I3(n29825), .O(n8361[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3803_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3803_11 (.CI(n29825), .I0(n8374[8]), .I1(n767_adj_3979), 
            .CO(n29826));
    SB_LUT4 add_3803_10_lut (.I0(GND_net), .I1(n8374[7]), .I2(n694_adj_3980), 
            .I3(n29824), .O(n8361[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3803_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_23_lut (.I0(GND_net), .I1(motor_state[21]), 
            .I2(n1_adj_4255[21]), .I3(n28163), .O(\PID_CONTROLLER.err_23__N_3641 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_23 (.CI(n28163), .I0(motor_state[21]), 
            .I1(n1_adj_4255[21]), .CO(n28164));
    SB_LUT4 state_23__I_0_add_2_22_lut (.I0(GND_net), .I1(motor_state[20]), 
            .I2(n1_adj_4255[20]), .I3(n28162), .O(\PID_CONTROLLER.err_23__N_3641 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_22 (.CI(n28162), .I0(motor_state[20]), 
            .I1(n1_adj_4255[20]), .CO(n28163));
    SB_LUT4 state_23__I_0_add_2_21_lut (.I0(GND_net), .I1(motor_state[19]), 
            .I2(n1_adj_4255[19]), .I3(n28161), .O(\PID_CONTROLLER.err_23__N_3641 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3803_10 (.CI(n29824), .I0(n8374[7]), .I1(n694_adj_3980), 
            .CO(n29825));
    SB_CARRY state_23__I_0_add_2_21 (.CI(n28161), .I0(motor_state[19]), 
            .I1(n1_adj_4255[19]), .CO(n28162));
    SB_LUT4 add_3803_9_lut (.I0(GND_net), .I1(n8374[6]), .I2(n621_adj_3984), 
            .I3(n29823), .O(n8361[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3803_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3803_9 (.CI(n29823), .I0(n8374[6]), .I1(n621_adj_3984), 
            .CO(n29824));
    SB_LUT4 add_3803_8_lut (.I0(GND_net), .I1(n8374[5]), .I2(n548_adj_3985), 
            .I3(n29822), .O(n8361[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3803_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3803_8 (.CI(n29822), .I0(n8374[5]), .I1(n548_adj_3985), 
            .CO(n29823));
    SB_LUT4 add_3803_7_lut (.I0(GND_net), .I1(n8374[4]), .I2(n475_adj_3986), 
            .I3(n29821), .O(n8361[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3803_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3803_7 (.CI(n29821), .I0(n8374[4]), .I1(n475_adj_3986), 
            .CO(n29822));
    SB_LUT4 add_3803_6_lut (.I0(GND_net), .I1(n8374[3]), .I2(n402_adj_3987), 
            .I3(n29820), .O(n8361[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3803_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3772_19_lut (.I0(GND_net), .I1(n7924[16]), .I2(GND_net), 
            .I3(n29455), .O(n7902[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_20_lut (.I0(GND_net), .I1(motor_state[18]), 
            .I2(n1_adj_4255[18]), .I3(n28160), .O(\PID_CONTROLLER.err_23__N_3641 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3772_19 (.CI(n29455), .I0(n7924[16]), .I1(GND_net), .CO(n29456));
    SB_CARRY add_3803_6 (.CI(n29820), .I0(n8374[3]), .I1(n402_adj_3987), 
            .CO(n29821));
    SB_LUT4 add_3803_5_lut (.I0(GND_net), .I1(n8374[2]), .I2(n329_adj_3989), 
            .I3(n29819), .O(n8361[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3803_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_20 (.CI(n28160), .I0(motor_state[18]), 
            .I1(n1_adj_4255[18]), .CO(n28161));
    SB_CARRY add_3803_5 (.CI(n29819), .I0(n8374[2]), .I1(n329_adj_3989), 
            .CO(n29820));
    SB_LUT4 add_3772_18_lut (.I0(GND_net), .I1(n7924[15]), .I2(GND_net), 
            .I3(n29454), .O(n7902[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3803_4_lut (.I0(GND_net), .I1(n8374[1]), .I2(n256_adj_3990), 
            .I3(n29818), .O(n8361[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3803_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3803_4 (.CI(n29818), .I0(n8374[1]), .I1(n256_adj_3990), 
            .CO(n29819));
    SB_LUT4 add_3803_3_lut (.I0(GND_net), .I1(n8374[0]), .I2(n183_adj_3991), 
            .I3(n29817), .O(n8361[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3803_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3803_3 (.CI(n29817), .I0(n8374[0]), .I1(n183_adj_3991), 
            .CO(n29818));
    SB_LUT4 add_3803_2_lut (.I0(GND_net), .I1(n41_adj_3992), .I2(n110_adj_3993), 
            .I3(GND_net), .O(n8361[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3803_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_19_lut (.I0(GND_net), .I1(motor_state[17]), 
            .I2(n1_adj_4255[17]), .I3(n28159), .O(\PID_CONTROLLER.err_23__N_3641 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_19 (.CI(n28159), .I0(motor_state[17]), 
            .I1(n1_adj_4255[17]), .CO(n28160));
    SB_LUT4 state_23__I_0_add_2_18_lut (.I0(GND_net), .I1(motor_state[16]), 
            .I2(n1_adj_4255[16]), .I3(n28158), .O(\PID_CONTROLLER.err_23__N_3641 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3803_2 (.CI(GND_net), .I0(n41_adj_3992), .I1(n110_adj_3993), 
            .CO(n29817));
    SB_CARRY state_23__I_0_add_2_18 (.CI(n28158), .I0(motor_state[16]), 
            .I1(n1_adj_4255[16]), .CO(n28159));
    SB_LUT4 add_3802_13_lut (.I0(GND_net), .I1(n8361[10]), .I2(n910_adj_3996), 
            .I3(n29816), .O(n8347[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3802_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_17_lut (.I0(GND_net), .I1(motor_state[15]), 
            .I2(n1_adj_4255[15]), .I3(n28157), .O(\PID_CONTROLLER.err_23__N_3641 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3802_12_lut (.I0(GND_net), .I1(n8361[9]), .I2(n837_adj_3998), 
            .I3(n29815), .O(n8347[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3802_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3802_12 (.CI(n29815), .I0(n8361[9]), .I1(n837_adj_3998), 
            .CO(n29816));
    SB_LUT4 add_3802_11_lut (.I0(GND_net), .I1(n8361[8]), .I2(n764_adj_3999), 
            .I3(n29814), .O(n8347[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3802_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_17 (.CI(n28157), .I0(motor_state[15]), 
            .I1(n1_adj_4255[15]), .CO(n28158));
    SB_CARRY add_3802_11 (.CI(n29814), .I0(n8361[8]), .I1(n764_adj_3999), 
            .CO(n29815));
    SB_LUT4 state_23__I_0_add_2_16_lut (.I0(GND_net), .I1(motor_state[14]), 
            .I2(n1_adj_4255[14]), .I3(n28156), .O(\PID_CONTROLLER.err_23__N_3641 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3802_10_lut (.I0(GND_net), .I1(n8361[7]), .I2(n691_adj_4001), 
            .I3(n29813), .O(n8347[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3802_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3802_10 (.CI(n29813), .I0(n8361[7]), .I1(n691_adj_4001), 
            .CO(n29814));
    SB_CARRY add_639_18 (.CI(n27968), .I0(n3048[16]), .I1(n3073[16]), 
            .CO(n27969));
    SB_LUT4 add_3802_9_lut (.I0(GND_net), .I1(n8361[6]), .I2(n618_adj_4002), 
            .I3(n29812), .O(n8347[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3802_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3802_9 (.CI(n29812), .I0(n8361[6]), .I1(n618_adj_4002), 
            .CO(n29813));
    SB_CARRY state_23__I_0_add_2_16 (.CI(n28156), .I0(motor_state[14]), 
            .I1(n1_adj_4255[14]), .CO(n28157));
    SB_LUT4 add_3802_8_lut (.I0(GND_net), .I1(n8361[5]), .I2(n545_adj_4003), 
            .I3(n29811), .O(n8347[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3802_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3802_8 (.CI(n29811), .I0(n8361[5]), .I1(n545_adj_4003), 
            .CO(n29812));
    SB_LUT4 add_3802_7_lut (.I0(GND_net), .I1(n8361[4]), .I2(n472_adj_4004), 
            .I3(n29810), .O(n8347[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3802_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3802_7 (.CI(n29810), .I0(n8361[4]), .I1(n472_adj_4004), 
            .CO(n29811));
    SB_LUT4 add_3802_6_lut (.I0(GND_net), .I1(n8361[3]), .I2(n399_adj_4005), 
            .I3(n29809), .O(n8347[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3802_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3802_6 (.CI(n29809), .I0(n8361[3]), .I1(n399_adj_4005), 
            .CO(n29810));
    SB_LUT4 add_3802_5_lut (.I0(GND_net), .I1(n8361[2]), .I2(n326_adj_4006), 
            .I3(n29808), .O(n8347[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3802_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3802_5 (.CI(n29808), .I0(n8361[2]), .I1(n326_adj_4006), 
            .CO(n29809));
    SB_LUT4 add_3802_4_lut (.I0(GND_net), .I1(n8361[1]), .I2(n253_adj_4007), 
            .I3(n29807), .O(n8347[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3802_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3802_4 (.CI(n29807), .I0(n8361[1]), .I1(n253_adj_4007), 
            .CO(n29808));
    SB_LUT4 add_3802_3_lut (.I0(GND_net), .I1(n8361[0]), .I2(n180_adj_4008), 
            .I3(n29806), .O(n8347[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3802_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3802_3 (.CI(n29806), .I0(n8361[0]), .I1(n180_adj_4008), 
            .CO(n29807));
    SB_LUT4 add_3802_2_lut (.I0(GND_net), .I1(n38_adj_4009), .I2(n107_adj_4010), 
            .I3(GND_net), .O(n8347[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3802_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3802_2 (.CI(GND_net), .I0(n38_adj_4009), .I1(n107_adj_4010), 
            .CO(n29806));
    SB_LUT4 add_3801_14_lut (.I0(GND_net), .I1(n8347[11]), .I2(n980_adj_4011), 
            .I3(n29805), .O(n8332[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3801_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3801_13_lut (.I0(GND_net), .I1(n8347[10]), .I2(n907_adj_4012), 
            .I3(n29804), .O(n8332[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3801_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3801_13 (.CI(n29804), .I0(n8347[10]), .I1(n907_adj_4012), 
            .CO(n29805));
    SB_LUT4 add_639_17_lut (.I0(GND_net), .I1(n3048[15]), .I2(n3073[15]), 
            .I3(n27967), .O(duty_23__N_3740[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3801_12_lut (.I0(GND_net), .I1(n8347[9]), .I2(n834_adj_4013), 
            .I3(n29803), .O(n8332[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3801_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3801_12 (.CI(n29803), .I0(n8347[9]), .I1(n834_adj_4013), 
            .CO(n29804));
    SB_LUT4 state_23__I_0_add_2_15_lut (.I0(GND_net), .I1(motor_state[13]), 
            .I2(n1_adj_4255[13]), .I3(n28155), .O(\PID_CONTROLLER.err_23__N_3641 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_15 (.CI(n28155), .I0(motor_state[13]), 
            .I1(n1_adj_4255[13]), .CO(n28156));
    SB_LUT4 add_3801_11_lut (.I0(GND_net), .I1(n8347[8]), .I2(n761_adj_4015), 
            .I3(n29802), .O(n8332[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3801_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3801_11 (.CI(n29802), .I0(n8347[8]), .I1(n761_adj_4015), 
            .CO(n29803));
    SB_LUT4 add_3801_10_lut (.I0(GND_net), .I1(n8347[7]), .I2(n688_adj_4016), 
            .I3(n29801), .O(n8332[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3801_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_14_lut (.I0(GND_net), .I1(motor_state[12]), 
            .I2(n1_adj_4255[12]), .I3(n28154), .O(\PID_CONTROLLER.err_23__N_3641 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3801_10 (.CI(n29801), .I0(n8347[7]), .I1(n688_adj_4016), 
            .CO(n29802));
    SB_CARRY state_23__I_0_add_2_14 (.CI(n28154), .I0(motor_state[12]), 
            .I1(n1_adj_4255[12]), .CO(n28155));
    SB_LUT4 add_3801_9_lut (.I0(GND_net), .I1(n8347[6]), .I2(n615_adj_4018), 
            .I3(n29800), .O(n8332[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3801_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3801_9 (.CI(n29800), .I0(n8347[6]), .I1(n615_adj_4018), 
            .CO(n29801));
    SB_LUT4 add_3801_8_lut (.I0(GND_net), .I1(n8347[5]), .I2(n542_adj_4019), 
            .I3(n29799), .O(n8332[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3801_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_13_lut (.I0(GND_net), .I1(motor_state[11]), 
            .I2(n1_adj_4255[11]), .I3(n28153), .O(\PID_CONTROLLER.err_23__N_3641 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3801_8 (.CI(n29799), .I0(n8347[5]), .I1(n542_adj_4019), 
            .CO(n29800));
    SB_CARRY state_23__I_0_add_2_13 (.CI(n28153), .I0(motor_state[11]), 
            .I1(n1_adj_4255[11]), .CO(n28154));
    SB_LUT4 add_3801_7_lut (.I0(GND_net), .I1(n8347[4]), .I2(n469_adj_4021), 
            .I3(n29798), .O(n8332[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3801_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_12_lut (.I0(GND_net), .I1(motor_state[10]), 
            .I2(n1_adj_4255[10]), .I3(n28152), .O(\PID_CONTROLLER.err_23__N_3641 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3801_7 (.CI(n29798), .I0(n8347[4]), .I1(n469_adj_4021), 
            .CO(n29799));
    SB_CARRY state_23__I_0_add_2_12 (.CI(n28152), .I0(motor_state[10]), 
            .I1(n1_adj_4255[10]), .CO(n28153));
    SB_LUT4 add_3801_6_lut (.I0(GND_net), .I1(n8347[3]), .I2(n396_adj_4023), 
            .I3(n29797), .O(n8332[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3801_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_11_lut (.I0(GND_net), .I1(motor_state[9]), 
            .I2(n1_adj_4255[9]), .I3(n28151), .O(\PID_CONTROLLER.err_23__N_3641 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_11 (.CI(n28151), .I0(motor_state[9]), .I1(n1_adj_4255[9]), 
            .CO(n28152));
    SB_CARRY add_3801_6 (.CI(n29797), .I0(n8347[3]), .I1(n396_adj_4023), 
            .CO(n29798));
    SB_LUT4 add_3801_5_lut (.I0(GND_net), .I1(n8347[2]), .I2(n323_adj_4025), 
            .I3(n29796), .O(n8332[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3801_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3801_5 (.CI(n29796), .I0(n8347[2]), .I1(n323_adj_4025), 
            .CO(n29797));
    SB_LUT4 add_3801_4_lut (.I0(GND_net), .I1(n8347[1]), .I2(n250_adj_4026), 
            .I3(n29795), .O(n8332[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3801_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_10_lut (.I0(GND_net), .I1(motor_state[8]), 
            .I2(n1_adj_4255[8]), .I3(n28150), .O(\PID_CONTROLLER.err_23__N_3641 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3801_4 (.CI(n29795), .I0(n8347[1]), .I1(n250_adj_4026), 
            .CO(n29796));
    SB_CARRY state_23__I_0_add_2_10 (.CI(n28150), .I0(motor_state[8]), .I1(n1_adj_4255[8]), 
            .CO(n28151));
    SB_LUT4 add_3801_3_lut (.I0(GND_net), .I1(n8347[0]), .I2(n177_adj_4028), 
            .I3(n29794), .O(n8332[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3801_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_9_lut (.I0(GND_net), .I1(motor_state[7]), 
            .I2(n1_adj_4255[7]), .I3(n28149), .O(\PID_CONTROLLER.err_23__N_3641 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3801_3 (.CI(n29794), .I0(n8347[0]), .I1(n177_adj_4028), 
            .CO(n29795));
    SB_CARRY state_23__I_0_add_2_9 (.CI(n28149), .I0(motor_state[7]), .I1(n1_adj_4255[7]), 
            .CO(n28150));
    SB_LUT4 add_3801_2_lut (.I0(GND_net), .I1(n35_adj_4030), .I2(n104_adj_4031), 
            .I3(GND_net), .O(n8332[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3801_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3801_2 (.CI(GND_net), .I0(n35_adj_4030), .I1(n104_adj_4031), 
            .CO(n29794));
    SB_LUT4 state_23__I_0_add_2_8_lut (.I0(GND_net), .I1(motor_state[6]), 
            .I2(n1_adj_4255[6]), .I3(n28148), .O(\PID_CONTROLLER.err_23__N_3641 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_8 (.CI(n28148), .I0(motor_state[6]), .I1(n1_adj_4255[6]), 
            .CO(n28149));
    SB_LUT4 state_23__I_0_add_2_7_lut (.I0(GND_net), .I1(motor_state[5]), 
            .I2(n1_adj_4255[5]), .I3(n28147), .O(\PID_CONTROLLER.err_23__N_3641 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3800_15_lut (.I0(GND_net), .I1(n8332[12]), .I2(n1050_adj_4034), 
            .I3(n29793), .O(n8316[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3800_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_7 (.CI(n28147), .I0(motor_state[5]), .I1(n1_adj_4255[5]), 
            .CO(n28148));
    SB_LUT4 add_3800_14_lut (.I0(GND_net), .I1(n8332[11]), .I2(n977_adj_4035), 
            .I3(n29792), .O(n8316[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3800_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3800_14 (.CI(n29792), .I0(n8332[11]), .I1(n977_adj_4035), 
            .CO(n29793));
    SB_LUT4 state_23__I_0_add_2_6_lut (.I0(GND_net), .I1(motor_state[4]), 
            .I2(n1_adj_4255[4]), .I3(n28146), .O(\PID_CONTROLLER.err_23__N_3641 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3800_13_lut (.I0(GND_net), .I1(n8332[10]), .I2(n904_adj_4037), 
            .I3(n29791), .O(n8316[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3800_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_6 (.CI(n28146), .I0(motor_state[4]), .I1(n1_adj_4255[4]), 
            .CO(n28147));
    SB_CARRY add_3800_13 (.CI(n29791), .I0(n8332[10]), .I1(n904_adj_4037), 
            .CO(n29792));
    SB_LUT4 add_3800_12_lut (.I0(GND_net), .I1(n8332[9]), .I2(n831_adj_4038), 
            .I3(n29790), .O(n8316[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3800_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3800_12 (.CI(n29790), .I0(n8332[9]), .I1(n831_adj_4038), 
            .CO(n29791));
    SB_LUT4 state_23__I_0_add_2_5_lut (.I0(GND_net), .I1(motor_state[3]), 
            .I2(n1_adj_4255[3]), .I3(n28145), .O(\PID_CONTROLLER.err_23__N_3641 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3800_11_lut (.I0(GND_net), .I1(n8332[8]), .I2(n758_adj_4040), 
            .I3(n29789), .O(n8316[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3800_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY state_23__I_0_add_2_5 (.CI(n28145), .I0(motor_state[3]), .I1(n1_adj_4255[3]), 
            .CO(n28146));
    SB_CARRY add_3800_11 (.CI(n29789), .I0(n8332[8]), .I1(n758_adj_4040), 
            .CO(n29790));
    SB_LUT4 add_3800_10_lut (.I0(GND_net), .I1(n8332[7]), .I2(n685_adj_4041), 
            .I3(n29788), .O(n8316[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3800_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3800_10 (.CI(n29788), .I0(n8332[7]), .I1(n685_adj_4041), 
            .CO(n29789));
    SB_LUT4 add_3800_9_lut (.I0(GND_net), .I1(n8332[6]), .I2(n612_adj_4042), 
            .I3(n29787), .O(n8316[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3800_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_4_lut (.I0(GND_net), .I1(motor_state[2]), 
            .I2(n1_adj_4255[2]), .I3(n28144), .O(\PID_CONTROLLER.err_23__N_3641 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3800_9 (.CI(n29787), .I0(n8332[6]), .I1(n612_adj_4042), 
            .CO(n29788));
    SB_CARRY state_23__I_0_add_2_4 (.CI(n28144), .I0(motor_state[2]), .I1(n1_adj_4255[2]), 
            .CO(n28145));
    SB_LUT4 state_23__I_0_add_2_3_lut (.I0(GND_net), .I1(motor_state[1]), 
            .I2(n1_adj_4255[1]), .I3(n28143), .O(\PID_CONTROLLER.err_23__N_3641 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3800_8_lut (.I0(GND_net), .I1(n8332[5]), .I2(n539_adj_4045), 
            .I3(n29786), .O(n8316[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3800_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3800_8 (.CI(n29786), .I0(n8332[5]), .I1(n539_adj_4045), 
            .CO(n29787));
    SB_CARRY state_23__I_0_add_2_3 (.CI(n28143), .I0(motor_state[1]), .I1(n1_adj_4255[1]), 
            .CO(n28144));
    SB_LUT4 add_3800_7_lut (.I0(GND_net), .I1(n8332[4]), .I2(n466_adj_4046), 
            .I3(n29785), .O(n8316[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3800_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 state_23__I_0_add_2_2_lut (.I0(GND_net), .I1(motor_state[0]), 
            .I2(n1_adj_4255[0]), .I3(VCC_net), .O(\PID_CONTROLLER.err_23__N_3641 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam state_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3800_7 (.CI(n29785), .I0(n8332[4]), .I1(n466_adj_4046), 
            .CO(n29786));
    SB_LUT4 add_3800_6_lut (.I0(GND_net), .I1(n8332[3]), .I2(n393_adj_4048), 
            .I3(n29784), .O(n8316[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3800_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3800_6 (.CI(n29784), .I0(n8332[3]), .I1(n393_adj_4048), 
            .CO(n29785));
    SB_CARRY state_23__I_0_add_2_2 (.CI(VCC_net), .I0(motor_state[0]), .I1(n1_adj_4255[0]), 
            .CO(n28143));
    SB_LUT4 add_3800_5_lut (.I0(GND_net), .I1(n8332[2]), .I2(n320_adj_4049), 
            .I3(n29783), .O(n8316[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3800_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3800_5 (.CI(n29783), .I0(n8332[2]), .I1(n320_adj_4049), 
            .CO(n29784));
    SB_LUT4 add_3800_4_lut (.I0(GND_net), .I1(n8332[1]), .I2(n247_adj_4050), 
            .I3(n29782), .O(n8316[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3800_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3800_4 (.CI(n29782), .I0(n8332[1]), .I1(n247_adj_4050), 
            .CO(n29783));
    SB_LUT4 add_3800_3_lut (.I0(GND_net), .I1(n8332[0]), .I2(n174_adj_4051), 
            .I3(n29781), .O(n8316[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3800_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3800_3 (.CI(n29781), .I0(n8332[0]), .I1(n174_adj_4051), 
            .CO(n29782));
    SB_LUT4 add_3800_2_lut (.I0(GND_net), .I1(n32_adj_4052), .I2(n101_adj_4053), 
            .I3(GND_net), .O(n8316[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3800_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3772_18 (.CI(n29454), .I0(n7924[15]), .I1(GND_net), .CO(n29455));
    SB_CARRY add_3800_2 (.CI(GND_net), .I0(n32_adj_4052), .I1(n101_adj_4053), 
            .CO(n29781));
    SB_LUT4 add_3799_16_lut (.I0(GND_net), .I1(n8316[13]), .I2(n1120_adj_4054), 
            .I3(n29780), .O(n8299[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3799_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3799_15_lut (.I0(GND_net), .I1(n8316[12]), .I2(n1047_adj_4055), 
            .I3(n29779), .O(n8299[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3799_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3799_15 (.CI(n29779), .I0(n8316[12]), .I1(n1047_adj_4055), 
            .CO(n29780));
    SB_CARRY add_639_17 (.CI(n27967), .I0(n3048[15]), .I1(n3073[15]), 
            .CO(n27968));
    SB_LUT4 add_3799_14_lut (.I0(GND_net), .I1(n8316[11]), .I2(n974_adj_4056), 
            .I3(n29778), .O(n8299[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3799_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3799_14 (.CI(n29778), .I0(n8316[11]), .I1(n974_adj_4056), 
            .CO(n29779));
    SB_LUT4 add_3799_13_lut (.I0(GND_net), .I1(n8316[10]), .I2(n901_adj_4057), 
            .I3(n29777), .O(n8299[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3799_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3799_13 (.CI(n29777), .I0(n8316[10]), .I1(n901_adj_4057), 
            .CO(n29778));
    SB_LUT4 add_3799_12_lut (.I0(GND_net), .I1(n8316[9]), .I2(n828_adj_4058), 
            .I3(n29776), .O(n8299[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3799_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3799_12 (.CI(n29776), .I0(n8316[9]), .I1(n828_adj_4058), 
            .CO(n29777));
    SB_LUT4 add_3799_11_lut (.I0(GND_net), .I1(n8316[8]), .I2(n755_adj_4059), 
            .I3(n29775), .O(n8299[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3799_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_639_16_lut (.I0(GND_net), .I1(n3048[14]), .I2(n3073[14]), 
            .I3(n27966), .O(duty_23__N_3740[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3799_11 (.CI(n29775), .I0(n8316[8]), .I1(n755_adj_4059), 
            .CO(n29776));
    SB_LUT4 add_3799_10_lut (.I0(GND_net), .I1(n8316[7]), .I2(n682_adj_4060), 
            .I3(n29774), .O(n8299[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3799_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3799_10 (.CI(n29774), .I0(n8316[7]), .I1(n682_adj_4060), 
            .CO(n29775));
    SB_LUT4 add_3799_9_lut (.I0(GND_net), .I1(n8316[6]), .I2(n609_adj_4061), 
            .I3(n29773), .O(n8299[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3799_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_639_16 (.CI(n27966), .I0(n3048[14]), .I1(n3073[14]), 
            .CO(n27967));
    SB_LUT4 add_3772_17_lut (.I0(GND_net), .I1(n7924[14]), .I2(GND_net), 
            .I3(n29453), .O(n7902[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3799_9 (.CI(n29773), .I0(n8316[6]), .I1(n609_adj_4061), 
            .CO(n29774));
    SB_LUT4 add_3799_8_lut (.I0(GND_net), .I1(n8316[5]), .I2(n536_adj_4062), 
            .I3(n29772), .O(n8299[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3799_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3799_8 (.CI(n29772), .I0(n8316[5]), .I1(n536_adj_4062), 
            .CO(n29773));
    SB_LUT4 add_3799_7_lut (.I0(GND_net), .I1(n8316[4]), .I2(n463_adj_4063), 
            .I3(n29771), .O(n8299[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3799_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3799_7 (.CI(n29771), .I0(n8316[4]), .I1(n463_adj_4063), 
            .CO(n29772));
    SB_LUT4 add_3799_6_lut (.I0(GND_net), .I1(n8316[3]), .I2(n390_adj_4064), 
            .I3(n29770), .O(n8299[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3799_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3799_6 (.CI(n29770), .I0(n8316[3]), .I1(n390_adj_4064), 
            .CO(n29771));
    SB_LUT4 add_3799_5_lut (.I0(GND_net), .I1(n8316[2]), .I2(n317_adj_4065), 
            .I3(n29769), .O(n8299[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3799_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3799_5 (.CI(n29769), .I0(n8316[2]), .I1(n317_adj_4065), 
            .CO(n29770));
    SB_LUT4 add_3799_4_lut (.I0(GND_net), .I1(n8316[1]), .I2(n244_adj_4066), 
            .I3(n29768), .O(n8299[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3799_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3799_4 (.CI(n29768), .I0(n8316[1]), .I1(n244_adj_4066), 
            .CO(n29769));
    SB_LUT4 add_3799_3_lut (.I0(GND_net), .I1(n8316[0]), .I2(n171_adj_4067), 
            .I3(n29767), .O(n8299[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3799_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_639_15_lut (.I0(GND_net), .I1(n3048[13]), .I2(n3073[13]), 
            .I3(n27965), .O(duty_23__N_3740[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3799_3 (.CI(n29767), .I0(n8316[0]), .I1(n171_adj_4067), 
            .CO(n29768));
    SB_LUT4 add_3799_2_lut (.I0(GND_net), .I1(n29_adj_4068), .I2(n98_adj_4069), 
            .I3(GND_net), .O(n8299[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3799_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_639_15 (.CI(n27965), .I0(n3048[13]), .I1(n3073[13]), 
            .CO(n27966));
    SB_CARRY add_3799_2 (.CI(GND_net), .I0(n29_adj_4068), .I1(n98_adj_4069), 
            .CO(n29767));
    SB_LUT4 add_3798_17_lut (.I0(GND_net), .I1(n8299[14]), .I2(GND_net), 
            .I3(n29766), .O(n8281[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3798_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3798_16_lut (.I0(GND_net), .I1(n8299[13]), .I2(n1117_adj_4070), 
            .I3(n29765), .O(n8281[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3798_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3798_16 (.CI(n29765), .I0(n8299[13]), .I1(n1117_adj_4070), 
            .CO(n29766));
    SB_LUT4 add_3798_15_lut (.I0(GND_net), .I1(n8299[12]), .I2(n1044_adj_4071), 
            .I3(n29764), .O(n8281[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3798_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_639_14_lut (.I0(GND_net), .I1(n3048[12]), .I2(n3073[12]), 
            .I3(n27964), .O(duty_23__N_3740[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3798_15 (.CI(n29764), .I0(n8299[12]), .I1(n1044_adj_4071), 
            .CO(n29765));
    SB_LUT4 add_3798_14_lut (.I0(GND_net), .I1(n8299[11]), .I2(n971_adj_4072), 
            .I3(n29763), .O(n8281[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3798_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3798_14 (.CI(n29763), .I0(n8299[11]), .I1(n971_adj_4072), 
            .CO(n29764));
    SB_LUT4 add_3798_13_lut (.I0(GND_net), .I1(n8299[10]), .I2(n898_adj_4073), 
            .I3(n29762), .O(n8281[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3798_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_639_14 (.CI(n27964), .I0(n3048[12]), .I1(n3073[12]), 
            .CO(n27965));
    SB_CARRY add_3798_13 (.CI(n29762), .I0(n8299[10]), .I1(n898_adj_4073), 
            .CO(n29763));
    SB_LUT4 add_3798_12_lut (.I0(GND_net), .I1(n8299[9]), .I2(n825_adj_4074), 
            .I3(n29761), .O(n8281[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3798_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3798_12 (.CI(n29761), .I0(n8299[9]), .I1(n825_adj_4074), 
            .CO(n29762));
    SB_CARRY add_3772_17 (.CI(n29453), .I0(n7924[14]), .I1(GND_net), .CO(n29454));
    SB_LUT4 add_3798_11_lut (.I0(GND_net), .I1(n8299[8]), .I2(n752_adj_4075), 
            .I3(n29760), .O(n8281[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3798_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3798_11 (.CI(n29760), .I0(n8299[8]), .I1(n752_adj_4075), 
            .CO(n29761));
    SB_LUT4 add_3798_10_lut (.I0(GND_net), .I1(n8299[7]), .I2(n679_adj_4076), 
            .I3(n29759), .O(n8281[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3798_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_639_13_lut (.I0(GND_net), .I1(n3048[11]), .I2(n3073[11]), 
            .I3(n27963), .O(duty_23__N_3740[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3798_10 (.CI(n29759), .I0(n8299[7]), .I1(n679_adj_4076), 
            .CO(n29760));
    SB_LUT4 add_3798_9_lut (.I0(GND_net), .I1(n8299[6]), .I2(n606_adj_4077), 
            .I3(n29758), .O(n8281[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3798_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3798_9 (.CI(n29758), .I0(n8299[6]), .I1(n606_adj_4077), 
            .CO(n29759));
    SB_LUT4 add_3798_8_lut (.I0(GND_net), .I1(n8299[5]), .I2(n533_adj_4078), 
            .I3(n29757), .O(n8281[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3798_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3798_8 (.CI(n29757), .I0(n8299[5]), .I1(n533_adj_4078), 
            .CO(n29758));
    SB_LUT4 add_3798_7_lut (.I0(GND_net), .I1(n8299[4]), .I2(n460_adj_4079), 
            .I3(n29756), .O(n8281[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3798_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3798_7 (.CI(n29756), .I0(n8299[4]), .I1(n460_adj_4079), 
            .CO(n29757));
    SB_LUT4 add_3798_6_lut (.I0(GND_net), .I1(n8299[3]), .I2(n387_adj_4080), 
            .I3(n29755), .O(n8281[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3798_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3798_6 (.CI(n29755), .I0(n8299[3]), .I1(n387_adj_4080), 
            .CO(n29756));
    SB_LUT4 add_3798_5_lut (.I0(GND_net), .I1(n8299[2]), .I2(n314_adj_4081), 
            .I3(n29754), .O(n8281[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3798_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3798_5 (.CI(n29754), .I0(n8299[2]), .I1(n314_adj_4081), 
            .CO(n29755));
    SB_LUT4 add_3798_4_lut (.I0(GND_net), .I1(n8299[1]), .I2(n241_adj_4082), 
            .I3(n29753), .O(n8281[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3798_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3798_4 (.CI(n29753), .I0(n8299[1]), .I1(n241_adj_4082), 
            .CO(n29754));
    SB_LUT4 add_3798_3_lut (.I0(GND_net), .I1(n8299[0]), .I2(n168_adj_4083), 
            .I3(n29752), .O(n8281[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3798_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3772_16_lut (.I0(GND_net), .I1(n7924[13]), .I2(n1105), 
            .I3(n29452), .O(n7902[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3798_3 (.CI(n29752), .I0(n8299[0]), .I1(n168_adj_4083), 
            .CO(n29753));
    SB_LUT4 add_3798_2_lut (.I0(GND_net), .I1(n26_adj_4084), .I2(n95_adj_4085), 
            .I3(GND_net), .O(n8281[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3798_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3798_2 (.CI(GND_net), .I0(n26_adj_4084), .I1(n95_adj_4085), 
            .CO(n29752));
    SB_LUT4 add_3797_18_lut (.I0(GND_net), .I1(n8281[15]), .I2(GND_net), 
            .I3(n29751), .O(n8262[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3797_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_639_13 (.CI(n27963), .I0(n3048[11]), .I1(n3073[11]), 
            .CO(n27964));
    SB_LUT4 add_3797_17_lut (.I0(GND_net), .I1(n8281[14]), .I2(GND_net), 
            .I3(n29750), .O(n8262[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3797_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3797_17 (.CI(n29750), .I0(n8281[14]), .I1(GND_net), .CO(n29751));
    SB_LUT4 add_639_12_lut (.I0(GND_net), .I1(n3048[10]), .I2(n3073[10]), 
            .I3(n27962), .O(duty_23__N_3740[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3797_16_lut (.I0(GND_net), .I1(n8281[13]), .I2(n1114_adj_4086), 
            .I3(n29749), .O(n8262[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3797_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3797_16 (.CI(n29749), .I0(n8281[13]), .I1(n1114_adj_4086), 
            .CO(n29750));
    SB_LUT4 add_3797_15_lut (.I0(GND_net), .I1(n8281[12]), .I2(n1041_adj_4087), 
            .I3(n29748), .O(n8262[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3797_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3797_15 (.CI(n29748), .I0(n8281[12]), .I1(n1041_adj_4087), 
            .CO(n29749));
    SB_LUT4 add_3797_14_lut (.I0(GND_net), .I1(n8281[11]), .I2(n968_adj_4088), 
            .I3(n29747), .O(n8262[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3797_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3797_14 (.CI(n29747), .I0(n8281[11]), .I1(n968_adj_4088), 
            .CO(n29748));
    SB_CARRY add_639_12 (.CI(n27962), .I0(n3048[10]), .I1(n3073[10]), 
            .CO(n27963));
    SB_LUT4 add_3797_13_lut (.I0(GND_net), .I1(n8281[10]), .I2(n895_adj_4089), 
            .I3(n29746), .O(n8262[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3797_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3797_13 (.CI(n29746), .I0(n8281[10]), .I1(n895_adj_4089), 
            .CO(n29747));
    SB_LUT4 add_3797_12_lut (.I0(GND_net), .I1(n8281[9]), .I2(n822_adj_4090), 
            .I3(n29745), .O(n8262[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3797_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3797_12 (.CI(n29745), .I0(n8281[9]), .I1(n822_adj_4090), 
            .CO(n29746));
    SB_LUT4 add_3797_11_lut (.I0(GND_net), .I1(n8281[8]), .I2(n749_adj_4091), 
            .I3(n29744), .O(n8262[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3797_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3797_11 (.CI(n29744), .I0(n8281[8]), .I1(n749_adj_4091), 
            .CO(n29745));
    SB_LUT4 add_3797_10_lut (.I0(GND_net), .I1(n8281[7]), .I2(n676_adj_4092), 
            .I3(n29743), .O(n8262[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3797_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3797_10 (.CI(n29743), .I0(n8281[7]), .I1(n676_adj_4092), 
            .CO(n29744));
    SB_LUT4 add_3797_9_lut (.I0(GND_net), .I1(n8281[6]), .I2(n603_adj_4093), 
            .I3(n29742), .O(n8262[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3797_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3797_9 (.CI(n29742), .I0(n8281[6]), .I1(n603_adj_4093), 
            .CO(n29743));
    SB_LUT4 add_3797_8_lut (.I0(GND_net), .I1(n8281[5]), .I2(n530_adj_4094), 
            .I3(n29741), .O(n8262[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3797_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3797_8 (.CI(n29741), .I0(n8281[5]), .I1(n530_adj_4094), 
            .CO(n29742));
    SB_LUT4 add_3797_7_lut (.I0(GND_net), .I1(n8281[4]), .I2(n457_adj_4095), 
            .I3(n29740), .O(n8262[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3797_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3797_7 (.CI(n29740), .I0(n8281[4]), .I1(n457_adj_4095), 
            .CO(n29741));
    SB_LUT4 add_3797_6_lut (.I0(GND_net), .I1(n8281[3]), .I2(n384_adj_4096), 
            .I3(n29739), .O(n8262[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3797_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3797_6 (.CI(n29739), .I0(n8281[3]), .I1(n384_adj_4096), 
            .CO(n29740));
    SB_LUT4 add_3797_5_lut (.I0(GND_net), .I1(n8281[2]), .I2(n311_adj_4097), 
            .I3(n29738), .O(n8262[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3797_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_639_11_lut (.I0(GND_net), .I1(n3048[9]), .I2(n3073[9]), 
            .I3(n27961), .O(duty_23__N_3740[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3797_5 (.CI(n29738), .I0(n8281[2]), .I1(n311_adj_4097), 
            .CO(n29739));
    SB_LUT4 add_3797_4_lut (.I0(GND_net), .I1(n8281[1]), .I2(n238_adj_4098), 
            .I3(n29737), .O(n8262[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3797_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3797_4 (.CI(n29737), .I0(n8281[1]), .I1(n238_adj_4098), 
            .CO(n29738));
    SB_LUT4 add_3797_3_lut (.I0(GND_net), .I1(n8281[0]), .I2(n165_adj_4099), 
            .I3(n29736), .O(n8262[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3797_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3772_16 (.CI(n29452), .I0(n7924[13]), .I1(n1105), .CO(n29453));
    SB_CARRY add_3797_3 (.CI(n29736), .I0(n8281[0]), .I1(n165_adj_4099), 
            .CO(n29737));
    SB_LUT4 add_3797_2_lut (.I0(GND_net), .I1(n23_adj_4100), .I2(n92_adj_4101), 
            .I3(GND_net), .O(n8262[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3797_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3797_2 (.CI(GND_net), .I0(n23_adj_4100), .I1(n92_adj_4101), 
            .CO(n29736));
    SB_LUT4 add_3796_19_lut (.I0(GND_net), .I1(n8262[16]), .I2(GND_net), 
            .I3(n29735), .O(n8242[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3796_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3796_18_lut (.I0(GND_net), .I1(n8262[15]), .I2(GND_net), 
            .I3(n29734), .O(n8242[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3796_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3796_18 (.CI(n29734), .I0(n8262[15]), .I1(GND_net), .CO(n29735));
    SB_LUT4 add_3796_17_lut (.I0(GND_net), .I1(n8262[14]), .I2(GND_net), 
            .I3(n29733), .O(n8242[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3796_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3796_17 (.CI(n29733), .I0(n8262[14]), .I1(GND_net), .CO(n29734));
    SB_LUT4 add_3796_16_lut (.I0(GND_net), .I1(n8262[13]), .I2(n1111_adj_4102), 
            .I3(n29732), .O(n8242[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3796_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_639_11 (.CI(n27961), .I0(n3048[9]), .I1(n3073[9]), .CO(n27962));
    SB_CARRY add_3796_16 (.CI(n29732), .I0(n8262[13]), .I1(n1111_adj_4102), 
            .CO(n29733));
    SB_LUT4 add_3796_15_lut (.I0(GND_net), .I1(n8262[12]), .I2(n1038_adj_4103), 
            .I3(n29731), .O(n8242[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3796_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_639_10_lut (.I0(GND_net), .I1(n3048[8]), .I2(n3073[8]), 
            .I3(n27960), .O(duty_23__N_3740[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3796_15 (.CI(n29731), .I0(n8262[12]), .I1(n1038_adj_4103), 
            .CO(n29732));
    SB_LUT4 add_3796_14_lut (.I0(GND_net), .I1(n8262[11]), .I2(n965_adj_4104), 
            .I3(n29730), .O(n8242[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3796_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3796_14 (.CI(n29730), .I0(n8262[11]), .I1(n965_adj_4104), 
            .CO(n29731));
    SB_LUT4 add_3796_13_lut (.I0(GND_net), .I1(n8262[10]), .I2(n892_adj_4105), 
            .I3(n29729), .O(n8242[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3796_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3796_13 (.CI(n29729), .I0(n8262[10]), .I1(n892_adj_4105), 
            .CO(n29730));
    SB_LUT4 add_3796_12_lut (.I0(GND_net), .I1(n8262[9]), .I2(n819_adj_4106), 
            .I3(n29728), .O(n8242[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3796_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3796_12 (.CI(n29728), .I0(n8262[9]), .I1(n819_adj_4106), 
            .CO(n29729));
    SB_LUT4 add_3772_15_lut (.I0(GND_net), .I1(n7924[12]), .I2(n1032), 
            .I3(n29451), .O(n7902[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3796_11_lut (.I0(GND_net), .I1(n8262[8]), .I2(n746_adj_4107), 
            .I3(n29727), .O(n8242[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3796_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3796_11 (.CI(n29727), .I0(n8262[8]), .I1(n746_adj_4107), 
            .CO(n29728));
    SB_LUT4 add_3796_10_lut (.I0(GND_net), .I1(n8262[7]), .I2(n673_adj_4108), 
            .I3(n29726), .O(n8242[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3796_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3796_10 (.CI(n29726), .I0(n8262[7]), .I1(n673_adj_4108), 
            .CO(n29727));
    SB_LUT4 add_3796_9_lut (.I0(GND_net), .I1(n8262[6]), .I2(n600_adj_4109), 
            .I3(n29725), .O(n8242[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3796_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3796_9 (.CI(n29725), .I0(n8262[6]), .I1(n600_adj_4109), 
            .CO(n29726));
    SB_LUT4 add_3796_8_lut (.I0(GND_net), .I1(n8262[5]), .I2(n527_adj_4110), 
            .I3(n29724), .O(n8242[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3796_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3796_8 (.CI(n29724), .I0(n8262[5]), .I1(n527_adj_4110), 
            .CO(n29725));
    SB_LUT4 add_3796_7_lut (.I0(GND_net), .I1(n8262[4]), .I2(n454_adj_4111), 
            .I3(n29723), .O(n8242[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3796_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3796_7 (.CI(n29723), .I0(n8262[4]), .I1(n454_adj_4111), 
            .CO(n29724));
    SB_LUT4 add_3796_6_lut (.I0(GND_net), .I1(n8262[3]), .I2(n381_adj_4112), 
            .I3(n29722), .O(n8242[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3796_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3796_6 (.CI(n29722), .I0(n8262[3]), .I1(n381_adj_4112), 
            .CO(n29723));
    SB_LUT4 add_3796_5_lut (.I0(GND_net), .I1(n8262[2]), .I2(n308_adj_4113), 
            .I3(n29721), .O(n8242[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3796_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3796_5 (.CI(n29721), .I0(n8262[2]), .I1(n308_adj_4113), 
            .CO(n29722));
    SB_LUT4 add_3796_4_lut (.I0(GND_net), .I1(n8262[1]), .I2(n235_adj_4114), 
            .I3(n29720), .O(n8242[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3796_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3796_4 (.CI(n29720), .I0(n8262[1]), .I1(n235_adj_4114), 
            .CO(n29721));
    SB_LUT4 add_3796_3_lut (.I0(GND_net), .I1(n8262[0]), .I2(n162_adj_4115), 
            .I3(n29719), .O(n8242[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3796_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3796_3 (.CI(n29719), .I0(n8262[0]), .I1(n162_adj_4115), 
            .CO(n29720));
    SB_LUT4 add_3796_2_lut (.I0(GND_net), .I1(n20_adj_4116), .I2(n89_adj_4117), 
            .I3(GND_net), .O(n8242[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3796_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3796_2 (.CI(GND_net), .I0(n20_adj_4116), .I1(n89_adj_4117), 
            .CO(n29719));
    SB_LUT4 add_3795_20_lut (.I0(GND_net), .I1(n8242[17]), .I2(GND_net), 
            .I3(n29718), .O(n8221[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3795_19_lut (.I0(GND_net), .I1(n8242[16]), .I2(GND_net), 
            .I3(n29717), .O(n8221[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_639_10 (.CI(n27960), .I0(n3048[8]), .I1(n3073[8]), .CO(n27961));
    SB_CARRY add_3795_19 (.CI(n29717), .I0(n8242[16]), .I1(GND_net), .CO(n29718));
    SB_LUT4 add_3795_18_lut (.I0(GND_net), .I1(n8242[15]), .I2(GND_net), 
            .I3(n29716), .O(n8221[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3795_18 (.CI(n29716), .I0(n8242[15]), .I1(GND_net), .CO(n29717));
    SB_LUT4 add_3795_17_lut (.I0(GND_net), .I1(n8242[14]), .I2(GND_net), 
            .I3(n29715), .O(n8221[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3795_17 (.CI(n29715), .I0(n8242[14]), .I1(GND_net), .CO(n29716));
    SB_LUT4 add_639_9_lut (.I0(GND_net), .I1(n3048[7]), .I2(n3073[7]), 
            .I3(n27959), .O(duty_23__N_3740[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3795_16_lut (.I0(GND_net), .I1(n8242[13]), .I2(n1108_adj_4118), 
            .I3(n29714), .O(n8221[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3795_16 (.CI(n29714), .I0(n8242[13]), .I1(n1108_adj_4118), 
            .CO(n29715));
    SB_LUT4 add_3795_15_lut (.I0(GND_net), .I1(n8242[12]), .I2(n1035_adj_4119), 
            .I3(n29713), .O(n8221[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3795_15 (.CI(n29713), .I0(n8242[12]), .I1(n1035_adj_4119), 
            .CO(n29714));
    SB_LUT4 add_3795_14_lut (.I0(GND_net), .I1(n8242[11]), .I2(n962_adj_4120), 
            .I3(n29712), .O(n8221[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3795_14 (.CI(n29712), .I0(n8242[11]), .I1(n962_adj_4120), 
            .CO(n29713));
    SB_LUT4 add_3795_13_lut (.I0(GND_net), .I1(n8242[10]), .I2(n889_adj_4121), 
            .I3(n29711), .O(n8221[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3795_13 (.CI(n29711), .I0(n8242[10]), .I1(n889_adj_4121), 
            .CO(n29712));
    SB_LUT4 add_3795_12_lut (.I0(GND_net), .I1(n8242[9]), .I2(n816_adj_4122), 
            .I3(n29710), .O(n8221[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_639_9 (.CI(n27959), .I0(n3048[7]), .I1(n3073[7]), .CO(n27960));
    SB_CARRY add_3795_12 (.CI(n29710), .I0(n8242[9]), .I1(n816_adj_4122), 
            .CO(n29711));
    SB_LUT4 add_3795_11_lut (.I0(GND_net), .I1(n8242[8]), .I2(n743_adj_4123), 
            .I3(n29709), .O(n8221[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3795_11 (.CI(n29709), .I0(n8242[8]), .I1(n743_adj_4123), 
            .CO(n29710));
    SB_CARRY add_3772_15 (.CI(n29451), .I0(n7924[12]), .I1(n1032), .CO(n29452));
    SB_LUT4 add_3795_10_lut (.I0(GND_net), .I1(n8242[7]), .I2(n670_adj_4124), 
            .I3(n29708), .O(n8221[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3795_10 (.CI(n29708), .I0(n8242[7]), .I1(n670_adj_4124), 
            .CO(n29709));
    SB_LUT4 add_3795_9_lut (.I0(GND_net), .I1(n8242[6]), .I2(n597_adj_4125), 
            .I3(n29707), .O(n8221[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3795_9 (.CI(n29707), .I0(n8242[6]), .I1(n597_adj_4125), 
            .CO(n29708));
    SB_LUT4 add_639_8_lut (.I0(GND_net), .I1(n3048[6]), .I2(n3073[6]), 
            .I3(n27958), .O(duty_23__N_3740[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_639_8 (.CI(n27958), .I0(n3048[6]), .I1(n3073[6]), .CO(n27959));
    SB_LUT4 i22916_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n27563), .I3(n8140[0]), .O(n4_adj_4126));   // verilog/motorControl.v(42[17:23])
    defparam i22916_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_977 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(n8140[0]), .I3(n27563), .O(n8134[1]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_977.LUT_INIT = 16'h8778;
    SB_LUT4 i22903_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.err [19]), .I3(\Kp[1] ), .O(n8134[0]));   // verilog/motorControl.v(42[17:23])
    defparam i22903_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_3772_14_lut (.I0(GND_net), .I1(n7924[11]), .I2(n959), 
            .I3(n29450), .O(n7902[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3772_14 (.CI(n29450), .I0(n7924[11]), .I1(n959), .CO(n29451));
    SB_LUT4 add_3772_13_lut (.I0(GND_net), .I1(n7924[10]), .I2(n886), 
            .I3(n29449), .O(n7902[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3795_8_lut (.I0(GND_net), .I1(n8242[5]), .I2(n524_adj_4127), 
            .I3(n29706), .O(n8221[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3795_8 (.CI(n29706), .I0(n8242[5]), .I1(n524_adj_4127), 
            .CO(n29707));
    SB_LUT4 add_3795_7_lut (.I0(GND_net), .I1(n8242[4]), .I2(n451_adj_4128), 
            .I3(n29705), .O(n8221[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3795_7 (.CI(n29705), .I0(n8242[4]), .I1(n451_adj_4128), 
            .CO(n29706));
    SB_LUT4 add_3795_6_lut (.I0(GND_net), .I1(n8242[3]), .I2(n378_adj_4129), 
            .I3(n29704), .O(n8221[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3795_6 (.CI(n29704), .I0(n8242[3]), .I1(n378_adj_4129), 
            .CO(n29705));
    SB_LUT4 add_3795_5_lut (.I0(GND_net), .I1(n8242[2]), .I2(n305_adj_4130), 
            .I3(n29703), .O(n8221[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3795_5 (.CI(n29703), .I0(n8242[2]), .I1(n305_adj_4130), 
            .CO(n29704));
    SB_LUT4 add_3795_4_lut (.I0(GND_net), .I1(n8242[1]), .I2(n232_adj_4131), 
            .I3(n29702), .O(n8221[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3795_4 (.CI(n29702), .I0(n8242[1]), .I1(n232_adj_4131), 
            .CO(n29703));
    SB_LUT4 i22905_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(\PID_CONTROLLER.err [19]), .I3(\Kp[1] ), .O(n27563));   // verilog/motorControl.v(42[17:23])
    defparam i22905_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_3795_3_lut (.I0(GND_net), .I1(n8242[0]), .I2(n159_adj_4132), 
            .I3(n29701), .O(n8221[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3795_3 (.CI(n29701), .I0(n8242[0]), .I1(n159_adj_4132), 
            .CO(n29702));
    SB_LUT4 add_3795_2_lut (.I0(GND_net), .I1(n17_adj_4133), .I2(n86_adj_4134), 
            .I3(GND_net), .O(n8221[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3795_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3795_2 (.CI(GND_net), .I0(n17_adj_4133), .I1(n86_adj_4134), 
            .CO(n29701));
    SB_LUT4 add_3794_21_lut (.I0(GND_net), .I1(n8221[18]), .I2(GND_net), 
            .I3(n29700), .O(n8199[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3794_20_lut (.I0(GND_net), .I1(n8221[17]), .I2(GND_net), 
            .I3(n29699), .O(n8199[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3794_20 (.CI(n29699), .I0(n8221[17]), .I1(GND_net), .CO(n29700));
    SB_LUT4 add_639_7_lut (.I0(GND_net), .I1(n3048[5]), .I2(n3073[5]), 
            .I3(n27957), .O(duty_23__N_3740[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3794_19_lut (.I0(GND_net), .I1(n8221[16]), .I2(GND_net), 
            .I3(n29698), .O(n8199[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3794_19 (.CI(n29698), .I0(n8221[16]), .I1(GND_net), .CO(n29699));
    SB_LUT4 add_3794_18_lut (.I0(GND_net), .I1(n8221[15]), .I2(GND_net), 
            .I3(n29697), .O(n8199[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3794_18 (.CI(n29697), .I0(n8221[15]), .I1(GND_net), .CO(n29698));
    SB_LUT4 add_3794_17_lut (.I0(GND_net), .I1(n8221[14]), .I2(GND_net), 
            .I3(n29696), .O(n8199[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22947_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n27597), .I3(n8145[0]), .O(n4_adj_4135));   // verilog/motorControl.v(42[17:23])
    defparam i22947_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_CARRY add_639_7 (.CI(n27957), .I0(n3048[5]), .I1(n3073[5]), .CO(n27958));
    SB_CARRY add_3794_17 (.CI(n29696), .I0(n8221[14]), .I1(GND_net), .CO(n29697));
    SB_LUT4 add_3794_16_lut (.I0(GND_net), .I1(n8221[13]), .I2(n1105_adj_4136), 
            .I3(n29695), .O(n8199[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3794_16 (.CI(n29695), .I0(n8221[13]), .I1(n1105_adj_4136), 
            .CO(n29696));
    SB_CARRY add_3772_13 (.CI(n29449), .I0(n7924[10]), .I1(n886), .CO(n29450));
    SB_LUT4 add_3794_15_lut (.I0(GND_net), .I1(n8221[12]), .I2(n1032_adj_4137), 
            .I3(n29694), .O(n8199[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3794_15 (.CI(n29694), .I0(n8221[12]), .I1(n1032_adj_4137), 
            .CO(n29695));
    SB_LUT4 add_3794_14_lut (.I0(GND_net), .I1(n8221[11]), .I2(n959_adj_4138), 
            .I3(n29693), .O(n8199[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3794_14 (.CI(n29693), .I0(n8221[11]), .I1(n959_adj_4138), 
            .CO(n29694));
    SB_LUT4 add_3794_13_lut (.I0(GND_net), .I1(n8221[10]), .I2(n886_adj_4139), 
            .I3(n29692), .O(n8199[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3794_13 (.CI(n29692), .I0(n8221[10]), .I1(n886_adj_4139), 
            .CO(n29693));
    SB_LUT4 add_3794_12_lut (.I0(GND_net), .I1(n8221[9]), .I2(n813), .I3(n29691), 
            .O(n8199[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3794_12 (.CI(n29691), .I0(n8221[9]), .I1(n813), .CO(n29692));
    SB_LUT4 add_3794_11_lut (.I0(GND_net), .I1(n8221[8]), .I2(n740), .I3(n29690), 
            .O(n8199[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3794_11 (.CI(n29690), .I0(n8221[8]), .I1(n740), .CO(n29691));
    SB_LUT4 add_3794_10_lut (.I0(GND_net), .I1(n8221[7]), .I2(n667), .I3(n29689), 
            .O(n8199[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3794_10 (.CI(n29689), .I0(n8221[7]), .I1(n667), .CO(n29690));
    SB_LUT4 add_3794_9_lut (.I0(GND_net), .I1(n8221[6]), .I2(n594), .I3(n29688), 
            .O(n8199[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3794_9 (.CI(n29688), .I0(n8221[6]), .I1(n594), .CO(n29689));
    SB_LUT4 add_3794_8_lut (.I0(GND_net), .I1(n8221[5]), .I2(n521), .I3(n29687), 
            .O(n8199[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3794_8 (.CI(n29687), .I0(n8221[5]), .I1(n521), .CO(n29688));
    SB_LUT4 add_3794_7_lut (.I0(GND_net), .I1(n8221[4]), .I2(n448), .I3(n29686), 
            .O(n8199[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3794_7 (.CI(n29686), .I0(n8221[4]), .I1(n448), .CO(n29687));
    SB_LUT4 add_3794_6_lut (.I0(GND_net), .I1(n8221[3]), .I2(n375), .I3(n29685), 
            .O(n8199[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3794_6 (.CI(n29685), .I0(n8221[3]), .I1(n375), .CO(n29686));
    SB_LUT4 add_3772_12_lut (.I0(GND_net), .I1(n7924[9]), .I2(n813_adj_4140), 
            .I3(n29448), .O(n7902[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3794_5_lut (.I0(GND_net), .I1(n8221[2]), .I2(n302), .I3(n29684), 
            .O(n8199[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3794_5 (.CI(n29684), .I0(n8221[2]), .I1(n302), .CO(n29685));
    SB_LUT4 i2_3_lut_4_lut_adj_978 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [20]), 
            .I2(n8145[0]), .I3(n27597), .O(n8140[1]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_978.LUT_INIT = 16'h8778;
    SB_LUT4 add_3794_4_lut (.I0(GND_net), .I1(n8221[1]), .I2(n229), .I3(n29683), 
            .O(n8199[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3794_4 (.CI(n29683), .I0(n8221[1]), .I1(n229), .CO(n29684));
    SB_LUT4 i22934_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n8140[0]));   // verilog/motorControl.v(42[17:23])
    defparam i22934_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 add_3794_3_lut (.I0(GND_net), .I1(n8221[0]), .I2(n156), .I3(n29682), 
            .O(n8199[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3794_3 (.CI(n29682), .I0(n8221[0]), .I1(n156), .CO(n29683));
    SB_LUT4 add_3794_2_lut (.I0(GND_net), .I1(n14_adj_4141), .I2(n83), 
            .I3(GND_net), .O(n8199[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3794_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3794_2 (.CI(GND_net), .I0(n14_adj_4141), .I1(n83), .CO(n29682));
    SB_CARRY add_3772_12 (.CI(n29448), .I0(n7924[9]), .I1(n813_adj_4140), 
            .CO(n29449));
    SB_LUT4 add_3793_22_lut (.I0(GND_net), .I1(n8199[19]), .I2(GND_net), 
            .I3(n29681), .O(n8176[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3793_21_lut (.I0(GND_net), .I1(n8199[18]), .I2(GND_net), 
            .I3(n29680), .O(n8176[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_21 (.CI(n29680), .I0(n8199[18]), .I1(GND_net), .CO(n29681));
    SB_LUT4 add_3793_20_lut (.I0(GND_net), .I1(n8199[17]), .I2(GND_net), 
            .I3(n29679), .O(n8176[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_20 (.CI(n29679), .I0(n8199[17]), .I1(GND_net), .CO(n29680));
    SB_LUT4 add_3793_19_lut (.I0(GND_net), .I1(n8199[16]), .I2(GND_net), 
            .I3(n29678), .O(n8176[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_19 (.CI(n29678), .I0(n8199[16]), .I1(GND_net), .CO(n29679));
    SB_LUT4 add_3793_18_lut (.I0(GND_net), .I1(n8199[15]), .I2(GND_net), 
            .I3(n29677), .O(n8176[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_18 (.CI(n29677), .I0(n8199[15]), .I1(GND_net), .CO(n29678));
    SB_LUT4 i22936_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [21]), 
            .I2(\PID_CONTROLLER.err [20]), .I3(\Kp[1] ), .O(n27597));   // verilog/motorControl.v(42[17:23])
    defparam i22936_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 add_3793_17_lut (.I0(GND_net), .I1(n8199[14]), .I2(GND_net), 
            .I3(n29676), .O(n8176[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_17 (.CI(n29676), .I0(n8199[14]), .I1(GND_net), .CO(n29677));
    SB_LUT4 add_3793_16_lut (.I0(GND_net), .I1(n8199[13]), .I2(n1102_adj_4142), 
            .I3(n29675), .O(n8176[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_16 (.CI(n29675), .I0(n8199[13]), .I1(n1102_adj_4142), 
            .CO(n29676));
    SB_LUT4 add_3793_15_lut (.I0(GND_net), .I1(n8199[12]), .I2(n1029_adj_4143), 
            .I3(n29674), .O(n8176[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_15 (.CI(n29674), .I0(n8199[12]), .I1(n1029_adj_4143), 
            .CO(n29675));
    SB_LUT4 add_3793_14_lut (.I0(GND_net), .I1(n8199[11]), .I2(n956_adj_4144), 
            .I3(n29673), .O(n8176[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_14 (.CI(n29673), .I0(n8199[11]), .I1(n956_adj_4144), 
            .CO(n29674));
    SB_LUT4 add_3793_13_lut (.I0(GND_net), .I1(n8199[10]), .I2(n883_adj_4145), 
            .I3(n29672), .O(n8176[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3772_11_lut (.I0(GND_net), .I1(n7924[8]), .I2(n740_adj_4146), 
            .I3(n29447), .O(n7902[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_13 (.CI(n29672), .I0(n8199[10]), .I1(n883_adj_4145), 
            .CO(n29673));
    SB_LUT4 add_3793_12_lut (.I0(GND_net), .I1(n8199[9]), .I2(n810_adj_4147), 
            .I3(n29671), .O(n8176[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_12 (.CI(n29671), .I0(n8199[9]), .I1(n810_adj_4147), 
            .CO(n29672));
    SB_LUT4 add_3793_11_lut (.I0(GND_net), .I1(n8199[8]), .I2(n737_adj_4148), 
            .I3(n29670), .O(n8176[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_11 (.CI(n29670), .I0(n8199[8]), .I1(n737_adj_4148), 
            .CO(n29671));
    SB_LUT4 add_3793_10_lut (.I0(GND_net), .I1(n8199[7]), .I2(n664_adj_4149), 
            .I3(n29669), .O(n8176[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_10 (.CI(n29669), .I0(n8199[7]), .I1(n664_adj_4149), 
            .CO(n29670));
    SB_LUT4 add_3793_9_lut (.I0(GND_net), .I1(n8199[6]), .I2(n591_adj_4150), 
            .I3(n29668), .O(n8176[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_9 (.CI(n29668), .I0(n8199[6]), .I1(n591_adj_4150), 
            .CO(n29669));
    SB_CARRY add_3772_11 (.CI(n29447), .I0(n7924[8]), .I1(n740_adj_4146), 
            .CO(n29448));
    SB_LUT4 add_3793_8_lut (.I0(GND_net), .I1(n8199[5]), .I2(n518_adj_4151), 
            .I3(n29667), .O(n8176[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_8 (.CI(n29667), .I0(n8199[5]), .I1(n518_adj_4151), 
            .CO(n29668));
    SB_LUT4 add_3793_7_lut (.I0(GND_net), .I1(n8199[4]), .I2(n445_adj_4152), 
            .I3(n29666), .O(n8176[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_7 (.CI(n29666), .I0(n8199[4]), .I1(n445_adj_4152), 
            .CO(n29667));
    SB_LUT4 add_3793_6_lut (.I0(GND_net), .I1(n8199[3]), .I2(n372_adj_4153), 
            .I3(n29665), .O(n8176[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_6 (.CI(n29665), .I0(n8199[3]), .I1(n372_adj_4153), 
            .CO(n29666));
    SB_LUT4 add_3793_5_lut (.I0(GND_net), .I1(n8199[2]), .I2(n299_adj_4154), 
            .I3(n29664), .O(n8176[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_5 (.CI(n29664), .I0(n8199[2]), .I1(n299_adj_4154), 
            .CO(n29665));
    SB_LUT4 add_3793_4_lut (.I0(GND_net), .I1(n8199[1]), .I2(n226_adj_4155), 
            .I3(n29663), .O(n8176[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_4 (.CI(n29663), .I0(n8199[1]), .I1(n226_adj_4155), 
            .CO(n29664));
    SB_LUT4 add_3793_3_lut (.I0(GND_net), .I1(n8199[0]), .I2(n153_adj_4156), 
            .I3(n29662), .O(n8176[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_3 (.CI(n29662), .I0(n8199[0]), .I1(n153_adj_4156), 
            .CO(n29663));
    SB_LUT4 add_3793_2_lut (.I0(GND_net), .I1(n11_adj_4157), .I2(n80_adj_4158), 
            .I3(GND_net), .O(n8176[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3793_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3793_2 (.CI(GND_net), .I0(n11_adj_4157), .I1(n80_adj_4158), 
            .CO(n29662));
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral [23]), .I1(n8152[21]), 
            .I2(GND_net), .I3(n29661), .O(n40677)) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_3772_10_lut (.I0(GND_net), .I1(n7924[7]), .I2(n667_adj_4159), 
            .I3(n29446), .O(n7902[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n8152[20]), .I2(GND_net), 
            .I3(n29660), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_23 (.CI(n29660), .I0(n8152[20]), .I1(GND_net), 
            .CO(n29661));
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n8152[19]), .I2(GND_net), 
            .I3(n29659), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_22 (.CI(n29659), .I0(n8152[19]), .I1(GND_net), 
            .CO(n29660));
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n8152[18]), .I2(GND_net), 
            .I3(n29658), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_21 (.CI(n29658), .I0(n8152[18]), .I1(GND_net), 
            .CO(n29659));
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n8152[17]), .I2(GND_net), 
            .I3(n29657), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_20 (.CI(n29657), .I0(n8152[17]), .I1(GND_net), 
            .CO(n29658));
    SB_CARRY add_3772_10 (.CI(n29446), .I0(n7924[7]), .I1(n667_adj_4159), 
            .CO(n29447));
    SB_LUT4 add_3772_9_lut (.I0(GND_net), .I1(n7924[6]), .I2(n594_adj_4161), 
            .I3(n29445), .O(n7902[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n8152[16]), .I2(GND_net), 
            .I3(n29656), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_19 (.CI(n29656), .I0(n8152[16]), .I1(GND_net), 
            .CO(n29657));
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n8152[15]), .I2(GND_net), 
            .I3(n29655), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_18 (.CI(n29655), .I0(n8152[15]), .I1(GND_net), 
            .CO(n29656));
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n8152[14]), .I2(GND_net), 
            .I3(n29654), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_17 (.CI(n29654), .I0(n8152[14]), .I1(GND_net), 
            .CO(n29655));
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n8152[13]), .I2(n1096_adj_4163), 
            .I3(n29653), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_16 (.CI(n29653), .I0(n8152[13]), .I1(n1096_adj_4163), 
            .CO(n29654));
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n8152[12]), .I2(n1023_adj_4165), 
            .I3(n29652), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3772_9 (.CI(n29445), .I0(n7924[6]), .I1(n594_adj_4161), 
            .CO(n29446));
    SB_CARRY mult_11_add_1225_15 (.CI(n29652), .I0(n8152[12]), .I1(n1023_adj_4165), 
            .CO(n29653));
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n8152[11]), .I2(n950_adj_4166), 
            .I3(n29651), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_14 (.CI(n29651), .I0(n8152[11]), .I1(n950_adj_4166), 
            .CO(n29652));
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n8152[10]), .I2(n877_adj_4167), 
            .I3(n29650), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_13 (.CI(n29650), .I0(n8152[10]), .I1(n877_adj_4167), 
            .CO(n29651));
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n8152[9]), .I2(n804_adj_4169), 
            .I3(n29649), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_12 (.CI(n29649), .I0(n8152[9]), .I1(n804_adj_4169), 
            .CO(n29650));
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n8152[8]), .I2(n731_adj_4170), 
            .I3(n29648), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_11 (.CI(n29648), .I0(n8152[8]), .I1(n731_adj_4170), 
            .CO(n29649));
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n8152[7]), .I2(n658_adj_4171), 
            .I3(n29647), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n29647), .I0(n8152[7]), .I1(n658_adj_4171), 
            .CO(n29648));
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n8152[6]), .I2(n585_adj_4173), 
            .I3(n29646), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3772_8_lut (.I0(GND_net), .I1(n7924[5]), .I2(n521_adj_4174), 
            .I3(n29444), .O(n7902[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_9 (.CI(n29646), .I0(n8152[6]), .I1(n585_adj_4173), 
            .CO(n29647));
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n8152[5]), .I2(n512_adj_4175), 
            .I3(n29645), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_8 (.CI(n29645), .I0(n8152[5]), .I1(n512_adj_4175), 
            .CO(n29646));
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n8152[4]), .I2(n439_adj_4176), 
            .I3(n29644), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_7 (.CI(n29644), .I0(n8152[4]), .I1(n439_adj_4176), 
            .CO(n29645));
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n8152[3]), .I2(n366_adj_4178), 
            .I3(n29643), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_6 (.CI(n29643), .I0(n8152[3]), .I1(n366_adj_4178), 
            .CO(n29644));
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n8152[2]), .I2(n293_adj_4179), 
            .I3(n29642), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_5 (.CI(n29642), .I0(n8152[2]), .I1(n293_adj_4179), 
            .CO(n29643));
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n8152[1]), .I2(n220_adj_4180), 
            .I3(n29641), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3772_8 (.CI(n29444), .I0(n7924[5]), .I1(n521_adj_4174), 
            .CO(n29445));
    SB_CARRY mult_11_add_1225_4 (.CI(n29641), .I0(n8152[1]), .I1(n220_adj_4180), 
            .CO(n29642));
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n8152[0]), .I2(n147_adj_4181), 
            .I3(n29640), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n29640), .I0(n8152[0]), .I1(n147_adj_4181), 
            .CO(n29641));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4182), .I2(n74_adj_4183), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_4182), .I1(n74_adj_4183), 
            .CO(n29640));
    SB_LUT4 add_3792_23_lut (.I0(GND_net), .I1(n8176[20]), .I2(GND_net), 
            .I3(n29639), .O(n8152[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3792_22_lut (.I0(GND_net), .I1(n8176[19]), .I2(GND_net), 
            .I3(n29638), .O(n8152[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_22 (.CI(n29638), .I0(n8176[19]), .I1(GND_net), .CO(n29639));
    SB_LUT4 add_3792_21_lut (.I0(GND_net), .I1(n8176[18]), .I2(GND_net), 
            .I3(n29637), .O(n8152[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_21 (.CI(n29637), .I0(n8176[18]), .I1(GND_net), .CO(n29638));
    SB_LUT4 add_3792_20_lut (.I0(GND_net), .I1(n8176[17]), .I2(GND_net), 
            .I3(n29636), .O(n8152[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_20 (.CI(n29636), .I0(n8176[17]), .I1(GND_net), .CO(n29637));
    SB_LUT4 add_3792_19_lut (.I0(GND_net), .I1(n8176[16]), .I2(GND_net), 
            .I3(n29635), .O(n8152[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_19 (.CI(n29635), .I0(n8176[16]), .I1(GND_net), .CO(n29636));
    SB_LUT4 add_3792_18_lut (.I0(GND_net), .I1(n8176[15]), .I2(GND_net), 
            .I3(n29634), .O(n8152[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_18 (.CI(n29634), .I0(n8176[15]), .I1(GND_net), .CO(n29635));
    SB_LUT4 add_3792_17_lut (.I0(GND_net), .I1(n8176[14]), .I2(GND_net), 
            .I3(n29633), .O(n8152[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_17 (.CI(n29633), .I0(n8176[14]), .I1(GND_net), .CO(n29634));
    SB_LUT4 add_3792_16_lut (.I0(GND_net), .I1(n8176[13]), .I2(n1099_adj_4184), 
            .I3(n29632), .O(n8152[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_16 (.CI(n29632), .I0(n8176[13]), .I1(n1099_adj_4184), 
            .CO(n29633));
    SB_LUT4 add_3792_15_lut (.I0(GND_net), .I1(n8176[12]), .I2(n1026_adj_4185), 
            .I3(n29631), .O(n8152[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_15 (.CI(n29631), .I0(n8176[12]), .I1(n1026_adj_4185), 
            .CO(n29632));
    SB_LUT4 add_3792_14_lut (.I0(GND_net), .I1(n8176[11]), .I2(n953_adj_4186), 
            .I3(n29630), .O(n8152[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_14 (.CI(n29630), .I0(n8176[11]), .I1(n953_adj_4186), 
            .CO(n29631));
    SB_LUT4 add_3772_7_lut (.I0(GND_net), .I1(n7924[4]), .I2(n448_adj_4187), 
            .I3(n29443), .O(n7902[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3792_13_lut (.I0(GND_net), .I1(n8176[10]), .I2(n880_adj_4188), 
            .I3(n29629), .O(n8152[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_13 (.CI(n29629), .I0(n8176[10]), .I1(n880_adj_4188), 
            .CO(n29630));
    SB_CARRY add_3772_7 (.CI(n29443), .I0(n7924[4]), .I1(n448_adj_4187), 
            .CO(n29444));
    SB_LUT4 add_639_6_lut (.I0(GND_net), .I1(n3048[4]), .I2(n3073[4]), 
            .I3(n27956), .O(duty_23__N_3740[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3792_12_lut (.I0(GND_net), .I1(n8176[9]), .I2(n807_adj_4189), 
            .I3(n29628), .O(n8152[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3772_6_lut (.I0(GND_net), .I1(n7924[3]), .I2(n375_adj_4190), 
            .I3(n29442), .O(n7902[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_12 (.CI(n29628), .I0(n8176[9]), .I1(n807_adj_4189), 
            .CO(n29629));
    SB_LUT4 add_3792_11_lut (.I0(GND_net), .I1(n8176[8]), .I2(n734_adj_4191), 
            .I3(n29627), .O(n8152[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_11 (.CI(n29627), .I0(n8176[8]), .I1(n734_adj_4191), 
            .CO(n29628));
    SB_CARRY add_639_6 (.CI(n27956), .I0(n3048[4]), .I1(n3073[4]), .CO(n27957));
    SB_LUT4 add_3792_10_lut (.I0(GND_net), .I1(n8176[7]), .I2(n661_adj_4192), 
            .I3(n29626), .O(n8152[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_10 (.CI(n29626), .I0(n8176[7]), .I1(n661_adj_4192), 
            .CO(n29627));
    SB_LUT4 add_3792_9_lut (.I0(GND_net), .I1(n8176[6]), .I2(n588_adj_4193), 
            .I3(n29625), .O(n8152[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_9 (.CI(n29625), .I0(n8176[6]), .I1(n588_adj_4193), 
            .CO(n29626));
    SB_LUT4 add_3792_8_lut (.I0(GND_net), .I1(n8176[5]), .I2(n515_adj_4194), 
            .I3(n29624), .O(n8152[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_8 (.CI(n29624), .I0(n8176[5]), .I1(n515_adj_4194), 
            .CO(n29625));
    SB_CARRY add_3772_6 (.CI(n29442), .I0(n7924[3]), .I1(n375_adj_4190), 
            .CO(n29443));
    SB_LUT4 add_3792_7_lut (.I0(GND_net), .I1(n8176[4]), .I2(n442_adj_4195), 
            .I3(n29623), .O(n8152[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3772_5_lut (.I0(GND_net), .I1(n7924[2]), .I2(n302_adj_4196), 
            .I3(n29441), .O(n7902[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3772_5 (.CI(n29441), .I0(n7924[2]), .I1(n302_adj_4196), 
            .CO(n29442));
    SB_LUT4 add_3772_4_lut (.I0(GND_net), .I1(n7924[1]), .I2(n229_adj_4197), 
            .I3(n29440), .O(n7902[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3772_4 (.CI(n29440), .I0(n7924[1]), .I1(n229_adj_4197), 
            .CO(n29441));
    SB_CARRY add_3792_7 (.CI(n29623), .I0(n8176[4]), .I1(n442_adj_4195), 
            .CO(n29624));
    SB_LUT4 add_3792_6_lut (.I0(GND_net), .I1(n8176[3]), .I2(n369_adj_4198), 
            .I3(n29622), .O(n8152[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_6 (.CI(n29622), .I0(n8176[3]), .I1(n369_adj_4198), 
            .CO(n29623));
    SB_LUT4 add_3792_5_lut (.I0(GND_net), .I1(n8176[2]), .I2(n296_adj_4199), 
            .I3(n29621), .O(n8152[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_5 (.CI(n29621), .I0(n8176[2]), .I1(n296_adj_4199), 
            .CO(n29622));
    SB_LUT4 add_3792_4_lut (.I0(GND_net), .I1(n8176[1]), .I2(n223_adj_4200), 
            .I3(n29620), .O(n8152[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_4 (.CI(n29620), .I0(n8176[1]), .I1(n223_adj_4200), 
            .CO(n29621));
    SB_LUT4 add_3792_3_lut (.I0(GND_net), .I1(n8176[0]), .I2(n150_adj_4201), 
            .I3(n29619), .O(n8152[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_3 (.CI(n29619), .I0(n8176[0]), .I1(n150_adj_4201), 
            .CO(n29620));
    SB_LUT4 add_3792_2_lut (.I0(GND_net), .I1(n8_adj_4202), .I2(n77_adj_4203), 
            .I3(GND_net), .O(n8152[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3792_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3792_2 (.CI(GND_net), .I0(n8_adj_4202), .I1(n77_adj_4203), 
            .CO(n29619));
    SB_LUT4 add_3786_7_lut (.I0(GND_net), .I1(n37305), .I2(n490_adj_4204), 
            .I3(n29618), .O(n8119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3786_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3786_6_lut (.I0(GND_net), .I1(n8127[3]), .I2(n417_adj_4205), 
            .I3(n29617), .O(n8119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3786_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3786_6 (.CI(n29617), .I0(n8127[3]), .I1(n417_adj_4205), 
            .CO(n29618));
    SB_LUT4 add_3786_5_lut (.I0(GND_net), .I1(n8127[2]), .I2(n344_adj_4206), 
            .I3(n29616), .O(n8119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3786_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3786_5 (.CI(n29616), .I0(n8127[2]), .I1(n344_adj_4206), 
            .CO(n29617));
    SB_LUT4 add_3786_4_lut (.I0(GND_net), .I1(n8127[1]), .I2(n271_adj_4207), 
            .I3(n29615), .O(n8119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3786_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3786_4 (.CI(n29615), .I0(n8127[1]), .I1(n271_adj_4207), 
            .CO(n29616));
    SB_LUT4 add_3786_3_lut (.I0(GND_net), .I1(n8127[0]), .I2(n198_adj_4208), 
            .I3(n29614), .O(n8119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3786_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3786_3 (.CI(n29614), .I0(n8127[0]), .I1(n198_adj_4208), 
            .CO(n29615));
    SB_LUT4 add_3786_2_lut (.I0(GND_net), .I1(n56_adj_4209), .I2(n125_adj_4210), 
            .I3(GND_net), .O(n8119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3786_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3786_2 (.CI(GND_net), .I0(n56_adj_4209), .I1(n125_adj_4210), 
            .CO(n29614));
    SB_LUT4 add_3785_8_lut (.I0(GND_net), .I1(n8119[5]), .I2(n560_adj_4211), 
            .I3(n29613), .O(n8110[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3785_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3785_7_lut (.I0(GND_net), .I1(n8119[4]), .I2(n487_adj_4212), 
            .I3(n29612), .O(n8110[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3785_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3785_7 (.CI(n29612), .I0(n8119[4]), .I1(n487_adj_4212), 
            .CO(n29613));
    SB_LUT4 add_3785_6_lut (.I0(GND_net), .I1(n8119[3]), .I2(n414_adj_4213), 
            .I3(n29611), .O(n8110[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3785_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3785_6 (.CI(n29611), .I0(n8119[3]), .I1(n414_adj_4213), 
            .CO(n29612));
    SB_LUT4 add_3772_3_lut (.I0(GND_net), .I1(n7924[0]), .I2(n156_adj_4214), 
            .I3(n29439), .O(n7902[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3785_5_lut (.I0(GND_net), .I1(n8119[2]), .I2(n341_adj_4215), 
            .I3(n29610), .O(n8110[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3785_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3772_3 (.CI(n29439), .I0(n7924[0]), .I1(n156_adj_4214), 
            .CO(n29440));
    SB_CARRY add_3785_5 (.CI(n29610), .I0(n8119[2]), .I1(n341_adj_4215), 
            .CO(n29611));
    SB_LUT4 add_3785_4_lut (.I0(GND_net), .I1(n8119[1]), .I2(n268_adj_4216), 
            .I3(n29609), .O(n8110[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3785_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3785_4 (.CI(n29609), .I0(n8119[1]), .I1(n268_adj_4216), 
            .CO(n29610));
    SB_LUT4 add_3772_2_lut (.I0(GND_net), .I1(n14_adj_4217), .I2(n83_adj_4218), 
            .I3(GND_net), .O(n7902[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3772_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3772_2 (.CI(GND_net), .I0(n14_adj_4217), .I1(n83_adj_4218), 
            .CO(n29439));
    SB_LUT4 add_3785_3_lut (.I0(GND_net), .I1(n8119[0]), .I2(n195_adj_4219), 
            .I3(n29608), .O(n8110[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3785_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3785_3 (.CI(n29608), .I0(n8119[0]), .I1(n195_adj_4219), 
            .CO(n29609));
    SB_LUT4 add_3785_2_lut (.I0(GND_net), .I1(n53_adj_4220), .I2(n122_adj_4221), 
            .I3(GND_net), .O(n8110[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3785_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3785_2 (.CI(GND_net), .I0(n53_adj_4220), .I1(n122_adj_4221), 
            .CO(n29608));
    SB_LUT4 add_3784_9_lut (.I0(GND_net), .I1(n8110[6]), .I2(n630_adj_4222), 
            .I3(n29607), .O(n8100[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3784_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3784_8_lut (.I0(GND_net), .I1(n8110[5]), .I2(n557_adj_4223), 
            .I3(n29606), .O(n8100[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3784_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3784_8 (.CI(n29606), .I0(n8110[5]), .I1(n557_adj_4223), 
            .CO(n29607));
    SB_LUT4 add_639_5_lut (.I0(GND_net), .I1(n3048[3]), .I2(n3073[3]), 
            .I3(n27955), .O(duty_23__N_3740[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_639_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3784_7_lut (.I0(GND_net), .I1(n8110[4]), .I2(n484_adj_4224), 
            .I3(n29605), .O(n8100[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3784_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3784_7 (.CI(n29605), .I0(n8110[4]), .I1(n484_adj_4224), 
            .CO(n29606));
    SB_LUT4 add_3784_6_lut (.I0(GND_net), .I1(n8110[3]), .I2(n411_adj_4225), 
            .I3(n29604), .O(n8100[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3784_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3784_6 (.CI(n29604), .I0(n8110[3]), .I1(n411_adj_4225), 
            .CO(n29605));
    SB_LUT4 add_3784_5_lut (.I0(GND_net), .I1(n8110[2]), .I2(n338_adj_4226), 
            .I3(n29603), .O(n8100[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3784_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3784_5 (.CI(n29603), .I0(n8110[2]), .I1(n338_adj_4226), 
            .CO(n29604));
    SB_LUT4 add_3784_4_lut (.I0(GND_net), .I1(n8110[1]), .I2(n265_adj_4227), 
            .I3(n29602), .O(n8100[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3784_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3784_4 (.CI(n29602), .I0(n8110[1]), .I1(n265_adj_4227), 
            .CO(n29603));
    SB_LUT4 add_3784_3_lut (.I0(GND_net), .I1(n8110[0]), .I2(n192_adj_4228), 
            .I3(n29601), .O(n8100[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3784_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3784_3 (.CI(n29601), .I0(n8110[0]), .I1(n192_adj_4228), 
            .CO(n29602));
    SB_LUT4 add_3784_2_lut (.I0(GND_net), .I1(n50_adj_4229), .I2(n119_adj_4230), 
            .I3(GND_net), .O(n8100[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3784_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3784_2 (.CI(GND_net), .I0(n50_adj_4229), .I1(n119_adj_4230), 
            .CO(n29601));
    SB_LUT4 add_3783_10_lut (.I0(GND_net), .I1(n8100[7]), .I2(n700_adj_4231), 
            .I3(n29600), .O(n8089[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3783_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_3783_9_lut (.I0(GND_net), .I1(n8100[6]), .I2(n627_adj_4232), 
            .I3(n29599), .O(n8089[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3783_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3783_9 (.CI(n29599), .I0(n8100[6]), .I1(n627_adj_4232), 
            .CO(n29600));
    SB_LUT4 add_3783_8_lut (.I0(GND_net), .I1(n8100[5]), .I2(n554_adj_4233), 
            .I3(n29598), .O(n8089[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3783_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3783_8 (.CI(n29598), .I0(n8100[5]), .I1(n554_adj_4233), 
            .CO(n29599));
    SB_LUT4 add_3783_7_lut (.I0(GND_net), .I1(n8100[4]), .I2(n481_adj_4234), 
            .I3(n29597), .O(n8089[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3783_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3783_7 (.CI(n29597), .I0(n8100[4]), .I1(n481_adj_4234), 
            .CO(n29598));
    SB_LUT4 add_3783_6_lut (.I0(GND_net), .I1(n8100[3]), .I2(n408_adj_4235), 
            .I3(n29596), .O(n8089[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3783_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3783_6 (.CI(n29596), .I0(n8100[3]), .I1(n408_adj_4235), 
            .CO(n29597));
    SB_LUT4 add_3783_5_lut (.I0(GND_net), .I1(n8100[2]), .I2(n335_adj_4236), 
            .I3(n29595), .O(n8089[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3783_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3783_5 (.CI(n29595), .I0(n8100[2]), .I1(n335_adj_4236), 
            .CO(n29596));
    SB_LUT4 add_3783_4_lut (.I0(GND_net), .I1(n8100[1]), .I2(n262_adj_4237), 
            .I3(n29594), .O(n8089[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3783_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3783_4 (.CI(n29594), .I0(n8100[1]), .I1(n262_adj_4237), 
            .CO(n29595));
    SB_CARRY add_639_5 (.CI(n27955), .I0(n3048[3]), .I1(n3073[3]), .CO(n27956));
    SB_LUT4 add_3783_3_lut (.I0(GND_net), .I1(n8100[0]), .I2(n189_adj_4238), 
            .I3(n29593), .O(n8089[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3783_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3783_3 (.CI(n29593), .I0(n8100[0]), .I1(n189_adj_4238), 
            .CO(n29594));
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty[4]), .I1(n257[4]), .I2(GND_net), 
            .I3(GND_net), .O(n9_adj_3926));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty[5]), .I1(n257[5]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_3930));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty[6]), .I1(n257[6]), .I2(GND_net), 
            .I3(GND_net), .O(n13_adj_3929));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty[7]), .I1(n257[7]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_3928));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty[10]), .I1(n257[10]), .I2(GND_net), 
            .I3(GND_net), .O(n21_adj_3923));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty[9]), .I1(n257[9]), .I2(GND_net), 
            .I3(GND_net), .O(n19_adj_3924));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i22885_3_lut_4_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n4_adj_4239), .I3(n8134[1]), .O(n6_adj_4240));   // verilog/motorControl.v(42[17:23])
    defparam i22885_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty[8]), .I1(n257[8]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_3925));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty[11]), .I1(n257[11]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_3942));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty[12]), .I1(n257[12]), .I2(GND_net), 
            .I3(GND_net), .O(n25_adj_3941));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty[13]), .I1(n257[13]), .I2(GND_net), 
            .I3(GND_net), .O(n27_adj_3927));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty[14]), .I1(n257[14]), .I2(GND_net), 
            .I3(GND_net), .O(n29_adj_3944));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty[16]), .I1(n257[16]), .I2(GND_net), 
            .I3(GND_net), .O(n33_adj_3931));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty[15]), .I1(n257[15]), .I2(GND_net), 
            .I3(GND_net), .O(n31_adj_3943));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty[17]), .I1(n257[17]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_3934));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty[18]), .I1(n257[18]), .I2(GND_net), 
            .I3(GND_net), .O(n37_adj_3945));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty[19]), .I1(n257[19]), .I2(GND_net), 
            .I3(GND_net), .O(n39_adj_3952));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty[21]), .I1(n257[21]), .I2(GND_net), 
            .I3(GND_net), .O(n43_adj_3946));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty[20]), .I1(n257[20]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_3953));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189_adj_4238));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_4237));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335_adj_4236));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_3_lut_4_lut_adj_979 (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n8134[1]), .I3(n4_adj_4239), .O(n8127[2]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_979.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408_adj_4235));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481_adj_4234));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554_adj_4233));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627_adj_4232));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700_adj_4231));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_4230));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_4229));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_4228));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_4227));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_4226));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_4225));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_4224));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i4_3_lut (.I0(n155[3]), .I1(n1_adj_4253[3]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[3]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_4223));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630_adj_4222));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_4221));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53_adj_4220));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195_adj_4219));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83_adj_4218));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4217));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_4216));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341_adj_4215));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156_adj_4214));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414_adj_4213));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487_adj_4212));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560_adj_4211));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_4210));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56_adj_4209));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198_adj_4208));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_4207));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344_adj_4206));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417_adj_4205));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n6_adj_4240), .I1(\Kp[4] ), .I2(n8134[2]), .I3(\PID_CONTROLLER.err [18]), 
            .O(n8127[3]));   // verilog/motorControl.v(42[17:23])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 i2_4_lut_adj_980 (.I0(n4_adj_4126), .I1(\Kp[3] ), .I2(n8140[1]), 
            .I3(\PID_CONTROLLER.err [19]), .O(n8134[2]));   // verilog/motorControl.v(42[17:23])
    defparam i2_4_lut_adj_980.LUT_INIT = 16'h965a;
    SB_LUT4 i22957_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n8145[0]));   // verilog/motorControl.v(42[17:23])
    defparam i22957_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[5]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490_adj_4204));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_981 (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [23]), 
            .I3(\PID_CONTROLLER.err [22]), .O(n12_adj_4241));   // verilog/motorControl.v(42[17:23])
    defparam i2_4_lut_adj_981.LUT_INIT = 16'h9c50;
    SB_LUT4 i22924_4_lut (.I0(n8140[1]), .I1(\Kp[3] ), .I2(n4_adj_4126), 
            .I3(\PID_CONTROLLER.err [19]), .O(n6_adj_4242));   // verilog/motorControl.v(42[17:23])
    defparam i22924_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(\PID_CONTROLLER.err [19]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n11_adj_4243));   // verilog/motorControl.v(42[17:23])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i22893_4_lut (.I0(n8134[2]), .I1(\Kp[4] ), .I2(n6_adj_4240), 
            .I3(\PID_CONTROLLER.err [18]), .O(n8_adj_4244));   // verilog/motorControl.v(42[17:23])
    defparam i22893_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i22959_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(\PID_CONTROLLER.err [22]), 
            .I3(\PID_CONTROLLER.err [21]), .O(n27622));   // verilog/motorControl.v(42[17:23])
    defparam i22959_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut (.I0(n8_adj_4244), .I1(n11_adj_4243), .I2(n6_adj_4242), 
            .I3(n12_adj_4241), .O(n18_adj_4245));   // verilog/motorControl.v(42[17:23])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut (.I0(\Kp[5] ), .I1(\Kp[3] ), .I2(\PID_CONTROLLER.err [18]), 
            .I3(\PID_CONTROLLER.err [20]), .O(n13_adj_4246));   // verilog/motorControl.v(42[17:23])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut (.I0(n13_adj_4246), .I1(n18_adj_4245), .I2(n27622), 
            .I3(n4_adj_4135), .O(n37305));   // verilog/motorControl.v(42[17:23])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77_adj_4203));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4202));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150_adj_4201));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223_adj_4200));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_4199));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_4198));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229_adj_4197));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302_adj_4196));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_4195));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_4194));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588_adj_4193));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661_adj_4192));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734_adj_4191));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[6]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_3_lut_4_lut_adj_982 (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n8134[0]), .I3(n27520), .O(n8127[1]));   // verilog/motorControl.v(42[17:23])
    defparam i2_3_lut_4_lut_adj_982.LUT_INIT = 16'h8778;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375_adj_4190));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22877_3_lut_4_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [18]), 
            .I2(n27520), .I3(n8134[0]), .O(n4_adj_4239));   // verilog/motorControl.v(42[17:23])
    defparam i22877_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807_adj_4189));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i5_3_lut (.I0(n155[4]), .I1(n1_adj_4253[4]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[4]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880_adj_4188));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_4187));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953_adj_4186));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026_adj_4185));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099_adj_4184));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74_adj_4183));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[7]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4182));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147_adj_4181));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_4180));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_4179));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_4178));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_4176));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_4175));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22866_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n27520));   // verilog/motorControl.v(42[17:23])
    defparam i22866_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_4174));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[8]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585_adj_4173));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[9]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658_adj_4171));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i22864_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [19]), 
            .I2(\PID_CONTROLLER.err [18]), .I3(\Kp[1] ), .O(n8127[0]));   // verilog/motorControl.v(42[17:23])
    defparam i22864_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731_adj_4170));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804_adj_4169));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[10]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877_adj_4167));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950_adj_4166));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023_adj_4165));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096_adj_4163));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[11]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[12]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594_adj_4161));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[13]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667_adj_4159));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80_adj_4158));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4157));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153_adj_4156));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226_adj_4155));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_4154));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_4153));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_4152));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_4151));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591_adj_4150));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664_adj_4149));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737_adj_4148));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810_adj_4147));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_4146));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883_adj_4145));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956_adj_4144));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029_adj_4143));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102_adj_4142));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4141));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_3907));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[14]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813_adj_4140));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_4139));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_4138));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_4137));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_4136));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i6_3_lut (.I0(n155[5]), .I1(n1_adj_4253[5]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[5]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_4134));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4133));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_4132));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_4131));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_4130));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4129));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_4128));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_4127));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[15]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_3904));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i7_3_lut (.I0(n155[6]), .I1(n1_adj_4253[6]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[6]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597_adj_4125));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670_adj_4124));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743_adj_4123));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816_adj_4122));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889_adj_4121));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962_adj_4120));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035_adj_4119));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108_adj_4118));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i8_3_lut (.I0(n155[7]), .I1(n1_adj_4253[7]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[7]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_4117));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4116));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4115));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4114));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4113));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36808_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n43653));   // verilog/motorControl.v(37[14] 56[8])
    defparam i36808_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_4112));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_4111));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_4110));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600_adj_4109));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673_adj_4108));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746_adj_4107));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819_adj_4106));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892_adj_4105));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965_adj_4104));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i9_3_lut (.I0(n155[8]), .I1(n1_adj_4253[8]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[8]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038_adj_4103));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111_adj_4102));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92_adj_4101));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4100));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165_adj_4099));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238_adj_4098));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i10_3_lut (.I0(n155[9]), .I1(n1_adj_4253[9]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[9]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311_adj_4097));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384_adj_4096));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457_adj_4095));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530_adj_4094));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603_adj_4093));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676_adj_4092));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749_adj_4091));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822_adj_4090));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895_adj_4089));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968_adj_4088));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041_adj_4087));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114_adj_4086));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i11_3_lut (.I0(n155[10]), .I1(n1_adj_4253[10]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[10]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95_adj_4085));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4084));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168_adj_4083));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241_adj_4082));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_4081));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_4080));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_4079));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_4078));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_4077));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i12_3_lut (.I0(n155[11]), .I1(n1_adj_4253[11]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[11]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679_adj_4076));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752_adj_4075));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825_adj_4074));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898_adj_4073));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_4072));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i13_3_lut (.I0(n155[12]), .I1(n1_adj_4253[12]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[12]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044_adj_4071));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117_adj_4070));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_4069));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4068));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i14_3_lut (.I0(n155[13]), .I1(n1_adj_4253[13]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[13]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34264_3_lut_4_lut (.I0(duty[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty[2]), .O(n41111));   // verilog/motorControl.v(46[19:35])
    defparam i34264_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(GND_net), .O(n6_adj_3948));   // verilog/motorControl.v(46[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_4067));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_4066));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317_adj_4065));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_4064));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_4063));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536_adj_4062));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609_adj_4061));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682_adj_4060));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i15_3_lut (.I0(n155[14]), .I1(n1_adj_4253[14]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[14]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755_adj_4059));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828_adj_4058));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901_adj_4057));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974_adj_4056));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047_adj_4055));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120_adj_4054));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_4053));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_4052));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_4051));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_4050));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_4049));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_4048));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i1_1_lut (.I0(setpoint[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[0]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_4046));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_4045));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i2_1_lut (.I0(setpoint[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[1]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i3_1_lut (.I0(setpoint[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[2]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612_adj_4042));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685_adj_4041));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758_adj_4040));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i4_1_lut (.I0(setpoint[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[3]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831_adj_4038));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_4037));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i5_1_lut (.I0(setpoint[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[4]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977_adj_4035));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050_adj_4034));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i6_1_lut (.I0(setpoint[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[5]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i7_1_lut (.I0(setpoint[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[6]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_4031));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4030));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i8_1_lut (.I0(setpoint[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[7]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177_adj_4028));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i9_1_lut (.I0(setpoint[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[8]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_4026));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_4025));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i10_1_lut (.I0(setpoint[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[9]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_4023));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i11_1_lut (.I0(setpoint[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[10]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_4021));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i12_1_lut (.I0(setpoint[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[11]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542_adj_4019));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615_adj_4018));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i13_1_lut (.I0(setpoint[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[12]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688_adj_4016));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761_adj_4015));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i14_1_lut (.I0(setpoint[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[13]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834_adj_4013));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i16_3_lut (.I0(n155[15]), .I1(n1_adj_4253[15]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[15]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907_adj_4012));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980_adj_4011));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107_adj_4010));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38_adj_4009));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180_adj_4008));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253_adj_4007));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_4006));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_4005));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_4004));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_4003));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618_adj_4002));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691_adj_4001));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i15_1_lut (.I0(setpoint[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[14]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764_adj_3999));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837_adj_3998));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i16_1_lut (.I0(setpoint[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[15]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910_adj_3996));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i17_1_lut (.I0(setpoint[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[16]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i18_1_lut (.I0(setpoint[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[17]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_3993));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_3992));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_3991));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256_adj_3990));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329_adj_3989));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i19_1_lut (.I0(setpoint[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[18]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402_adj_3987));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475_adj_3986));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548_adj_3985));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621_adj_3984));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i20_1_lut (.I0(setpoint[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[19]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i21_1_lut (.I0(setpoint[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[20]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i22_1_lut (.I0(setpoint[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[21]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694_adj_3980));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767_adj_3979));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840_adj_3978));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_3977));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_3976));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186_adj_3975));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259_adj_3974));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332_adj_3973));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 state_23__I_0_inv_0_i23_1_lut (.I0(setpoint[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[22]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 state_23__I_0_inv_0_i24_1_lut (.I0(setpoint[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4255[23]));   // verilog/motorControl.v(38[14:30])
    defparam state_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405_adj_3970));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478_adj_3969));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551_adj_3968));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624_adj_3967));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697_adj_3966));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770_adj_3965));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i17_3_lut (.I0(n155[16]), .I1(n1_adj_4253[16]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[16]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116_adj_3964));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47_adj_3963));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262_adj_3962));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_3961));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_3960));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_3959));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i18_3_lut (.I0(n155[17]), .I1(n1_adj_4253[17]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[17]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122_adj_3958));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_3957));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125_adj_3956));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_3955));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_983 (.I0(n6_adj_3937), .I1(\Ki[4] ), .I2(n8431[2]), 
            .I3(\PID_CONTROLLER.integral [18]), .O(n8424[3]));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut_adj_983.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i138_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23117_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [22]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n8442[0]));   // verilog/motorControl.v(42[26:37])
    defparam i23117_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 mult_11_i89_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i42_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_984 (.I0(n4_adj_3939), .I1(\Ki[3] ), .I2(n8437[1]), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n8431[2]));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut_adj_984.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(42[26:37])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_985 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral [23]), 
            .I3(\PID_CONTROLLER.integral [20]), .O(n12_adj_4247));   // verilog/motorControl.v(42[26:37])
    defparam i2_4_lut_adj_985.LUT_INIT = 16'h9c50;
    SB_LUT4 i23053_4_lut (.I0(n8431[2]), .I1(\Ki[4] ), .I2(n6_adj_3937), 
            .I3(\PID_CONTROLLER.integral [18]), .O(n8_adj_4248));   // verilog/motorControl.v(42[26:37])
    defparam i23053_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i1_4_lut_adj_986 (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n11_adj_4249));   // verilog/motorControl.v(42[26:37])
    defparam i1_4_lut_adj_986.LUT_INIT = 16'h6ca0;
    SB_LUT4 i23084_4_lut (.I0(n8437[1]), .I1(\Ki[3] ), .I2(n4_adj_3939), 
            .I3(\PID_CONTROLLER.integral [19]), .O(n6_adj_4250));   // verilog/motorControl.v(42[26:37])
    defparam i23084_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 i23119_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [22]), 
            .I3(\PID_CONTROLLER.integral [21]), .O(n27792));   // verilog/motorControl.v(42[26:37])
    defparam i23119_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut_adj_987 (.I0(n6_adj_4250), .I1(n11_adj_4249), .I2(n8_adj_4248), 
            .I3(n12_adj_4247), .O(n18_adj_4251));   // verilog/motorControl.v(42[26:37])
    defparam i8_4_lut_adj_987.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_988 (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(\PID_CONTROLLER.integral [22]), .O(n13_adj_4252));   // verilog/motorControl.v(42[26:37])
    defparam i3_4_lut_adj_988.LUT_INIT = 16'h6ca0;
    SB_LUT4 i9_4_lut_adj_989 (.I0(n13_adj_4252), .I1(n18_adj_4251), .I2(n27792), 
            .I3(n4_adj_3938), .O(n36379));   // verilog/motorControl.v(42[26:37])
    defparam i9_4_lut_adj_989.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i19_3_lut (.I0(n155[18]), .I1(n1_adj_4253[18]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[18]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[20]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_637_i20_3_lut (.I0(n155[19]), .I1(n1_adj_4253[19]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[19]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i21_3_lut (.I0(n155[20]), .I1(n1_adj_4253[20]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[20]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i22_3_lut (.I0(n155[21]), .I1(n1_adj_4253[21]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[21]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4254[21]));   // verilog/motorControl.v(39[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mux_637_i23_3_lut (.I0(n155[22]), .I1(n1_adj_4253[22]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[22]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_3940));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i23063_2_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(\Ki[1] ), .I3(\PID_CONTROLLER.integral [19]), .O(n8431[0]));   // verilog/motorControl.v(42[26:37])
    defparam i23063_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i24_3_lut (.I0(duty_23__N_3740[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[23]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i23_3_lut (.I0(duty_23__N_3740[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[22]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i22_3_lut (.I0(duty_23__N_3740[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[21]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i21_3_lut (.I0(duty_23__N_3740[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[20]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i20_3_lut (.I0(duty_23__N_3740[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[19]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i19_3_lut (.I0(duty_23__N_3740[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[18]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i18_3_lut (.I0(duty_23__N_3740[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[17]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i17_3_lut (.I0(duty_23__N_3740[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[16]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i16_3_lut (.I0(duty_23__N_3740[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[15]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i15_3_lut (.I0(duty_23__N_3740[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[14]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i14_3_lut (.I0(duty_23__N_3740[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[13]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i13_3_lut (.I0(duty_23__N_3740[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[12]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i12_3_lut (.I0(duty_23__N_3740[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[11]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i11_3_lut (.I0(duty_23__N_3740[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[10]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i10_3_lut (.I0(duty_23__N_3740[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[9]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i9_3_lut (.I0(duty_23__N_3740[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[8]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i8_3_lut (.I0(duty_23__N_3740[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[7]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i7_3_lut (.I0(duty_23__N_3740[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[6]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i6_3_lut (.I0(duty_23__N_3740[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[5]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i5_3_lut (.I0(duty_23__N_3740[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[4]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i4_3_lut (.I0(duty_23__N_3740[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[3]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_29_i3_3_lut (.I0(duty_23__N_3740[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[2]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(\PID_CONTROLLER.err [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_29_i2_3_lut (.I0(duty_23__N_3740[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3764), .I3(GND_net), .O(duty_23__N_3617[1]));   // verilog/motorControl.v(46[16] 48[10])
    defparam duty_23__I_0_29_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34109_2_lut_4_lut (.I0(duty[21]), .I1(n257[21]), .I2(duty[9]), 
            .I3(n257[9]), .O(n40955));
    defparam i34109_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i34170_2_lut_4_lut (.I0(duty[16]), .I1(n257[16]), .I2(duty[7]), 
            .I3(n257[7]), .O(n41016));
    defparam i34170_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mux_637_i24_3_lut_3_lut (.I0(PWMLimit[23]), .I1(n256_adj_3900), 
            .I2(n40677), .I3(GND_net), .O(n3073[23]));   // verilog/motorControl.v(47[19:28])
    defparam mux_637_i24_3_lut_3_lut.LUT_INIT = 16'h7474;
    SB_LUT4 duty_23__I_0_i8_3_lut_3_lut (.I0(duty[4]), .I1(duty[8]), .I2(PWMLimit[8]), 
            .I3(GND_net), .O(n8_adj_3893));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34273_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty[21]), .I2(PWMLimit[9]), 
            .I3(duty[9]), .O(n41120));
    defparam i34273_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i16_3_lut_3_lut (.I0(duty[9]), .I1(duty[21]), .I2(PWMLimit[21]), 
            .I3(GND_net), .O(n16_adj_3889));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i16_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(\PID_CONTROLLER.err [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_3921));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 duty_23__I_0_i10_3_lut_3_lut (.I0(duty[5]), .I1(duty[6]), .I2(PWMLimit[6]), 
            .I3(GND_net), .O(n10_adj_3896));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34298_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty[16]), .I2(PWMLimit[7]), 
            .I3(duty[7]), .O(n41145));
    defparam i34298_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_3882));   // verilog/motorControl.v(39[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 duty_23__I_0_i12_3_lut_3_lut (.I0(duty[7]), .I1(duty[16]), .I2(PWMLimit[16]), 
            .I3(GND_net), .O(n12_adj_3880));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(\PID_CONTROLLER.err [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(42[17:23])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i19555_2_lut_2_lut (.I0(n256_adj_3900), .I1(n6308[0]), .I2(GND_net), 
            .I3(GND_net), .O(n3048[23]));   // verilog/motorControl.v(46[19:35])
    defparam i19555_2_lut_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 mux_637_i3_3_lut (.I0(n155[2]), .I1(PWMLimit[2]), .I2(n256_adj_3900), 
            .I3(GND_net), .O(n3073[2]));   // verilog/motorControl.v(46[16] 48[10])
    defparam mux_637_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i34415_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty[3]), .I2(duty[2]), 
            .I3(PWMLimit[2]), .O(n41262));   // verilog/motorControl.v(44[10:25])
    defparam i34415_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_0_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty[3]), 
            .I2(duty[2]), .I3(GND_net), .O(n6_adj_3888));   // verilog/motorControl.v(44[10:25])
    defparam duty_23__I_0_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    
endmodule
//
// Verilog Description of module \quad(DEBOUNCE_TICKS=100)_U1 
//

module \quad(DEBOUNCE_TICKS=100)_U1  (n18176, encoder0_position, clk32MHz, 
            n18177, n18178, n18179, n18165, n18166, n18167, n18168, 
            n18169, n18170, n18171, n18172, n18173, n18174, n18175, 
            n18163, n18164, n18161, n18162, n18159, n18160, n18157, 
            n18158, data_o, GND_net, n2992, n17594, count_enable, 
            n18213, reg_B, n36518, PIN_2_c_0, PIN_1_c_1, n17597) /* synthesis lattice_noprune=1, syn_preserve=0, syn_module_defined=1, syn_noprune=0 */ ;
    input n18176;
    output [23:0]encoder0_position;
    input clk32MHz;
    input n18177;
    input n18178;
    input n18179;
    input n18165;
    input n18166;
    input n18167;
    input n18168;
    input n18169;
    input n18170;
    input n18171;
    input n18172;
    input n18173;
    input n18174;
    input n18175;
    input n18163;
    input n18164;
    input n18161;
    input n18162;
    input n18159;
    input n18160;
    input n18157;
    input n18158;
    output [1:0]data_o;
    input GND_net;
    output [23:0]n2992;
    input n17594;
    output count_enable;
    input n18213;
    output [1:0]reg_B;
    output n36518;
    input PIN_2_c_0;
    input PIN_1_c_1;
    input n17597;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    
    wire B_delayed, count_direction, A_delayed, n2988, n27999, n27998, 
        n27997, n27996, n27995, n27994, n27993, n27992, n27991, 
        n27990, n27989, n27988, n27987, n27986, n27985, n27984, 
        n27983, n27982, n27981, n27980, n27979, n27978, n27977, 
        n27976;
    
    SB_DFF count_i0_i20 (.Q(encoder0_position[20]), .C(clk32MHz), .D(n18176));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i21 (.Q(encoder0_position[21]), .C(clk32MHz), .D(n18177));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i22 (.Q(encoder0_position[22]), .C(clk32MHz), .D(n18178));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i23 (.Q(encoder0_position[23]), .C(clk32MHz), .D(n18179));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i9 (.Q(encoder0_position[9]), .C(clk32MHz), .D(n18165));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i10 (.Q(encoder0_position[10]), .C(clk32MHz), .D(n18166));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i11 (.Q(encoder0_position[11]), .C(clk32MHz), .D(n18167));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i12 (.Q(encoder0_position[12]), .C(clk32MHz), .D(n18168));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i13 (.Q(encoder0_position[13]), .C(clk32MHz), .D(n18169));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i14 (.Q(encoder0_position[14]), .C(clk32MHz), .D(n18170));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i15 (.Q(encoder0_position[15]), .C(clk32MHz), .D(n18171));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i16 (.Q(encoder0_position[16]), .C(clk32MHz), .D(n18172));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i17 (.Q(encoder0_position[17]), .C(clk32MHz), .D(n18173));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i18 (.Q(encoder0_position[18]), .C(clk32MHz), .D(n18174));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i19 (.Q(encoder0_position[19]), .C(clk32MHz), .D(n18175));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i7 (.Q(encoder0_position[7]), .C(clk32MHz), .D(n18163));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i8 (.Q(encoder0_position[8]), .C(clk32MHz), .D(n18164));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i5 (.Q(encoder0_position[5]), .C(clk32MHz), .D(n18161));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i6 (.Q(encoder0_position[6]), .C(clk32MHz), .D(n18162));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i3 (.Q(encoder0_position[3]), .C(clk32MHz), .D(n18159));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i4 (.Q(encoder0_position[4]), .C(clk32MHz), .D(n18160));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i1 (.Q(encoder0_position[1]), .C(clk32MHz), .D(n18157));   // quad.v(35[10] 41[6])
    SB_DFF count_i0_i2 (.Q(encoder0_position[2]), .C(clk32MHz), .D(n18158));   // quad.v(35[10] 41[6])
    SB_LUT4 quadA_debounced_I_0_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(count_direction));   // quad.v(26[26:53])
    defparam quadA_debounced_I_0_2_lut.LUT_INIT = 16'h6666;
    SB_DFF B_delayed_16 (.Q(B_delayed), .C(clk32MHz), .D(data_o[0]));   // quad.v(23[10:54])
    SB_DFF A_delayed_15 (.Q(A_delayed), .C(clk32MHz), .D(data_o[1]));   // quad.v(22[10:54])
    SB_LUT4 add_631_25_lut (.I0(GND_net), .I1(encoder0_position[23]), .I2(n2988), 
            .I3(n27999), .O(n2992[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_631_24_lut (.I0(GND_net), .I1(encoder0_position[22]), .I2(n2988), 
            .I3(n27998), .O(n2992[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_24 (.CI(n27998), .I0(encoder0_position[22]), .I1(n2988), 
            .CO(n27999));
    SB_LUT4 add_631_23_lut (.I0(GND_net), .I1(encoder0_position[21]), .I2(n2988), 
            .I3(n27997), .O(n2992[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_23 (.CI(n27997), .I0(encoder0_position[21]), .I1(n2988), 
            .CO(n27998));
    SB_LUT4 add_631_22_lut (.I0(GND_net), .I1(encoder0_position[20]), .I2(n2988), 
            .I3(n27996), .O(n2992[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_22 (.CI(n27996), .I0(encoder0_position[20]), .I1(n2988), 
            .CO(n27997));
    SB_LUT4 add_631_21_lut (.I0(GND_net), .I1(encoder0_position[19]), .I2(n2988), 
            .I3(n27995), .O(n2992[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_21 (.CI(n27995), .I0(encoder0_position[19]), .I1(n2988), 
            .CO(n27996));
    SB_LUT4 add_631_20_lut (.I0(GND_net), .I1(encoder0_position[18]), .I2(n2988), 
            .I3(n27994), .O(n2992[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_20 (.CI(n27994), .I0(encoder0_position[18]), .I1(n2988), 
            .CO(n27995));
    SB_LUT4 add_631_19_lut (.I0(GND_net), .I1(encoder0_position[17]), .I2(n2988), 
            .I3(n27993), .O(n2992[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_19 (.CI(n27993), .I0(encoder0_position[17]), .I1(n2988), 
            .CO(n27994));
    SB_LUT4 add_631_18_lut (.I0(GND_net), .I1(encoder0_position[16]), .I2(n2988), 
            .I3(n27992), .O(n2992[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_18 (.CI(n27992), .I0(encoder0_position[16]), .I1(n2988), 
            .CO(n27993));
    SB_LUT4 add_631_17_lut (.I0(GND_net), .I1(encoder0_position[15]), .I2(n2988), 
            .I3(n27991), .O(n2992[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_17 (.CI(n27991), .I0(encoder0_position[15]), .I1(n2988), 
            .CO(n27992));
    SB_LUT4 add_631_16_lut (.I0(GND_net), .I1(encoder0_position[14]), .I2(n2988), 
            .I3(n27990), .O(n2992[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_16 (.CI(n27990), .I0(encoder0_position[14]), .I1(n2988), 
            .CO(n27991));
    SB_LUT4 add_631_15_lut (.I0(GND_net), .I1(encoder0_position[13]), .I2(n2988), 
            .I3(n27989), .O(n2992[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_15 (.CI(n27989), .I0(encoder0_position[13]), .I1(n2988), 
            .CO(n27990));
    SB_LUT4 add_631_14_lut (.I0(GND_net), .I1(encoder0_position[12]), .I2(n2988), 
            .I3(n27988), .O(n2992[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_14 (.CI(n27988), .I0(encoder0_position[12]), .I1(n2988), 
            .CO(n27989));
    SB_LUT4 add_631_13_lut (.I0(GND_net), .I1(encoder0_position[11]), .I2(n2988), 
            .I3(n27987), .O(n2992[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_13 (.CI(n27987), .I0(encoder0_position[11]), .I1(n2988), 
            .CO(n27988));
    SB_LUT4 add_631_12_lut (.I0(GND_net), .I1(encoder0_position[10]), .I2(n2988), 
            .I3(n27986), .O(n2992[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_12 (.CI(n27986), .I0(encoder0_position[10]), .I1(n2988), 
            .CO(n27987));
    SB_LUT4 add_631_11_lut (.I0(GND_net), .I1(encoder0_position[9]), .I2(n2988), 
            .I3(n27985), .O(n2992[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_11 (.CI(n27985), .I0(encoder0_position[9]), .I1(n2988), 
            .CO(n27986));
    SB_LUT4 add_631_10_lut (.I0(GND_net), .I1(encoder0_position[8]), .I2(n2988), 
            .I3(n27984), .O(n2992[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_10 (.CI(n27984), .I0(encoder0_position[8]), .I1(n2988), 
            .CO(n27985));
    SB_LUT4 add_631_9_lut (.I0(GND_net), .I1(encoder0_position[7]), .I2(n2988), 
            .I3(n27983), .O(n2992[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_9 (.CI(n27983), .I0(encoder0_position[7]), .I1(n2988), 
            .CO(n27984));
    SB_LUT4 add_631_8_lut (.I0(GND_net), .I1(encoder0_position[6]), .I2(n2988), 
            .I3(n27982), .O(n2992[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_8 (.CI(n27982), .I0(encoder0_position[6]), .I1(n2988), 
            .CO(n27983));
    SB_LUT4 add_631_7_lut (.I0(GND_net), .I1(encoder0_position[5]), .I2(n2988), 
            .I3(n27981), .O(n2992[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_7 (.CI(n27981), .I0(encoder0_position[5]), .I1(n2988), 
            .CO(n27982));
    SB_DFF count_i0_i0 (.Q(encoder0_position[0]), .C(clk32MHz), .D(n17594));   // quad.v(35[10] 41[6])
    SB_LUT4 add_631_6_lut (.I0(GND_net), .I1(encoder0_position[4]), .I2(n2988), 
            .I3(n27980), .O(n2992[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_6 (.CI(n27980), .I0(encoder0_position[4]), .I1(n2988), 
            .CO(n27981));
    SB_LUT4 add_631_5_lut (.I0(GND_net), .I1(encoder0_position[3]), .I2(n2988), 
            .I3(n27979), .O(n2992[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_5 (.CI(n27979), .I0(encoder0_position[3]), .I1(n2988), 
            .CO(n27980));
    SB_LUT4 add_631_4_lut (.I0(GND_net), .I1(encoder0_position[2]), .I2(n2988), 
            .I3(n27978), .O(n2992[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_4 (.CI(n27978), .I0(encoder0_position[2]), .I1(n2988), 
            .CO(n27979));
    SB_LUT4 add_631_3_lut (.I0(GND_net), .I1(encoder0_position[1]), .I2(n2988), 
            .I3(n27977), .O(n2992[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_3 (.CI(n27977), .I0(encoder0_position[1]), .I1(n2988), 
            .CO(n27978));
    SB_LUT4 add_631_2_lut (.I0(GND_net), .I1(encoder0_position[0]), .I2(count_direction), 
            .I3(n27976), .O(n2992[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_631_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_631_2 (.CI(n27976), .I0(encoder0_position[0]), .I1(count_direction), 
            .CO(n27977));
    SB_CARRY add_631_1 (.CI(GND_net), .I0(n2988), .I1(n2988), .CO(n27976));
    SB_LUT4 i3_4_lut (.I0(data_o[1]), .I1(A_delayed), .I2(B_delayed), 
            .I3(data_o[0]), .O(count_enable));   // quad.v(25[23:80])
    defparam i3_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i937_1_lut_2_lut (.I0(data_o[1]), .I1(B_delayed), .I2(GND_net), 
            .I3(GND_net), .O(n2988));   // quad.v(37[5] 40[8])
    defparam i937_1_lut_2_lut.LUT_INIT = 16'h9999;
    \grp_debouncer(2,5)_U0  debounce (.n18213(n18213), .data_o({data_o}), 
            .clk32MHz(clk32MHz), .reg_B({reg_B}), .GND_net(GND_net), .n36518(n36518), 
            .PIN_2_c_0(PIN_2_c_0), .PIN_1_c_1(PIN_1_c_1), .n17597(n17597)) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;   // quad.v(15[24] 19[4])
    
endmodule
//
// Verilog Description of module \grp_debouncer(2,5)_U0 
//

module \grp_debouncer(2,5)_U0  (n18213, data_o, clk32MHz, reg_B, GND_net, 
            n36518, PIN_2_c_0, PIN_1_c_1, n17597) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input n18213;
    output [1:0]data_o;
    input clk32MHz;
    output [1:0]reg_B;
    input GND_net;
    output n36518;
    input PIN_2_c_0;
    input PIN_1_c_1;
    input n17597;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(34[6:14])
    wire [1:0]reg_A;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(142[12:17])
    
    wire n2, cnt_next_2__N_3821;
    wire [2:0]cnt_reg;   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(149[12:19])
    wire [2:0]n17;
    
    SB_DFF reg_out_i0_i1 (.Q(data_o[1]), .C(clk32MHz), .D(n18213));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_LUT4 reg_B_1__I_0_i2_2_lut (.I0(reg_B[1]), .I1(reg_A[1]), .I2(GND_net), 
            .I3(GND_net), .O(n2));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(193[46:60])
    defparam reg_B_1__I_0_i2_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_4_lut (.I0(reg_B[0]), .I1(n36518), .I2(reg_A[0]), .I3(n2), 
            .O(cnt_next_2__N_3821));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[40:72])
    defparam i2_4_lut.LUT_INIT = 16'hff7b;
    SB_LUT4 i22812_1_lut (.I0(cnt_reg[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22812_1_lut.LUT_INIT = 16'h5555;
    SB_DFF reg_B_i0 (.Q(reg_B[0]), .C(clk32MHz), .D(reg_A[0]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFFSR cnt_reg_1226__i0 (.Q(cnt_reg[0]), .C(clk32MHz), .D(n17[0]), 
            .R(cnt_next_2__N_3821));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i2_3_lut (.I0(cnt_reg[0]), .I1(cnt_reg[2]), .I2(cnt_reg[1]), 
            .I3(GND_net), .O(n36518));
    defparam i2_3_lut.LUT_INIT = 16'hf7f7;
    SB_DFF reg_B_i1 (.Q(reg_B[1]), .C(clk32MHz), .D(reg_A[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i0 (.Q(reg_A[0]), .C(clk32MHz), .D(PIN_2_c_0));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_A_i1 (.Q(reg_A[1]), .C(clk32MHz), .D(PIN_1_c_1));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(178[9] 184[16])
    SB_DFF reg_out_i0_i0 (.Q(data_o[0]), .C(clk32MHz), .D(n17597));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(186[9] 190[16])
    SB_DFFSR cnt_reg_1226__i1 (.Q(cnt_reg[1]), .C(clk32MHz), .D(n17[1]), 
            .R(cnt_next_2__N_3821));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_DFFSR cnt_reg_1226__i2 (.Q(cnt_reg[2]), .C(clk32MHz), .D(n17[2]), 
            .R(cnt_next_2__N_3821));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    SB_LUT4 i22821_3_lut (.I0(cnt_reg[2]), .I1(cnt_reg[1]), .I2(cnt_reg[0]), 
            .I3(GND_net), .O(n17[2]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22821_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i22814_2_lut (.I0(cnt_reg[1]), .I1(cnt_reg[0]), .I2(GND_net), 
            .I3(GND_net), .O(n17[1]));   // vhdl/spi_master_slave/trunk/rtl/spi_master_slave/grp_debouncer.vhd(168[78:85])
    defparam i22814_2_lut.LUT_INIT = 16'h6666;
    
endmodule
//
// Verilog Description of module \pwm(32000000,20000,32000000,23,1) 
//

module \pwm(32000000,20000,32000000,23,1)  (GND_net, VCC_net, \half_duty_new[0] , 
            CLK_c, PIN_19_c_0, pwm_setpoint, n18253, \half_duty[0][1] , 
            n18254, \half_duty[0][2] , n18255, \half_duty[0][3] , n18256, 
            \half_duty[0][4] , n18258, \half_duty[0][6] , n18259, \half_duty[0][7] , 
            \half_duty[0][0] , n1170, \half_duty_new[1] , \half_duty_new[2] , 
            \half_duty_new[3] , \half_duty_new[4] , \half_duty_new[6] , 
            \half_duty_new[7] , n17617) /* synthesis lattice_noprune=1, syn_preserve=0, syn_noprune=0 */ ;
    input GND_net;
    input VCC_net;
    output \half_duty_new[0] ;
    input CLK_c;
    output PIN_19_c_0;
    input [22:0]pwm_setpoint;
    input n18253;
    output \half_duty[0][1] ;
    input n18254;
    output \half_duty[0][2] ;
    input n18255;
    output \half_duty[0][3] ;
    input n18256;
    output \half_duty[0][4] ;
    input n18258;
    output \half_duty[0][6] ;
    input n18259;
    output \half_duty[0][7] ;
    output \half_duty[0][0] ;
    output n1170;
    output \half_duty_new[1] ;
    output \half_duty_new[2] ;
    output \half_duty_new[3] ;
    output \half_duty_new[4] ;
    output \half_duty_new[6] ;
    output \half_duty_new[7] ;
    input n17617;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n42887, n27879;
    wire [10:0]\count[0] ;   // vhdl/pwm.vhd(51[11:16])
    
    wire n27882, pwm_out_0__N_586, n27880;
    wire [9:0]half_duty_new_9__N_664;
    
    wire n8;
    wire [10:0]pwm_out_0__N_587;
    
    wire n27878, pwm_out_0__N_582, n17199, n27881, n42891, n27877;
    wire [22:0]n5649;
    
    wire n27836, n42885, n27876, n27837, n22753;
    wire [9:0]\half_duty[0] ;   // vhdl/pwm.vhd(55[11:20])
    wire [10:0]n49;
    
    wire pause_counter_0__N_612, n27835, pause_counter_0, n35811, n27824, 
        n5, n27875, n4, n27874, n27825, n27834, n3, n27873, 
        n2, n27872, n28611, n28610, n28609, n28608, n28607, n28606, 
        n28605, n28604, n28603, n28602, n27823, n27833, n1, n27832, 
        n27822, n27831, n20, n13, n22, n10, n38571, n13_adj_3823, 
        n3_adj_3824, n18, n16, n17, n15;
    wire [9:0]half_duty_new;   // vhdl/pwm.vhd(53[12:25])
    
    wire n27830, n27821, n27829, n28267, n28266, n28265, n28264, 
        n28263, n28262, n28261, n28260, n28259, n28258, n28257, 
        n28256, n28255, n28254, n28253, n28252, n28251, n28250, 
        n28249, n28248, n28247, n28246, n27820, n27828, n27827, 
        n27826, n27840, n27839, n27838, n38553, n12, n18_adj_3825, 
        n19;
    
    SB_LUT4 pwm_out_0__I_20_10_lut (.I0(\count[0] [8]), .I1(GND_net), .I2(VCC_net), 
            .I3(n27879), .O(n42887)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_10_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_13 (.CI(n27882), .I0(GND_net), .I1(VCC_net), 
            .CO(pwm_out_0__N_586));
    SB_CARRY pwm_out_0__I_20_10 (.CI(n27879), .I0(GND_net), .I1(VCC_net), 
            .CO(n27880));
    SB_DFF half_duty_new_i1 (.Q(\half_duty_new[0] ), .C(CLK_c), .D(half_duty_new_9__N_664[0]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 pwm_out_0__I_20_9_lut (.I0(\count[0] [7]), .I1(GND_net), .I2(pwm_out_0__N_587[7]), 
            .I3(n27878), .O(n8)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_9_lut.LUT_INIT = 16'h6996;
    SB_DFFE pwm_out_0__39 (.Q(PIN_19_c_0), .C(CLK_c), .E(n17199), .D(pwm_out_0__N_582));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_CARRY pwm_out_0__I_20_12 (.CI(n27881), .I0(VCC_net), .I1(VCC_net), 
            .CO(n27882));
    SB_CARRY pwm_out_0__I_20_9 (.CI(n27878), .I0(GND_net), .I1(pwm_out_0__N_587[7]), 
            .CO(n27879));
    SB_LUT4 pwm_out_0__I_20_8_lut (.I0(\count[0] [6]), .I1(VCC_net), .I2(pwm_out_0__N_587[6]), 
            .I3(n27877), .O(n42891)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_8_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_2096_19_lut (.I0(GND_net), .I1(pwm_setpoint[17]), .I2(pwm_setpoint[21]), 
            .I3(n27836), .O(n5649[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_out_0__I_20_8 (.CI(n27877), .I0(VCC_net), .I1(pwm_out_0__N_587[6]), 
            .CO(n27878));
    SB_LUT4 pwm_out_0__I_20_7_lut (.I0(\count[0] [5]), .I1(GND_net), .I2(pwm_out_0__N_587[5]), 
            .I3(n27876), .O(n42885)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_7_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_2096_19 (.CI(n27836), .I0(pwm_setpoint[17]), .I1(pwm_setpoint[21]), 
            .CO(n27837));
    SB_DFF half_duty_0___i2 (.Q(\half_duty[0][1] ), .C(CLK_c), .D(n18253));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i3 (.Q(\half_duty[0][2] ), .C(CLK_c), .D(n18254));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i4 (.Q(\half_duty[0][3] ), .C(CLK_c), .D(n18255));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i5 (.Q(\half_duty[0][4] ), .C(CLK_c), .D(n18256));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i6 (.Q(\half_duty[0] [5]), .C(CLK_c), .D(n22753));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i7 (.Q(\half_duty[0][6] ), .C(CLK_c), .D(n18258));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_0___i8 (.Q(\half_duty[0][7] ), .C(CLK_c), .D(n18259));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 half_duty_0__9__I_0_i1_1_lut (.I0(\half_duty[0][0] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[0]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY pwm_out_0__I_20_7 (.CI(n27876), .I0(GND_net), .I1(pwm_out_0__N_587[5]), 
            .CO(n27877));
    SB_DFFESR count_0__1224__i10 (.Q(\count[0] [10]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[10]), .R(n1170));   // vhdl/pwm.vhd(77[18:26])
    SB_LUT4 add_2096_18_lut (.I0(GND_net), .I1(pwm_setpoint[16]), .I2(pwm_setpoint[20]), 
            .I3(n27835), .O(n5649[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_18_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR count_0__1224__i9 (.Q(\count[0] [9]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[9]), .R(n1170));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1224__i8 (.Q(\count[0] [8]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[8]), .R(n1170));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1224__i7 (.Q(\count[0] [7]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[7]), .R(n1170));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1224__i6 (.Q(\count[0] [6]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[6]), .R(n1170));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1224__i5 (.Q(\count[0] [5]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[5]), .R(n1170));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1224__i4 (.Q(\count[0] [4]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[4]), .R(n1170));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1224__i3 (.Q(\count[0] [3]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[3]), .R(n1170));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1224__i2 (.Q(\count[0] [2]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[2]), .R(n1170));   // vhdl/pwm.vhd(77[18:26])
    SB_DFFESR count_0__1224__i1 (.Q(\count[0] [1]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[1]), .R(n1170));   // vhdl/pwm.vhd(77[18:26])
    SB_LUT4 i36782_2_lut (.I0(pause_counter_0), .I1(pwm_out_0__N_582), .I2(GND_net), 
            .I3(GND_net), .O(n35811));
    defparam i36782_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 add_2096_7_lut (.I0(GND_net), .I1(pwm_setpoint[5]), .I2(pwm_setpoint[9]), 
            .I3(n27824), .O(n5649[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_out_0__I_20_11 (.CI(n27880), .I0(VCC_net), .I1(VCC_net), 
            .CO(n27881));
    SB_LUT4 pwm_out_0__I_20_6_lut (.I0(\count[0] [4]), .I1(GND_net), .I2(pwm_out_0__N_587[4]), 
            .I3(n27875), .O(n5)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_6 (.CI(n27875), .I0(GND_net), .I1(pwm_out_0__N_587[4]), 
            .CO(n27876));
    SB_CARRY add_2096_18 (.CI(n27835), .I0(pwm_setpoint[16]), .I1(pwm_setpoint[20]), 
            .CO(n27836));
    SB_LUT4 pwm_out_0__I_20_5_lut (.I0(\count[0] [3]), .I1(GND_net), .I2(pwm_out_0__N_587[3]), 
            .I3(n27874), .O(n4)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_5_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_5 (.CI(n27874), .I0(GND_net), .I1(pwm_out_0__N_587[3]), 
            .CO(n27875));
    SB_CARRY add_2096_7 (.CI(n27824), .I0(pwm_setpoint[5]), .I1(pwm_setpoint[9]), 
            .CO(n27825));
    SB_LUT4 add_2096_17_lut (.I0(GND_net), .I1(pwm_setpoint[15]), .I2(pwm_setpoint[19]), 
            .I3(n27834), .O(n5649[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2096_17 (.CI(n27834), .I0(pwm_setpoint[15]), .I1(pwm_setpoint[19]), 
            .CO(n27835));
    SB_LUT4 pwm_out_0__I_20_4_lut (.I0(\count[0] [2]), .I1(GND_net), .I2(pwm_out_0__N_587[2]), 
            .I3(n27873), .O(n3)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY pwm_out_0__I_20_4 (.CI(n27873), .I0(GND_net), .I1(pwm_out_0__N_587[2]), 
            .CO(n27874));
    SB_LUT4 pwm_out_0__I_20_3_lut (.I0(\count[0] [1]), .I1(GND_net), .I2(pwm_out_0__N_587[1]), 
            .I3(n27872), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 count_0__1224_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [10]), 
            .I3(n28611), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1224_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 count_0__1224_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [9]), 
            .I3(n28610), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1224_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1224_add_4_11 (.CI(n28610), .I0(GND_net), .I1(\count[0] [9]), 
            .CO(n28611));
    SB_LUT4 count_0__1224_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [8]), 
            .I3(n28609), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1224_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1224_add_4_10 (.CI(n28609), .I0(GND_net), .I1(\count[0] [8]), 
            .CO(n28610));
    SB_LUT4 count_0__1224_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [7]), 
            .I3(n28608), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1224_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1224_add_4_9 (.CI(n28608), .I0(GND_net), .I1(\count[0] [7]), 
            .CO(n28609));
    SB_LUT4 count_0__1224_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [6]), 
            .I3(n28607), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1224_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1224_add_4_8 (.CI(n28607), .I0(GND_net), .I1(\count[0] [6]), 
            .CO(n28608));
    SB_LUT4 count_0__1224_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [5]), 
            .I3(n28606), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1224_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1224_add_4_7 (.CI(n28606), .I0(GND_net), .I1(\count[0] [5]), 
            .CO(n28607));
    SB_LUT4 count_0__1224_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [4]), 
            .I3(n28605), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1224_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1224_add_4_6 (.CI(n28605), .I0(GND_net), .I1(\count[0] [4]), 
            .CO(n28606));
    SB_LUT4 count_0__1224_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [3]), 
            .I3(n28604), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1224_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1224_add_4_5 (.CI(n28604), .I0(GND_net), .I1(\count[0] [3]), 
            .CO(n28605));
    SB_LUT4 count_0__1224_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [2]), 
            .I3(n28603), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1224_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1224_add_4_4 (.CI(n28603), .I0(GND_net), .I1(\count[0] [2]), 
            .CO(n28604));
    SB_LUT4 count_0__1224_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [1]), 
            .I3(n28602), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1224_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1224_add_4_3 (.CI(n28602), .I0(GND_net), .I1(\count[0] [1]), 
            .CO(n28603));
    SB_LUT4 count_0__1224_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(\count[0] [0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam count_0__1224_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY count_0__1224_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(\count[0] [0]), 
            .CO(n28602));
    SB_LUT4 add_2096_6_lut (.I0(GND_net), .I1(pwm_setpoint[4]), .I2(pwm_setpoint[8]), 
            .I3(n27823), .O(n5649[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2096_16_lut (.I0(GND_net), .I1(pwm_setpoint[14]), .I2(pwm_setpoint[18]), 
            .I3(n27833), .O(n5649[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_16_lut.LUT_INIT = 16'hC33C;
    SB_DFF pause_counter_0__38 (.Q(pause_counter_0), .C(CLK_c), .D(n35811));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_CARRY pwm_out_0__I_20_3 (.CI(n27872), .I0(GND_net), .I1(pwm_out_0__N_587[1]), 
            .CO(n27873));
    SB_LUT4 half_duty_0__9__I_0_i2_1_lut (.I0(\half_duty[0][1] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[1]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 pwm_out_0__I_20_2_lut (.I0(\count[0] [0]), .I1(GND_net), .I2(pwm_out_0__N_587[0]), 
            .I3(VCC_net), .O(n1)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_2_lut.LUT_INIT = 16'h6996;
    SB_LUT4 half_duty_0__9__I_0_i3_1_lut (.I0(\half_duty[0][2] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[2]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY pwm_out_0__I_20_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_out_0__N_587[0]), 
            .CO(n27872));
    SB_CARRY add_2096_6 (.CI(n27823), .I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .CO(n27824));
    SB_CARRY add_2096_16 (.CI(n27833), .I0(pwm_setpoint[14]), .I1(pwm_setpoint[18]), 
            .CO(n27834));
    SB_LUT4 add_2096_15_lut (.I0(GND_net), .I1(pwm_setpoint[13]), .I2(pwm_setpoint[17]), 
            .I3(n27832), .O(n5649[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_15_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR count_0__1224__i0 (.Q(\count[0] [0]), .C(CLK_c), .E(pause_counter_0__N_612), 
            .D(n49[0]), .R(n1170));   // vhdl/pwm.vhd(77[18:26])
    SB_LUT4 add_2096_5_lut (.I0(GND_net), .I1(pwm_setpoint[3]), .I2(pwm_setpoint[7]), 
            .I3(n27822), .O(n5649[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 half_duty_0__9__I_0_i4_1_lut (.I0(\half_duty[0][3] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[3]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 half_duty_0__9__I_0_i5_1_lut (.I0(\half_duty[0][4] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[4]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2096_15 (.CI(n27832), .I0(pwm_setpoint[13]), .I1(pwm_setpoint[17]), 
            .CO(n27833));
    SB_LUT4 pause_counter_0__I_0_48_1_lut (.I0(pause_counter_0), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pause_counter_0__N_612));   // vhdl/pwm.vhd(72[7:27])
    defparam pause_counter_0__I_0_48_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_2096_14_lut (.I0(GND_net), .I1(pwm_setpoint[12]), .I2(pwm_setpoint[16]), 
            .I3(n27831), .O(n5649[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2096_5 (.CI(n27822), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[7]), 
            .CO(n27823));
    SB_LUT4 half_duty_0__9__I_0_i6_1_lut (.I0(\half_duty[0] [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[5]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_2096_14 (.CI(n27831), .I0(pwm_setpoint[12]), .I1(pwm_setpoint[16]), 
            .CO(n27832));
    SB_LUT4 i18035_1_lut (.I0(\half_duty[0][6] ), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(pwm_out_0__N_587[6]));   // vhdl/pwm.vhd(59[5] 95[12])
    defparam i18035_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i8_4_lut (.I0(n4), .I1(n42887), .I2(n42891), .I3(pwm_out_0__N_586), 
            .O(n20));
    defparam i8_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i1_2_lut (.I0(\count[0] [10]), .I1(n5), .I2(GND_net), .I3(GND_net), 
            .O(n13));
    defparam i1_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i10_4_lut (.I0(n13), .I1(n20), .I2(n8), .I3(n42885), .O(n22));
    defparam i10_4_lut.LUT_INIT = 16'h0008;
    SB_LUT4 i31799_4_lut (.I0(n2), .I1(n3), .I2(n10), .I3(n1), .O(n38571));
    defparam i31799_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut (.I0(n38571), .I1(pause_counter_0), .I2(pwm_out_0__N_582), 
            .I3(n22), .O(n17199));
    defparam i1_4_lut.LUT_INIT = 16'h1303;
    SB_LUT4 i2_4_lut (.I0(\count[0] [6]), .I1(\count[0] [5]), .I2(\half_duty[0][6] ), 
            .I3(\half_duty[0] [5]), .O(n13_adj_3823));   // vhdl/pwm.vhd(80[8:31])
    defparam i2_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 half_duty_0__9__I_0_47_i3_2_lut (.I0(\half_duty[0][2] ), .I1(\count[0] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_3824));   // vhdl/pwm.vhd(80[8:31])
    defparam half_duty_0__9__I_0_47_i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut (.I0(n13_adj_3823), .I1(\half_duty[0][7] ), .I2(\count[0] [9]), 
            .I3(\count[0] [7]), .O(n18));   // vhdl/pwm.vhd(80[8:31])
    defparam i7_4_lut.LUT_INIT = 16'hfbfe;
    SB_LUT4 i5_3_lut (.I0(\count[0] [8]), .I1(\count[0] [0]), .I2(\half_duty[0][0] ), 
            .I3(GND_net), .O(n16));   // vhdl/pwm.vhd(80[8:31])
    defparam i5_3_lut.LUT_INIT = 16'hbebe;
    SB_LUT4 i6_4_lut (.I0(\half_duty[0][3] ), .I1(n3_adj_3824), .I2(\count[0] [3]), 
            .I3(\count[0] [10]), .O(n17));   // vhdl/pwm.vhd(80[8:31])
    defparam i6_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i4_4_lut (.I0(\half_duty[0][4] ), .I1(\half_duty[0][1] ), .I2(\count[0] [4]), 
            .I3(\count[0] [1]), .O(n15));   // vhdl/pwm.vhd(80[8:31])
    defparam i4_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i10_4_lut_adj_969 (.I0(n15), .I1(n17), .I2(n16), .I3(n18), 
            .O(pwm_out_0__N_582));   // vhdl/pwm.vhd(80[8:31])
    defparam i10_4_lut_adj_969.LUT_INIT = 16'hfffe;
    SB_LUT4 half_duty_0__9__I_0_i8_1_lut (.I0(\half_duty[0][7] ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(pwm_out_0__N_587[7]));   // vhdl/pwm.vhd(84[22:28])
    defparam half_duty_0__9__I_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_DFF half_duty_new_i2 (.Q(\half_duty_new[1] ), .C(CLK_c), .D(half_duty_new_9__N_664[1]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i3 (.Q(\half_duty_new[2] ), .C(CLK_c), .D(half_duty_new_9__N_664[2]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i4 (.Q(\half_duty_new[3] ), .C(CLK_c), .D(half_duty_new_9__N_664[3]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i5 (.Q(\half_duty_new[4] ), .C(CLK_c), .D(half_duty_new_9__N_664[4]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i6 (.Q(half_duty_new[5]), .C(CLK_c), .D(half_duty_new_9__N_664[5]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i7 (.Q(\half_duty_new[6] ), .C(CLK_c), .D(half_duty_new_9__N_664[6]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_DFF half_duty_new_i8 (.Q(\half_duty_new[7] ), .C(CLK_c), .D(half_duty_new_9__N_664[7]));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_LUT4 add_2096_13_lut (.I0(GND_net), .I1(pwm_setpoint[11]), .I2(pwm_setpoint[15]), 
            .I3(n27830), .O(n5649[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2096_4_lut (.I0(GND_net), .I1(pwm_setpoint[2]), .I2(pwm_setpoint[6]), 
            .I3(n27821), .O(n5649[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2096_13 (.CI(n27830), .I0(pwm_setpoint[11]), .I1(pwm_setpoint[15]), 
            .CO(n27831));
    SB_LUT4 add_2096_12_lut (.I0(GND_net), .I1(pwm_setpoint[10]), .I2(pwm_setpoint[14]), 
            .I3(n27829), .O(n5649[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF half_duty_0___i1 (.Q(\half_duty[0][0] ), .C(CLK_c), .D(n17617));   // vhdl/pwm.vhd(59[5] 95[12])
    SB_CARRY add_2096_4 (.CI(n27821), .I0(pwm_setpoint[2]), .I1(pwm_setpoint[6]), 
            .CO(n27822));
    SB_LUT4 add_2086_24_lut (.I0(GND_net), .I1(n5649[22]), .I2(pwm_setpoint[22]), 
            .I3(n28267), .O(half_duty_new_9__N_664[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2086_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2086_23_lut (.I0(GND_net), .I1(n5649[21]), .I2(pwm_setpoint[21]), 
            .I3(n28266), .O(half_duty_new_9__N_664[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2086_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2086_23 (.CI(n28266), .I0(n5649[21]), .I1(pwm_setpoint[21]), 
            .CO(n28267));
    SB_LUT4 add_2086_22_lut (.I0(GND_net), .I1(n5649[20]), .I2(pwm_setpoint[20]), 
            .I3(n28265), .O(half_duty_new_9__N_664[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2086_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2086_22 (.CI(n28265), .I0(n5649[20]), .I1(pwm_setpoint[20]), 
            .CO(n28266));
    SB_LUT4 add_2086_21_lut (.I0(GND_net), .I1(n5649[19]), .I2(pwm_setpoint[19]), 
            .I3(n28264), .O(half_duty_new_9__N_664[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2086_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2086_21 (.CI(n28264), .I0(n5649[19]), .I1(pwm_setpoint[19]), 
            .CO(n28265));
    SB_LUT4 add_2086_20_lut (.I0(GND_net), .I1(n5649[18]), .I2(pwm_setpoint[18]), 
            .I3(n28263), .O(half_duty_new_9__N_664[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2086_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2086_20 (.CI(n28263), .I0(n5649[18]), .I1(pwm_setpoint[18]), 
            .CO(n28264));
    SB_LUT4 add_2086_19_lut (.I0(GND_net), .I1(n5649[17]), .I2(pwm_setpoint[17]), 
            .I3(n28262), .O(half_duty_new_9__N_664[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2086_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2086_19 (.CI(n28262), .I0(n5649[17]), .I1(pwm_setpoint[17]), 
            .CO(n28263));
    SB_LUT4 add_2086_18_lut (.I0(GND_net), .I1(n5649[16]), .I2(pwm_setpoint[16]), 
            .I3(n28261), .O(half_duty_new_9__N_664[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2086_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2086_18 (.CI(n28261), .I0(n5649[16]), .I1(pwm_setpoint[16]), 
            .CO(n28262));
    SB_LUT4 add_2086_17_lut (.I0(GND_net), .I1(n5649[15]), .I2(pwm_setpoint[15]), 
            .I3(n28260), .O(half_duty_new_9__N_664[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2086_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2086_17 (.CI(n28260), .I0(n5649[15]), .I1(pwm_setpoint[15]), 
            .CO(n28261));
    SB_CARRY add_2086_16 (.CI(n28259), .I0(n5649[14]), .I1(pwm_setpoint[14]), 
            .CO(n28260));
    SB_CARRY add_2086_15 (.CI(n28258), .I0(n5649[13]), .I1(pwm_setpoint[13]), 
            .CO(n28259));
    SB_CARRY add_2086_14 (.CI(n28257), .I0(n5649[12]), .I1(pwm_setpoint[12]), 
            .CO(n28258));
    SB_CARRY add_2086_13 (.CI(n28256), .I0(n5649[11]), .I1(pwm_setpoint[11]), 
            .CO(n28257));
    SB_CARRY add_2086_12 (.CI(n28255), .I0(n5649[10]), .I1(pwm_setpoint[10]), 
            .CO(n28256));
    SB_CARRY add_2086_11 (.CI(n28254), .I0(n5649[9]), .I1(pwm_setpoint[9]), 
            .CO(n28255));
    SB_CARRY add_2086_10 (.CI(n28253), .I0(n5649[8]), .I1(pwm_setpoint[8]), 
            .CO(n28254));
    SB_CARRY add_2086_9 (.CI(n28252), .I0(n5649[7]), .I1(pwm_setpoint[7]), 
            .CO(n28253));
    SB_CARRY add_2086_8 (.CI(n28251), .I0(n5649[6]), .I1(pwm_setpoint[6]), 
            .CO(n28252));
    SB_CARRY add_2086_7 (.CI(n28250), .I0(n5649[5]), .I1(pwm_setpoint[5]), 
            .CO(n28251));
    SB_CARRY add_2086_6 (.CI(n28249), .I0(n5649[4]), .I1(pwm_setpoint[4]), 
            .CO(n28250));
    SB_CARRY add_2086_5 (.CI(n28248), .I0(n5649[3]), .I1(pwm_setpoint[3]), 
            .CO(n28249));
    SB_CARRY add_2086_4 (.CI(n28247), .I0(n5649[2]), .I1(pwm_setpoint[2]), 
            .CO(n28248));
    SB_CARRY add_2086_3 (.CI(n28246), .I0(n5649[1]), .I1(pwm_setpoint[1]), 
            .CO(n28247));
    SB_CARRY add_2086_2 (.CI(GND_net), .I0(pwm_setpoint[3]), .I1(pwm_setpoint[0]), 
            .CO(n28246));
    SB_CARRY add_2096_12 (.CI(n27829), .I0(pwm_setpoint[10]), .I1(pwm_setpoint[14]), 
            .CO(n27830));
    SB_LUT4 add_2096_3_lut (.I0(GND_net), .I1(pwm_setpoint[1]), .I2(pwm_setpoint[5]), 
            .I3(n27820), .O(n5649[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2096_11_lut (.I0(GND_net), .I1(pwm_setpoint[9]), .I2(pwm_setpoint[13]), 
            .I3(n27828), .O(n5649[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2096_11 (.CI(n27828), .I0(pwm_setpoint[9]), .I1(pwm_setpoint[13]), 
            .CO(n27829));
    SB_LUT4 add_2096_10_lut (.I0(GND_net), .I1(pwm_setpoint[8]), .I2(pwm_setpoint[12]), 
            .I3(n27827), .O(n5649[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2096_3 (.CI(n27820), .I0(pwm_setpoint[1]), .I1(pwm_setpoint[5]), 
            .CO(n27821));
    SB_LUT4 add_2096_2_lut (.I0(GND_net), .I1(pwm_setpoint[0]), .I2(pwm_setpoint[4]), 
            .I3(GND_net), .O(n5649[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2096_10 (.CI(n27827), .I0(pwm_setpoint[8]), .I1(pwm_setpoint[12]), 
            .CO(n27828));
    SB_LUT4 add_2096_9_lut (.I0(GND_net), .I1(pwm_setpoint[7]), .I2(pwm_setpoint[11]), 
            .I3(n27826), .O(n5649[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2096_9 (.CI(n27826), .I0(pwm_setpoint[7]), .I1(pwm_setpoint[11]), 
            .CO(n27827));
    SB_LUT4 add_2096_8_lut (.I0(GND_net), .I1(pwm_setpoint[6]), .I2(pwm_setpoint[10]), 
            .I3(n27825), .O(n5649[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2096_2 (.CI(GND_net), .I0(pwm_setpoint[0]), .I1(pwm_setpoint[4]), 
            .CO(n27820));
    SB_CARRY add_2096_8 (.CI(n27825), .I0(pwm_setpoint[6]), .I1(pwm_setpoint[10]), 
            .CO(n27826));
    SB_LUT4 add_2096_23_lut (.I0(GND_net), .I1(pwm_setpoint[21]), .I2(GND_net), 
            .I3(n27840), .O(n5649[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_2096_22_lut (.I0(GND_net), .I1(pwm_setpoint[20]), .I2(GND_net), 
            .I3(n27839), .O(n5649[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2096_22 (.CI(n27839), .I0(pwm_setpoint[20]), .I1(GND_net), 
            .CO(n27840));
    SB_LUT4 add_2096_21_lut (.I0(GND_net), .I1(pwm_setpoint[19]), .I2(GND_net), 
            .I3(n27838), .O(n5649[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2096_21 (.CI(n27838), .I0(pwm_setpoint[19]), .I1(GND_net), 
            .CO(n27839));
    SB_LUT4 add_2096_20_lut (.I0(GND_net), .I1(pwm_setpoint[18]), .I2(pwm_setpoint[22]), 
            .I3(n27837), .O(n5649[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_2096_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_2096_20 (.CI(n27837), .I0(pwm_setpoint[18]), .I1(pwm_setpoint[22]), 
            .CO(n27838));
    SB_LUT4 pwm_out_0__I_20_11_lut (.I0(\count[0] [9]), .I1(VCC_net), .I2(VCC_net), 
            .I3(n27880), .O(n10)) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_out_0__I_20_11_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i18027_3_lut (.I0(\half_duty[0] [5]), .I1(half_duty_new[5]), 
            .I2(n1170), .I3(GND_net), .O(n22753));
    defparam i18027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i31784_2_lut (.I0(\count[0] [8]), .I1(\count[0] [6]), .I2(GND_net), 
            .I3(GND_net), .O(n38553));
    defparam i31784_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_970 (.I0(\count[0] [4]), .I1(\count[0] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n12));
    defparam i1_2_lut_adj_970.LUT_INIT = 16'h8888;
    SB_LUT4 i7_4_lut_adj_971 (.I0(n38553), .I1(\count[0] [3]), .I2(\count[0] [10]), 
            .I3(pause_counter_0), .O(n18_adj_3825));
    defparam i7_4_lut_adj_971.LUT_INIT = 16'h0040;
    SB_LUT4 i8_4_lut_adj_972 (.I0(\count[0] [9]), .I1(\count[0] [0]), .I2(\count[0] [1]), 
            .I3(\count[0] [2]), .O(n19));
    defparam i8_4_lut_adj_972.LUT_INIT = 16'h8000;
    SB_LUT4 i10_4_lut_adj_973 (.I0(n19), .I1(\count[0] [7]), .I2(n18_adj_3825), 
            .I3(n12), .O(n1170));
    defparam i10_4_lut_adj_973.LUT_INIT = 16'h2000;
    
endmodule
