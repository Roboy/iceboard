// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Feb 17 2020 11:47:54

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    TX,
    SDA,
    SCL,
    RX,
    NEOPXL,
    LED,
    INLC,
    INLB,
    INLA,
    INHC,
    INHB,
    INHA,
    HALL3,
    HALL2,
    HALL1,
    FAULT_N,
    ENCODER1_B,
    ENCODER1_A,
    ENCODER0_B,
    ENCODER0_A,
    DE,
    CS_MISO,
    CS_CLK,
    CS,
    CLK);

    output USBPU;
    output TX;
    input SDA;
    input SCL;
    input RX;
    output NEOPXL;
    output LED;
    output INLC;
    output INLB;
    output INLA;
    output INHC;
    output INHB;
    output INHA;
    input HALL3;
    input HALL2;
    input HALL1;
    input FAULT_N;
    input ENCODER1_B;
    input ENCODER1_A;
    input ENCODER0_B;
    input ENCODER0_A;
    output DE;
    input CS_MISO;
    output CS_CLK;
    output CS;
    input CLK;

    wire N__56752;
    wire N__56751;
    wire N__56750;
    wire N__56743;
    wire N__56742;
    wire N__56741;
    wire N__56734;
    wire N__56733;
    wire N__56732;
    wire N__56725;
    wire N__56724;
    wire N__56723;
    wire N__56716;
    wire N__56715;
    wire N__56714;
    wire N__56707;
    wire N__56706;
    wire N__56705;
    wire N__56698;
    wire N__56697;
    wire N__56696;
    wire N__56689;
    wire N__56688;
    wire N__56687;
    wire N__56680;
    wire N__56679;
    wire N__56678;
    wire N__56671;
    wire N__56670;
    wire N__56669;
    wire N__56662;
    wire N__56661;
    wire N__56660;
    wire N__56653;
    wire N__56652;
    wire N__56651;
    wire N__56644;
    wire N__56643;
    wire N__56642;
    wire N__56635;
    wire N__56634;
    wire N__56633;
    wire N__56626;
    wire N__56625;
    wire N__56624;
    wire N__56617;
    wire N__56616;
    wire N__56615;
    wire N__56608;
    wire N__56607;
    wire N__56606;
    wire N__56599;
    wire N__56598;
    wire N__56597;
    wire N__56590;
    wire N__56589;
    wire N__56588;
    wire N__56571;
    wire N__56568;
    wire N__56565;
    wire N__56562;
    wire N__56559;
    wire N__56556;
    wire N__56553;
    wire N__56550;
    wire N__56547;
    wire N__56544;
    wire N__56541;
    wire N__56538;
    wire N__56535;
    wire N__56532;
    wire N__56529;
    wire N__56526;
    wire N__56523;
    wire N__56522;
    wire N__56521;
    wire N__56520;
    wire N__56519;
    wire N__56518;
    wire N__56517;
    wire N__56516;
    wire N__56515;
    wire N__56514;
    wire N__56513;
    wire N__56512;
    wire N__56511;
    wire N__56510;
    wire N__56509;
    wire N__56508;
    wire N__56497;
    wire N__56494;
    wire N__56491;
    wire N__56488;
    wire N__56485;
    wire N__56476;
    wire N__56469;
    wire N__56466;
    wire N__56461;
    wire N__56450;
    wire N__56447;
    wire N__56442;
    wire N__56441;
    wire N__56440;
    wire N__56439;
    wire N__56436;
    wire N__56433;
    wire N__56432;
    wire N__56431;
    wire N__56428;
    wire N__56425;
    wire N__56416;
    wire N__56413;
    wire N__56410;
    wire N__56407;
    wire N__56406;
    wire N__56405;
    wire N__56404;
    wire N__56403;
    wire N__56398;
    wire N__56395;
    wire N__56392;
    wire N__56389;
    wire N__56384;
    wire N__56381;
    wire N__56378;
    wire N__56373;
    wire N__56364;
    wire N__56363;
    wire N__56360;
    wire N__56359;
    wire N__56356;
    wire N__56355;
    wire N__56354;
    wire N__56353;
    wire N__56344;
    wire N__56341;
    wire N__56338;
    wire N__56333;
    wire N__56328;
    wire N__56327;
    wire N__56326;
    wire N__56325;
    wire N__56324;
    wire N__56323;
    wire N__56322;
    wire N__56321;
    wire N__56320;
    wire N__56319;
    wire N__56316;
    wire N__56307;
    wire N__56304;
    wire N__56297;
    wire N__56294;
    wire N__56287;
    wire N__56284;
    wire N__56277;
    wire N__56274;
    wire N__56271;
    wire N__56268;
    wire N__56265;
    wire N__56262;
    wire N__56261;
    wire N__56260;
    wire N__56259;
    wire N__56258;
    wire N__56257;
    wire N__56256;
    wire N__56255;
    wire N__56254;
    wire N__56253;
    wire N__56252;
    wire N__56251;
    wire N__56250;
    wire N__56249;
    wire N__56248;
    wire N__56247;
    wire N__56246;
    wire N__56245;
    wire N__56244;
    wire N__56243;
    wire N__56242;
    wire N__56241;
    wire N__56240;
    wire N__56239;
    wire N__56238;
    wire N__56237;
    wire N__56236;
    wire N__56235;
    wire N__56234;
    wire N__56233;
    wire N__56232;
    wire N__56231;
    wire N__56230;
    wire N__56229;
    wire N__56228;
    wire N__56227;
    wire N__56226;
    wire N__56225;
    wire N__56224;
    wire N__56223;
    wire N__56222;
    wire N__56221;
    wire N__56220;
    wire N__56219;
    wire N__56218;
    wire N__56217;
    wire N__56216;
    wire N__56215;
    wire N__56214;
    wire N__56213;
    wire N__56212;
    wire N__56211;
    wire N__56210;
    wire N__56209;
    wire N__56208;
    wire N__56207;
    wire N__56206;
    wire N__56205;
    wire N__56204;
    wire N__56203;
    wire N__56202;
    wire N__56201;
    wire N__56200;
    wire N__56199;
    wire N__56070;
    wire N__56067;
    wire N__56064;
    wire N__56063;
    wire N__56060;
    wire N__56057;
    wire N__56056;
    wire N__56053;
    wire N__56050;
    wire N__56047;
    wire N__56040;
    wire N__56037;
    wire N__56034;
    wire N__56031;
    wire N__56030;
    wire N__56029;
    wire N__56026;
    wire N__56023;
    wire N__56020;
    wire N__56015;
    wire N__56012;
    wire N__56009;
    wire N__56006;
    wire N__56001;
    wire N__55998;
    wire N__55995;
    wire N__55994;
    wire N__55993;
    wire N__55990;
    wire N__55985;
    wire N__55980;
    wire N__55977;
    wire N__55974;
    wire N__55971;
    wire N__55968;
    wire N__55965;
    wire N__55962;
    wire N__55959;
    wire N__55956;
    wire N__55955;
    wire N__55952;
    wire N__55949;
    wire N__55946;
    wire N__55941;
    wire N__55938;
    wire N__55937;
    wire N__55934;
    wire N__55931;
    wire N__55928;
    wire N__55923;
    wire N__55920;
    wire N__55917;
    wire N__55916;
    wire N__55913;
    wire N__55912;
    wire N__55911;
    wire N__55908;
    wire N__55905;
    wire N__55902;
    wire N__55899;
    wire N__55898;
    wire N__55897;
    wire N__55894;
    wire N__55891;
    wire N__55888;
    wire N__55885;
    wire N__55882;
    wire N__55881;
    wire N__55878;
    wire N__55875;
    wire N__55872;
    wire N__55869;
    wire N__55866;
    wire N__55863;
    wire N__55860;
    wire N__55857;
    wire N__55850;
    wire N__55841;
    wire N__55836;
    wire N__55835;
    wire N__55832;
    wire N__55829;
    wire N__55826;
    wire N__55821;
    wire N__55820;
    wire N__55817;
    wire N__55814;
    wire N__55811;
    wire N__55806;
    wire N__55805;
    wire N__55802;
    wire N__55799;
    wire N__55796;
    wire N__55791;
    wire N__55790;
    wire N__55787;
    wire N__55784;
    wire N__55779;
    wire N__55776;
    wire N__55775;
    wire N__55772;
    wire N__55769;
    wire N__55766;
    wire N__55761;
    wire N__55760;
    wire N__55757;
    wire N__55754;
    wire N__55751;
    wire N__55748;
    wire N__55745;
    wire N__55742;
    wire N__55739;
    wire N__55734;
    wire N__55731;
    wire N__55728;
    wire N__55725;
    wire N__55722;
    wire N__55719;
    wire N__55716;
    wire N__55715;
    wire N__55712;
    wire N__55709;
    wire N__55706;
    wire N__55701;
    wire N__55698;
    wire N__55695;
    wire N__55694;
    wire N__55691;
    wire N__55688;
    wire N__55685;
    wire N__55680;
    wire N__55677;
    wire N__55674;
    wire N__55671;
    wire N__55668;
    wire N__55667;
    wire N__55664;
    wire N__55661;
    wire N__55658;
    wire N__55653;
    wire N__55650;
    wire N__55647;
    wire N__55646;
    wire N__55643;
    wire N__55640;
    wire N__55637;
    wire N__55632;
    wire N__55629;
    wire N__55626;
    wire N__55625;
    wire N__55622;
    wire N__55619;
    wire N__55616;
    wire N__55611;
    wire N__55608;
    wire N__55605;
    wire N__55602;
    wire N__55599;
    wire N__55596;
    wire N__55593;
    wire N__55592;
    wire N__55591;
    wire N__55588;
    wire N__55583;
    wire N__55580;
    wire N__55575;
    wire N__55572;
    wire N__55569;
    wire N__55566;
    wire N__55563;
    wire N__55562;
    wire N__55559;
    wire N__55558;
    wire N__55557;
    wire N__55556;
    wire N__55555;
    wire N__55554;
    wire N__55553;
    wire N__55552;
    wire N__55551;
    wire N__55550;
    wire N__55549;
    wire N__55548;
    wire N__55547;
    wire N__55546;
    wire N__55545;
    wire N__55544;
    wire N__55543;
    wire N__55542;
    wire N__55541;
    wire N__55540;
    wire N__55539;
    wire N__55538;
    wire N__55537;
    wire N__55536;
    wire N__55535;
    wire N__55534;
    wire N__55533;
    wire N__55532;
    wire N__55531;
    wire N__55530;
    wire N__55529;
    wire N__55528;
    wire N__55527;
    wire N__55526;
    wire N__55521;
    wire N__55518;
    wire N__55515;
    wire N__55512;
    wire N__55509;
    wire N__55506;
    wire N__55503;
    wire N__55500;
    wire N__55497;
    wire N__55496;
    wire N__55495;
    wire N__55494;
    wire N__55493;
    wire N__55492;
    wire N__55491;
    wire N__55490;
    wire N__55487;
    wire N__55486;
    wire N__55485;
    wire N__55482;
    wire N__55479;
    wire N__55478;
    wire N__55477;
    wire N__55476;
    wire N__55473;
    wire N__55470;
    wire N__55463;
    wire N__55456;
    wire N__55455;
    wire N__55454;
    wire N__55453;
    wire N__55450;
    wire N__55447;
    wire N__55446;
    wire N__55445;
    wire N__55444;
    wire N__55441;
    wire N__55438;
    wire N__55437;
    wire N__55436;
    wire N__55435;
    wire N__55434;
    wire N__55433;
    wire N__55432;
    wire N__55431;
    wire N__55428;
    wire N__55427;
    wire N__55426;
    wire N__55425;
    wire N__55422;
    wire N__55421;
    wire N__55420;
    wire N__55419;
    wire N__55418;
    wire N__55415;
    wire N__55412;
    wire N__55409;
    wire N__55406;
    wire N__55403;
    wire N__55400;
    wire N__55397;
    wire N__55394;
    wire N__55393;
    wire N__55392;
    wire N__55389;
    wire N__55380;
    wire N__55371;
    wire N__55368;
    wire N__55361;
    wire N__55358;
    wire N__55357;
    wire N__55356;
    wire N__55355;
    wire N__55352;
    wire N__55351;
    wire N__55350;
    wire N__55349;
    wire N__55348;
    wire N__55347;
    wire N__55346;
    wire N__55345;
    wire N__55344;
    wire N__55341;
    wire N__55340;
    wire N__55333;
    wire N__55322;
    wire N__55319;
    wire N__55312;
    wire N__55305;
    wire N__55294;
    wire N__55289;
    wire N__55288;
    wire N__55287;
    wire N__55286;
    wire N__55285;
    wire N__55284;
    wire N__55283;
    wire N__55282;
    wire N__55281;
    wire N__55280;
    wire N__55279;
    wire N__55278;
    wire N__55277;
    wire N__55276;
    wire N__55275;
    wire N__55270;
    wire N__55263;
    wire N__55252;
    wire N__55241;
    wire N__55240;
    wire N__55237;
    wire N__55228;
    wire N__55219;
    wire N__55218;
    wire N__55215;
    wire N__55214;
    wire N__55213;
    wire N__55212;
    wire N__55211;
    wire N__55210;
    wire N__55209;
    wire N__55206;
    wire N__55205;
    wire N__55204;
    wire N__55203;
    wire N__55192;
    wire N__55183;
    wire N__55174;
    wire N__55167;
    wire N__55166;
    wire N__55165;
    wire N__55164;
    wire N__55161;
    wire N__55160;
    wire N__55159;
    wire N__55158;
    wire N__55157;
    wire N__55152;
    wire N__55151;
    wire N__55148;
    wire N__55141;
    wire N__55132;
    wire N__55131;
    wire N__55130;
    wire N__55129;
    wire N__55128;
    wire N__55127;
    wire N__55126;
    wire N__55125;
    wire N__55122;
    wire N__55121;
    wire N__55120;
    wire N__55119;
    wire N__55118;
    wire N__55117;
    wire N__55110;
    wire N__55101;
    wire N__55098;
    wire N__55097;
    wire N__55096;
    wire N__55093;
    wire N__55092;
    wire N__55091;
    wire N__55088;
    wire N__55087;
    wire N__55086;
    wire N__55085;
    wire N__55084;
    wire N__55083;
    wire N__55082;
    wire N__55081;
    wire N__55080;
    wire N__55079;
    wire N__55078;
    wire N__55077;
    wire N__55076;
    wire N__55073;
    wire N__55070;
    wire N__55067;
    wire N__55066;
    wire N__55065;
    wire N__55064;
    wire N__55063;
    wire N__55062;
    wire N__55061;
    wire N__55060;
    wire N__55059;
    wire N__55058;
    wire N__55057;
    wire N__55056;
    wire N__55055;
    wire N__55046;
    wire N__55045;
    wire N__55042;
    wire N__55041;
    wire N__55040;
    wire N__55039;
    wire N__55038;
    wire N__55037;
    wire N__55036;
    wire N__55035;
    wire N__55034;
    wire N__55033;
    wire N__55032;
    wire N__55031;
    wire N__55030;
    wire N__55023;
    wire N__55020;
    wire N__55011;
    wire N__55004;
    wire N__54995;
    wire N__54988;
    wire N__54985;
    wire N__54974;
    wire N__54967;
    wire N__54964;
    wire N__54959;
    wire N__54958;
    wire N__54957;
    wire N__54956;
    wire N__54955;
    wire N__54954;
    wire N__54953;
    wire N__54952;
    wire N__54947;
    wire N__54944;
    wire N__54937;
    wire N__54932;
    wire N__54925;
    wire N__54922;
    wire N__54915;
    wire N__54908;
    wire N__54903;
    wire N__54894;
    wire N__54893;
    wire N__54892;
    wire N__54891;
    wire N__54890;
    wire N__54887;
    wire N__54884;
    wire N__54883;
    wire N__54882;
    wire N__54881;
    wire N__54880;
    wire N__54879;
    wire N__54878;
    wire N__54877;
    wire N__54876;
    wire N__54875;
    wire N__54874;
    wire N__54873;
    wire N__54872;
    wire N__54871;
    wire N__54870;
    wire N__54869;
    wire N__54868;
    wire N__54867;
    wire N__54866;
    wire N__54865;
    wire N__54864;
    wire N__54863;
    wire N__54862;
    wire N__54861;
    wire N__54860;
    wire N__54857;
    wire N__54854;
    wire N__54851;
    wire N__54848;
    wire N__54845;
    wire N__54842;
    wire N__54839;
    wire N__54836;
    wire N__54833;
    wire N__54830;
    wire N__54823;
    wire N__54820;
    wire N__54817;
    wire N__54814;
    wire N__54813;
    wire N__54810;
    wire N__54807;
    wire N__54804;
    wire N__54801;
    wire N__54798;
    wire N__54795;
    wire N__54794;
    wire N__54793;
    wire N__54792;
    wire N__54789;
    wire N__54788;
    wire N__54787;
    wire N__54786;
    wire N__54785;
    wire N__54784;
    wire N__54783;
    wire N__54780;
    wire N__54777;
    wire N__54776;
    wire N__54773;
    wire N__54770;
    wire N__54767;
    wire N__54764;
    wire N__54763;
    wire N__54762;
    wire N__54759;
    wire N__54758;
    wire N__54757;
    wire N__54756;
    wire N__54753;
    wire N__54750;
    wire N__54747;
    wire N__54746;
    wire N__54745;
    wire N__54744;
    wire N__54743;
    wire N__54740;
    wire N__54737;
    wire N__54736;
    wire N__54733;
    wire N__54732;
    wire N__54731;
    wire N__54730;
    wire N__54729;
    wire N__54728;
    wire N__54727;
    wire N__54726;
    wire N__54725;
    wire N__54724;
    wire N__54723;
    wire N__54722;
    wire N__54721;
    wire N__54714;
    wire N__54713;
    wire N__54710;
    wire N__54709;
    wire N__54708;
    wire N__54707;
    wire N__54706;
    wire N__54705;
    wire N__54702;
    wire N__54701;
    wire N__54700;
    wire N__54695;
    wire N__54690;
    wire N__54677;
    wire N__54668;
    wire N__54663;
    wire N__54662;
    wire N__54661;
    wire N__54658;
    wire N__54657;
    wire N__54656;
    wire N__54655;
    wire N__54654;
    wire N__54653;
    wire N__54652;
    wire N__54651;
    wire N__54650;
    wire N__54649;
    wire N__54648;
    wire N__54647;
    wire N__54646;
    wire N__54645;
    wire N__54644;
    wire N__54643;
    wire N__54640;
    wire N__54627;
    wire N__54624;
    wire N__54621;
    wire N__54618;
    wire N__54615;
    wire N__54608;
    wire N__54603;
    wire N__54596;
    wire N__54593;
    wire N__54592;
    wire N__54591;
    wire N__54590;
    wire N__54589;
    wire N__54588;
    wire N__54587;
    wire N__54586;
    wire N__54583;
    wire N__54582;
    wire N__54581;
    wire N__54580;
    wire N__54579;
    wire N__54578;
    wire N__54577;
    wire N__54576;
    wire N__54575;
    wire N__54574;
    wire N__54573;
    wire N__54572;
    wire N__54569;
    wire N__54566;
    wire N__54565;
    wire N__54564;
    wire N__54561;
    wire N__54558;
    wire N__54557;
    wire N__54556;
    wire N__54553;
    wire N__54550;
    wire N__54547;
    wire N__54544;
    wire N__54541;
    wire N__54538;
    wire N__54535;
    wire N__54534;
    wire N__54531;
    wire N__54528;
    wire N__54525;
    wire N__54522;
    wire N__54519;
    wire N__54516;
    wire N__54515;
    wire N__54512;
    wire N__54509;
    wire N__54508;
    wire N__54507;
    wire N__54506;
    wire N__54499;
    wire N__54492;
    wire N__54483;
    wire N__54480;
    wire N__54477;
    wire N__54466;
    wire N__54457;
    wire N__54452;
    wire N__54447;
    wire N__54446;
    wire N__54445;
    wire N__54444;
    wire N__54443;
    wire N__54438;
    wire N__54431;
    wire N__54424;
    wire N__54423;
    wire N__54422;
    wire N__54421;
    wire N__54418;
    wire N__54417;
    wire N__54416;
    wire N__54415;
    wire N__54414;
    wire N__54407;
    wire N__54402;
    wire N__54391;
    wire N__54382;
    wire N__54381;
    wire N__54380;
    wire N__54379;
    wire N__54376;
    wire N__54375;
    wire N__54374;
    wire N__54373;
    wire N__54370;
    wire N__54369;
    wire N__54368;
    wire N__54367;
    wire N__54364;
    wire N__54357;
    wire N__54352;
    wire N__54351;
    wire N__54348;
    wire N__54347;
    wire N__54346;
    wire N__54345;
    wire N__54342;
    wire N__54339;
    wire N__54336;
    wire N__54333;
    wire N__54330;
    wire N__54329;
    wire N__54328;
    wire N__54327;
    wire N__54326;
    wire N__54325;
    wire N__54324;
    wire N__54321;
    wire N__54318;
    wire N__54315;
    wire N__54312;
    wire N__54309;
    wire N__54306;
    wire N__54297;
    wire N__54294;
    wire N__54293;
    wire N__54292;
    wire N__54289;
    wire N__54288;
    wire N__54287;
    wire N__54284;
    wire N__54283;
    wire N__54280;
    wire N__54275;
    wire N__54270;
    wire N__54263;
    wire N__54258;
    wire N__54253;
    wire N__54252;
    wire N__54249;
    wire N__54248;
    wire N__54247;
    wire N__54246;
    wire N__54245;
    wire N__54244;
    wire N__54243;
    wire N__54242;
    wire N__54241;
    wire N__54240;
    wire N__54237;
    wire N__54236;
    wire N__54233;
    wire N__54230;
    wire N__54223;
    wire N__54218;
    wire N__54215;
    wire N__54212;
    wire N__54205;
    wire N__54186;
    wire N__54177;
    wire N__54168;
    wire N__54163;
    wire N__54154;
    wire N__54145;
    wire N__54140;
    wire N__54131;
    wire N__54122;
    wire N__54113;
    wire N__54106;
    wire N__54095;
    wire N__54090;
    wire N__54083;
    wire N__54076;
    wire N__54075;
    wire N__54074;
    wire N__54067;
    wire N__54058;
    wire N__54053;
    wire N__54050;
    wire N__54043;
    wire N__54036;
    wire N__54025;
    wire N__54024;
    wire N__54023;
    wire N__54022;
    wire N__54021;
    wire N__54020;
    wire N__54017;
    wire N__54014;
    wire N__54011;
    wire N__54010;
    wire N__54001;
    wire N__53994;
    wire N__53983;
    wire N__53982;
    wire N__53979;
    wire N__53978;
    wire N__53977;
    wire N__53976;
    wire N__53975;
    wire N__53972;
    wire N__53969;
    wire N__53968;
    wire N__53967;
    wire N__53960;
    wire N__53957;
    wire N__53950;
    wire N__53945;
    wire N__53936;
    wire N__53935;
    wire N__53932;
    wire N__53929;
    wire N__53926;
    wire N__53923;
    wire N__53920;
    wire N__53919;
    wire N__53918;
    wire N__53917;
    wire N__53910;
    wire N__53903;
    wire N__53898;
    wire N__53891;
    wire N__53880;
    wire N__53875;
    wire N__53868;
    wire N__53865;
    wire N__53856;
    wire N__53855;
    wire N__53852;
    wire N__53851;
    wire N__53850;
    wire N__53847;
    wire N__53846;
    wire N__53843;
    wire N__53842;
    wire N__53841;
    wire N__53838;
    wire N__53835;
    wire N__53834;
    wire N__53831;
    wire N__53828;
    wire N__53825;
    wire N__53820;
    wire N__53819;
    wire N__53818;
    wire N__53817;
    wire N__53816;
    wire N__53815;
    wire N__53814;
    wire N__53813;
    wire N__53810;
    wire N__53799;
    wire N__53792;
    wire N__53791;
    wire N__53790;
    wire N__53789;
    wire N__53788;
    wire N__53787;
    wire N__53786;
    wire N__53785;
    wire N__53778;
    wire N__53761;
    wire N__53758;
    wire N__53753;
    wire N__53742;
    wire N__53737;
    wire N__53728;
    wire N__53717;
    wire N__53710;
    wire N__53705;
    wire N__53696;
    wire N__53689;
    wire N__53686;
    wire N__53677;
    wire N__53674;
    wire N__53667;
    wire N__53660;
    wire N__53659;
    wire N__53656;
    wire N__53653;
    wire N__53650;
    wire N__53649;
    wire N__53648;
    wire N__53647;
    wire N__53646;
    wire N__53635;
    wire N__53630;
    wire N__53625;
    wire N__53616;
    wire N__53605;
    wire N__53594;
    wire N__53589;
    wire N__53586;
    wire N__53579;
    wire N__53572;
    wire N__53565;
    wire N__53562;
    wire N__53557;
    wire N__53552;
    wire N__53547;
    wire N__53542;
    wire N__53537;
    wire N__53528;
    wire N__53519;
    wire N__53516;
    wire N__53513;
    wire N__53506;
    wire N__53497;
    wire N__53494;
    wire N__53491;
    wire N__53488;
    wire N__53485;
    wire N__53482;
    wire N__53477;
    wire N__53472;
    wire N__53461;
    wire N__53450;
    wire N__53445;
    wire N__53440;
    wire N__53435;
    wire N__53430;
    wire N__53421;
    wire N__53418;
    wire N__53415;
    wire N__53408;
    wire N__53403;
    wire N__53396;
    wire N__53385;
    wire N__53384;
    wire N__53381;
    wire N__53378;
    wire N__53377;
    wire N__53374;
    wire N__53371;
    wire N__53368;
    wire N__53365;
    wire N__53358;
    wire N__53355;
    wire N__53352;
    wire N__53349;
    wire N__53346;
    wire N__53345;
    wire N__53342;
    wire N__53339;
    wire N__53336;
    wire N__53331;
    wire N__53328;
    wire N__53327;
    wire N__53324;
    wire N__53321;
    wire N__53318;
    wire N__53313;
    wire N__53310;
    wire N__53309;
    wire N__53306;
    wire N__53303;
    wire N__53300;
    wire N__53295;
    wire N__53292;
    wire N__53289;
    wire N__53286;
    wire N__53285;
    wire N__53282;
    wire N__53279;
    wire N__53276;
    wire N__53271;
    wire N__53268;
    wire N__53265;
    wire N__53264;
    wire N__53261;
    wire N__53258;
    wire N__53255;
    wire N__53250;
    wire N__53247;
    wire N__53246;
    wire N__53243;
    wire N__53240;
    wire N__53237;
    wire N__53232;
    wire N__53229;
    wire N__53226;
    wire N__53223;
    wire N__53222;
    wire N__53221;
    wire N__53218;
    wire N__53215;
    wire N__53212;
    wire N__53209;
    wire N__53206;
    wire N__53203;
    wire N__53200;
    wire N__53193;
    wire N__53190;
    wire N__53187;
    wire N__53184;
    wire N__53181;
    wire N__53180;
    wire N__53179;
    wire N__53176;
    wire N__53175;
    wire N__53174;
    wire N__53173;
    wire N__53172;
    wire N__53171;
    wire N__53168;
    wire N__53167;
    wire N__53166;
    wire N__53163;
    wire N__53162;
    wire N__53159;
    wire N__53156;
    wire N__53153;
    wire N__53150;
    wire N__53145;
    wire N__53134;
    wire N__53121;
    wire N__53118;
    wire N__53115;
    wire N__53114;
    wire N__53113;
    wire N__53110;
    wire N__53107;
    wire N__53104;
    wire N__53101;
    wire N__53096;
    wire N__53091;
    wire N__53088;
    wire N__53085;
    wire N__53084;
    wire N__53083;
    wire N__53080;
    wire N__53075;
    wire N__53070;
    wire N__53067;
    wire N__53064;
    wire N__53061;
    wire N__53058;
    wire N__53055;
    wire N__53052;
    wire N__53051;
    wire N__53050;
    wire N__53047;
    wire N__53042;
    wire N__53039;
    wire N__53034;
    wire N__53031;
    wire N__53028;
    wire N__53025;
    wire N__53022;
    wire N__53021;
    wire N__53018;
    wire N__53017;
    wire N__53014;
    wire N__53011;
    wire N__53008;
    wire N__53005;
    wire N__53002;
    wire N__52995;
    wire N__52992;
    wire N__52989;
    wire N__52986;
    wire N__52983;
    wire N__52980;
    wire N__52979;
    wire N__52976;
    wire N__52973;
    wire N__52972;
    wire N__52969;
    wire N__52966;
    wire N__52963;
    wire N__52960;
    wire N__52953;
    wire N__52950;
    wire N__52947;
    wire N__52944;
    wire N__52941;
    wire N__52938;
    wire N__52937;
    wire N__52934;
    wire N__52931;
    wire N__52930;
    wire N__52927;
    wire N__52924;
    wire N__52921;
    wire N__52918;
    wire N__52911;
    wire N__52908;
    wire N__52905;
    wire N__52902;
    wire N__52899;
    wire N__52896;
    wire N__52895;
    wire N__52892;
    wire N__52889;
    wire N__52886;
    wire N__52885;
    wire N__52880;
    wire N__52877;
    wire N__52874;
    wire N__52869;
    wire N__52866;
    wire N__52863;
    wire N__52860;
    wire N__52859;
    wire N__52856;
    wire N__52853;
    wire N__52852;
    wire N__52849;
    wire N__52846;
    wire N__52843;
    wire N__52840;
    wire N__52833;
    wire N__52830;
    wire N__52827;
    wire N__52824;
    wire N__52821;
    wire N__52820;
    wire N__52817;
    wire N__52814;
    wire N__52813;
    wire N__52810;
    wire N__52807;
    wire N__52804;
    wire N__52799;
    wire N__52794;
    wire N__52791;
    wire N__52788;
    wire N__52785;
    wire N__52782;
    wire N__52781;
    wire N__52778;
    wire N__52775;
    wire N__52774;
    wire N__52771;
    wire N__52768;
    wire N__52765;
    wire N__52762;
    wire N__52755;
    wire N__52752;
    wire N__52749;
    wire N__52746;
    wire N__52745;
    wire N__52742;
    wire N__52739;
    wire N__52736;
    wire N__52733;
    wire N__52732;
    wire N__52727;
    wire N__52724;
    wire N__52719;
    wire N__52716;
    wire N__52713;
    wire N__52710;
    wire N__52709;
    wire N__52706;
    wire N__52703;
    wire N__52700;
    wire N__52697;
    wire N__52692;
    wire N__52689;
    wire N__52686;
    wire N__52683;
    wire N__52680;
    wire N__52679;
    wire N__52678;
    wire N__52675;
    wire N__52670;
    wire N__52665;
    wire N__52662;
    wire N__52659;
    wire N__52656;
    wire N__52653;
    wire N__52652;
    wire N__52649;
    wire N__52646;
    wire N__52641;
    wire N__52638;
    wire N__52635;
    wire N__52632;
    wire N__52629;
    wire N__52626;
    wire N__52623;
    wire N__52620;
    wire N__52619;
    wire N__52616;
    wire N__52613;
    wire N__52608;
    wire N__52605;
    wire N__52602;
    wire N__52601;
    wire N__52598;
    wire N__52595;
    wire N__52592;
    wire N__52589;
    wire N__52584;
    wire N__52581;
    wire N__52578;
    wire N__52577;
    wire N__52574;
    wire N__52571;
    wire N__52568;
    wire N__52565;
    wire N__52562;
    wire N__52559;
    wire N__52554;
    wire N__52551;
    wire N__52548;
    wire N__52545;
    wire N__52542;
    wire N__52539;
    wire N__52536;
    wire N__52533;
    wire N__52532;
    wire N__52529;
    wire N__52526;
    wire N__52525;
    wire N__52522;
    wire N__52519;
    wire N__52516;
    wire N__52509;
    wire N__52506;
    wire N__52503;
    wire N__52500;
    wire N__52497;
    wire N__52496;
    wire N__52493;
    wire N__52490;
    wire N__52487;
    wire N__52484;
    wire N__52479;
    wire N__52476;
    wire N__52475;
    wire N__52472;
    wire N__52469;
    wire N__52466;
    wire N__52463;
    wire N__52460;
    wire N__52457;
    wire N__52454;
    wire N__52451;
    wire N__52446;
    wire N__52443;
    wire N__52440;
    wire N__52439;
    wire N__52436;
    wire N__52433;
    wire N__52430;
    wire N__52427;
    wire N__52424;
    wire N__52421;
    wire N__52416;
    wire N__52413;
    wire N__52410;
    wire N__52409;
    wire N__52408;
    wire N__52405;
    wire N__52402;
    wire N__52399;
    wire N__52394;
    wire N__52389;
    wire N__52386;
    wire N__52383;
    wire N__52380;
    wire N__52377;
    wire N__52374;
    wire N__52371;
    wire N__52368;
    wire N__52365;
    wire N__52362;
    wire N__52359;
    wire N__52356;
    wire N__52353;
    wire N__52350;
    wire N__52349;
    wire N__52348;
    wire N__52347;
    wire N__52344;
    wire N__52343;
    wire N__52342;
    wire N__52339;
    wire N__52338;
    wire N__52337;
    wire N__52336;
    wire N__52333;
    wire N__52332;
    wire N__52331;
    wire N__52328;
    wire N__52327;
    wire N__52324;
    wire N__52319;
    wire N__52314;
    wire N__52311;
    wire N__52304;
    wire N__52301;
    wire N__52296;
    wire N__52281;
    wire N__52280;
    wire N__52277;
    wire N__52276;
    wire N__52273;
    wire N__52270;
    wire N__52267;
    wire N__52264;
    wire N__52261;
    wire N__52258;
    wire N__52255;
    wire N__52248;
    wire N__52247;
    wire N__52246;
    wire N__52243;
    wire N__52240;
    wire N__52237;
    wire N__52230;
    wire N__52227;
    wire N__52224;
    wire N__52221;
    wire N__52218;
    wire N__52215;
    wire N__52214;
    wire N__52211;
    wire N__52208;
    wire N__52205;
    wire N__52202;
    wire N__52199;
    wire N__52194;
    wire N__52191;
    wire N__52188;
    wire N__52185;
    wire N__52182;
    wire N__52179;
    wire N__52178;
    wire N__52177;
    wire N__52174;
    wire N__52171;
    wire N__52168;
    wire N__52165;
    wire N__52158;
    wire N__52155;
    wire N__52152;
    wire N__52149;
    wire N__52148;
    wire N__52145;
    wire N__52142;
    wire N__52141;
    wire N__52138;
    wire N__52135;
    wire N__52132;
    wire N__52125;
    wire N__52122;
    wire N__52119;
    wire N__52116;
    wire N__52113;
    wire N__52110;
    wire N__52109;
    wire N__52106;
    wire N__52105;
    wire N__52102;
    wire N__52099;
    wire N__52096;
    wire N__52089;
    wire N__52086;
    wire N__52083;
    wire N__52080;
    wire N__52077;
    wire N__52076;
    wire N__52075;
    wire N__52072;
    wire N__52069;
    wire N__52066;
    wire N__52063;
    wire N__52060;
    wire N__52057;
    wire N__52050;
    wire N__52047;
    wire N__52044;
    wire N__52041;
    wire N__52038;
    wire N__52035;
    wire N__52034;
    wire N__52031;
    wire N__52028;
    wire N__52027;
    wire N__52024;
    wire N__52021;
    wire N__52018;
    wire N__52011;
    wire N__52008;
    wire N__52005;
    wire N__52002;
    wire N__51999;
    wire N__51996;
    wire N__51993;
    wire N__51992;
    wire N__51989;
    wire N__51986;
    wire N__51985;
    wire N__51982;
    wire N__51979;
    wire N__51976;
    wire N__51969;
    wire N__51966;
    wire N__51963;
    wire N__51960;
    wire N__51957;
    wire N__51954;
    wire N__51953;
    wire N__51950;
    wire N__51947;
    wire N__51944;
    wire N__51943;
    wire N__51940;
    wire N__51937;
    wire N__51934;
    wire N__51927;
    wire N__51924;
    wire N__51921;
    wire N__51918;
    wire N__51915;
    wire N__51912;
    wire N__51909;
    wire N__51906;
    wire N__51905;
    wire N__51904;
    wire N__51901;
    wire N__51896;
    wire N__51891;
    wire N__51888;
    wire N__51885;
    wire N__51882;
    wire N__51879;
    wire N__51876;
    wire N__51873;
    wire N__51870;
    wire N__51867;
    wire N__51866;
    wire N__51863;
    wire N__51860;
    wire N__51855;
    wire N__51854;
    wire N__51851;
    wire N__51848;
    wire N__51843;
    wire N__51840;
    wire N__51837;
    wire N__51834;
    wire N__51833;
    wire N__51830;
    wire N__51827;
    wire N__51824;
    wire N__51821;
    wire N__51816;
    wire N__51815;
    wire N__51812;
    wire N__51809;
    wire N__51804;
    wire N__51801;
    wire N__51798;
    wire N__51795;
    wire N__51792;
    wire N__51791;
    wire N__51788;
    wire N__51785;
    wire N__51782;
    wire N__51781;
    wire N__51778;
    wire N__51775;
    wire N__51772;
    wire N__51765;
    wire N__51762;
    wire N__51759;
    wire N__51756;
    wire N__51753;
    wire N__51750;
    wire N__51747;
    wire N__51746;
    wire N__51743;
    wire N__51740;
    wire N__51735;
    wire N__51732;
    wire N__51729;
    wire N__51728;
    wire N__51725;
    wire N__51722;
    wire N__51717;
    wire N__51714;
    wire N__51711;
    wire N__51710;
    wire N__51707;
    wire N__51706;
    wire N__51703;
    wire N__51700;
    wire N__51697;
    wire N__51694;
    wire N__51689;
    wire N__51686;
    wire N__51683;
    wire N__51678;
    wire N__51675;
    wire N__51672;
    wire N__51669;
    wire N__51666;
    wire N__51663;
    wire N__51662;
    wire N__51659;
    wire N__51658;
    wire N__51655;
    wire N__51652;
    wire N__51649;
    wire N__51642;
    wire N__51639;
    wire N__51636;
    wire N__51633;
    wire N__51630;
    wire N__51627;
    wire N__51626;
    wire N__51623;
    wire N__51622;
    wire N__51619;
    wire N__51616;
    wire N__51613;
    wire N__51606;
    wire N__51603;
    wire N__51600;
    wire N__51597;
    wire N__51594;
    wire N__51591;
    wire N__51590;
    wire N__51587;
    wire N__51584;
    wire N__51581;
    wire N__51578;
    wire N__51573;
    wire N__51570;
    wire N__51567;
    wire N__51564;
    wire N__51561;
    wire N__51558;
    wire N__51557;
    wire N__51554;
    wire N__51551;
    wire N__51548;
    wire N__51545;
    wire N__51542;
    wire N__51539;
    wire N__51538;
    wire N__51535;
    wire N__51532;
    wire N__51529;
    wire N__51526;
    wire N__51519;
    wire N__51516;
    wire N__51513;
    wire N__51510;
    wire N__51507;
    wire N__51504;
    wire N__51503;
    wire N__51500;
    wire N__51497;
    wire N__51494;
    wire N__51489;
    wire N__51486;
    wire N__51483;
    wire N__51480;
    wire N__51477;
    wire N__51476;
    wire N__51473;
    wire N__51470;
    wire N__51467;
    wire N__51466;
    wire N__51461;
    wire N__51458;
    wire N__51455;
    wire N__51450;
    wire N__51447;
    wire N__51444;
    wire N__51441;
    wire N__51440;
    wire N__51437;
    wire N__51434;
    wire N__51431;
    wire N__51428;
    wire N__51425;
    wire N__51420;
    wire N__51417;
    wire N__51414;
    wire N__51411;
    wire N__51408;
    wire N__51405;
    wire N__51402;
    wire N__51399;
    wire N__51396;
    wire N__51393;
    wire N__51392;
    wire N__51389;
    wire N__51388;
    wire N__51385;
    wire N__51382;
    wire N__51379;
    wire N__51372;
    wire N__51369;
    wire N__51366;
    wire N__51363;
    wire N__51360;
    wire N__51357;
    wire N__51356;
    wire N__51353;
    wire N__51350;
    wire N__51347;
    wire N__51342;
    wire N__51339;
    wire N__51336;
    wire N__51333;
    wire N__51332;
    wire N__51329;
    wire N__51326;
    wire N__51325;
    wire N__51322;
    wire N__51319;
    wire N__51316;
    wire N__51309;
    wire N__51306;
    wire N__51303;
    wire N__51300;
    wire N__51297;
    wire N__51296;
    wire N__51293;
    wire N__51292;
    wire N__51291;
    wire N__51288;
    wire N__51285;
    wire N__51280;
    wire N__51273;
    wire N__51270;
    wire N__51267;
    wire N__51266;
    wire N__51265;
    wire N__51264;
    wire N__51261;
    wire N__51256;
    wire N__51253;
    wire N__51250;
    wire N__51247;
    wire N__51244;
    wire N__51241;
    wire N__51238;
    wire N__51231;
    wire N__51228;
    wire N__51227;
    wire N__51224;
    wire N__51221;
    wire N__51220;
    wire N__51217;
    wire N__51216;
    wire N__51213;
    wire N__51210;
    wire N__51207;
    wire N__51204;
    wire N__51201;
    wire N__51192;
    wire N__51189;
    wire N__51188;
    wire N__51187;
    wire N__51186;
    wire N__51185;
    wire N__51182;
    wire N__51181;
    wire N__51178;
    wire N__51177;
    wire N__51174;
    wire N__51173;
    wire N__51170;
    wire N__51169;
    wire N__51168;
    wire N__51167;
    wire N__51166;
    wire N__51165;
    wire N__51164;
    wire N__51161;
    wire N__51144;
    wire N__51143;
    wire N__51140;
    wire N__51139;
    wire N__51136;
    wire N__51135;
    wire N__51132;
    wire N__51131;
    wire N__51128;
    wire N__51127;
    wire N__51126;
    wire N__51125;
    wire N__51122;
    wire N__51121;
    wire N__51120;
    wire N__51119;
    wire N__51118;
    wire N__51117;
    wire N__51116;
    wire N__51115;
    wire N__51110;
    wire N__51093;
    wire N__51084;
    wire N__51075;
    wire N__51068;
    wire N__51057;
    wire N__51054;
    wire N__51051;
    wire N__51050;
    wire N__51049;
    wire N__51046;
    wire N__51043;
    wire N__51040;
    wire N__51039;
    wire N__51038;
    wire N__51037;
    wire N__51034;
    wire N__51031;
    wire N__51028;
    wire N__51025;
    wire N__51022;
    wire N__51019;
    wire N__51016;
    wire N__51013;
    wire N__51006;
    wire N__50997;
    wire N__50994;
    wire N__50991;
    wire N__50988;
    wire N__50985;
    wire N__50982;
    wire N__50981;
    wire N__50980;
    wire N__50977;
    wire N__50974;
    wire N__50971;
    wire N__50964;
    wire N__50961;
    wire N__50958;
    wire N__50955;
    wire N__50952;
    wire N__50951;
    wire N__50950;
    wire N__50947;
    wire N__50944;
    wire N__50941;
    wire N__50934;
    wire N__50933;
    wire N__50930;
    wire N__50927;
    wire N__50924;
    wire N__50919;
    wire N__50916;
    wire N__50913;
    wire N__50910;
    wire N__50909;
    wire N__50908;
    wire N__50907;
    wire N__50906;
    wire N__50905;
    wire N__50902;
    wire N__50901;
    wire N__50900;
    wire N__50899;
    wire N__50896;
    wire N__50895;
    wire N__50894;
    wire N__50893;
    wire N__50892;
    wire N__50885;
    wire N__50882;
    wire N__50879;
    wire N__50874;
    wire N__50873;
    wire N__50870;
    wire N__50869;
    wire N__50868;
    wire N__50867;
    wire N__50864;
    wire N__50863;
    wire N__50858;
    wire N__50853;
    wire N__50850;
    wire N__50847;
    wire N__50842;
    wire N__50839;
    wire N__50838;
    wire N__50837;
    wire N__50836;
    wire N__50835;
    wire N__50834;
    wire N__50833;
    wire N__50832;
    wire N__50829;
    wire N__50822;
    wire N__50819;
    wire N__50816;
    wire N__50811;
    wire N__50806;
    wire N__50801;
    wire N__50798;
    wire N__50795;
    wire N__50792;
    wire N__50789;
    wire N__50782;
    wire N__50773;
    wire N__50754;
    wire N__50751;
    wire N__50750;
    wire N__50747;
    wire N__50744;
    wire N__50743;
    wire N__50740;
    wire N__50737;
    wire N__50734;
    wire N__50731;
    wire N__50728;
    wire N__50725;
    wire N__50718;
    wire N__50715;
    wire N__50712;
    wire N__50709;
    wire N__50706;
    wire N__50705;
    wire N__50704;
    wire N__50701;
    wire N__50700;
    wire N__50697;
    wire N__50694;
    wire N__50691;
    wire N__50686;
    wire N__50679;
    wire N__50676;
    wire N__50675;
    wire N__50674;
    wire N__50671;
    wire N__50670;
    wire N__50667;
    wire N__50664;
    wire N__50661;
    wire N__50658;
    wire N__50655;
    wire N__50652;
    wire N__50647;
    wire N__50640;
    wire N__50637;
    wire N__50634;
    wire N__50631;
    wire N__50630;
    wire N__50629;
    wire N__50626;
    wire N__50625;
    wire N__50622;
    wire N__50619;
    wire N__50616;
    wire N__50613;
    wire N__50610;
    wire N__50601;
    wire N__50598;
    wire N__50597;
    wire N__50594;
    wire N__50591;
    wire N__50588;
    wire N__50587;
    wire N__50586;
    wire N__50583;
    wire N__50580;
    wire N__50575;
    wire N__50568;
    wire N__50565;
    wire N__50562;
    wire N__50559;
    wire N__50558;
    wire N__50557;
    wire N__50554;
    wire N__50551;
    wire N__50548;
    wire N__50545;
    wire N__50544;
    wire N__50541;
    wire N__50538;
    wire N__50535;
    wire N__50532;
    wire N__50527;
    wire N__50520;
    wire N__50517;
    wire N__50514;
    wire N__50511;
    wire N__50510;
    wire N__50509;
    wire N__50506;
    wire N__50505;
    wire N__50502;
    wire N__50499;
    wire N__50496;
    wire N__50491;
    wire N__50484;
    wire N__50481;
    wire N__50478;
    wire N__50477;
    wire N__50476;
    wire N__50473;
    wire N__50470;
    wire N__50467;
    wire N__50464;
    wire N__50463;
    wire N__50460;
    wire N__50457;
    wire N__50454;
    wire N__50451;
    wire N__50446;
    wire N__50439;
    wire N__50436;
    wire N__50433;
    wire N__50430;
    wire N__50429;
    wire N__50426;
    wire N__50423;
    wire N__50420;
    wire N__50419;
    wire N__50418;
    wire N__50413;
    wire N__50410;
    wire N__50407;
    wire N__50400;
    wire N__50397;
    wire N__50396;
    wire N__50393;
    wire N__50392;
    wire N__50391;
    wire N__50388;
    wire N__50385;
    wire N__50382;
    wire N__50379;
    wire N__50376;
    wire N__50371;
    wire N__50368;
    wire N__50365;
    wire N__50362;
    wire N__50355;
    wire N__50352;
    wire N__50351;
    wire N__50348;
    wire N__50347;
    wire N__50344;
    wire N__50341;
    wire N__50338;
    wire N__50335;
    wire N__50332;
    wire N__50329;
    wire N__50322;
    wire N__50319;
    wire N__50318;
    wire N__50317;
    wire N__50314;
    wire N__50311;
    wire N__50310;
    wire N__50307;
    wire N__50304;
    wire N__50301;
    wire N__50298;
    wire N__50295;
    wire N__50292;
    wire N__50289;
    wire N__50286;
    wire N__50277;
    wire N__50274;
    wire N__50271;
    wire N__50270;
    wire N__50267;
    wire N__50266;
    wire N__50265;
    wire N__50262;
    wire N__50259;
    wire N__50254;
    wire N__50251;
    wire N__50246;
    wire N__50241;
    wire N__50238;
    wire N__50237;
    wire N__50234;
    wire N__50233;
    wire N__50232;
    wire N__50229;
    wire N__50226;
    wire N__50221;
    wire N__50218;
    wire N__50215;
    wire N__50212;
    wire N__50205;
    wire N__50202;
    wire N__50199;
    wire N__50198;
    wire N__50195;
    wire N__50192;
    wire N__50191;
    wire N__50188;
    wire N__50185;
    wire N__50182;
    wire N__50181;
    wire N__50178;
    wire N__50173;
    wire N__50170;
    wire N__50165;
    wire N__50160;
    wire N__50157;
    wire N__50154;
    wire N__50153;
    wire N__50152;
    wire N__50151;
    wire N__50148;
    wire N__50145;
    wire N__50142;
    wire N__50139;
    wire N__50134;
    wire N__50131;
    wire N__50126;
    wire N__50121;
    wire N__50118;
    wire N__50117;
    wire N__50114;
    wire N__50111;
    wire N__50108;
    wire N__50107;
    wire N__50106;
    wire N__50103;
    wire N__50100;
    wire N__50097;
    wire N__50094;
    wire N__50091;
    wire N__50086;
    wire N__50079;
    wire N__50076;
    wire N__50073;
    wire N__50072;
    wire N__50071;
    wire N__50070;
    wire N__50067;
    wire N__50062;
    wire N__50059;
    wire N__50056;
    wire N__50053;
    wire N__50050;
    wire N__50047;
    wire N__50044;
    wire N__50037;
    wire N__50034;
    wire N__50033;
    wire N__50030;
    wire N__50027;
    wire N__50026;
    wire N__50023;
    wire N__50020;
    wire N__50017;
    wire N__50010;
    wire N__50007;
    wire N__50004;
    wire N__50001;
    wire N__50000;
    wire N__49999;
    wire N__49996;
    wire N__49991;
    wire N__49986;
    wire N__49983;
    wire N__49980;
    wire N__49979;
    wire N__49976;
    wire N__49973;
    wire N__49970;
    wire N__49967;
    wire N__49962;
    wire N__49959;
    wire N__49956;
    wire N__49953;
    wire N__49950;
    wire N__49947;
    wire N__49944;
    wire N__49943;
    wire N__49942;
    wire N__49941;
    wire N__49938;
    wire N__49935;
    wire N__49934;
    wire N__49931;
    wire N__49930;
    wire N__49929;
    wire N__49928;
    wire N__49925;
    wire N__49924;
    wire N__49923;
    wire N__49922;
    wire N__49919;
    wire N__49916;
    wire N__49913;
    wire N__49904;
    wire N__49901;
    wire N__49894;
    wire N__49881;
    wire N__49878;
    wire N__49877;
    wire N__49876;
    wire N__49875;
    wire N__49872;
    wire N__49869;
    wire N__49868;
    wire N__49867;
    wire N__49864;
    wire N__49861;
    wire N__49860;
    wire N__49855;
    wire N__49854;
    wire N__49851;
    wire N__49848;
    wire N__49843;
    wire N__49842;
    wire N__49841;
    wire N__49838;
    wire N__49835;
    wire N__49832;
    wire N__49827;
    wire N__49824;
    wire N__49817;
    wire N__49806;
    wire N__49805;
    wire N__49802;
    wire N__49801;
    wire N__49798;
    wire N__49795;
    wire N__49792;
    wire N__49789;
    wire N__49782;
    wire N__49779;
    wire N__49776;
    wire N__49773;
    wire N__49770;
    wire N__49767;
    wire N__49764;
    wire N__49763;
    wire N__49762;
    wire N__49759;
    wire N__49756;
    wire N__49753;
    wire N__49748;
    wire N__49743;
    wire N__49740;
    wire N__49737;
    wire N__49736;
    wire N__49735;
    wire N__49732;
    wire N__49729;
    wire N__49726;
    wire N__49723;
    wire N__49720;
    wire N__49717;
    wire N__49712;
    wire N__49707;
    wire N__49704;
    wire N__49703;
    wire N__49700;
    wire N__49699;
    wire N__49696;
    wire N__49693;
    wire N__49690;
    wire N__49687;
    wire N__49684;
    wire N__49681;
    wire N__49674;
    wire N__49671;
    wire N__49668;
    wire N__49665;
    wire N__49664;
    wire N__49661;
    wire N__49658;
    wire N__49657;
    wire N__49654;
    wire N__49651;
    wire N__49648;
    wire N__49641;
    wire N__49638;
    wire N__49635;
    wire N__49632;
    wire N__49629;
    wire N__49626;
    wire N__49625;
    wire N__49624;
    wire N__49623;
    wire N__49622;
    wire N__49621;
    wire N__49612;
    wire N__49611;
    wire N__49610;
    wire N__49607;
    wire N__49606;
    wire N__49605;
    wire N__49604;
    wire N__49603;
    wire N__49602;
    wire N__49601;
    wire N__49600;
    wire N__49599;
    wire N__49598;
    wire N__49597;
    wire N__49594;
    wire N__49593;
    wire N__49592;
    wire N__49591;
    wire N__49590;
    wire N__49589;
    wire N__49586;
    wire N__49581;
    wire N__49580;
    wire N__49577;
    wire N__49574;
    wire N__49569;
    wire N__49566;
    wire N__49561;
    wire N__49560;
    wire N__49557;
    wire N__49554;
    wire N__49553;
    wire N__49552;
    wire N__49549;
    wire N__49548;
    wire N__49547;
    wire N__49546;
    wire N__49543;
    wire N__49542;
    wire N__49541;
    wire N__49540;
    wire N__49539;
    wire N__49538;
    wire N__49535;
    wire N__49528;
    wire N__49523;
    wire N__49518;
    wire N__49517;
    wire N__49514;
    wire N__49513;
    wire N__49508;
    wire N__49505;
    wire N__49500;
    wire N__49497;
    wire N__49496;
    wire N__49495;
    wire N__49494;
    wire N__49493;
    wire N__49488;
    wire N__49485;
    wire N__49482;
    wire N__49469;
    wire N__49466;
    wire N__49463;
    wire N__49460;
    wire N__49457;
    wire N__49452;
    wire N__49447;
    wire N__49440;
    wire N__49437;
    wire N__49430;
    wire N__49427;
    wire N__49420;
    wire N__49417;
    wire N__49412;
    wire N__49407;
    wire N__49380;
    wire N__49377;
    wire N__49376;
    wire N__49373;
    wire N__49370;
    wire N__49369;
    wire N__49366;
    wire N__49363;
    wire N__49360;
    wire N__49353;
    wire N__49350;
    wire N__49347;
    wire N__49344;
    wire N__49341;
    wire N__49338;
    wire N__49335;
    wire N__49332;
    wire N__49329;
    wire N__49328;
    wire N__49325;
    wire N__49322;
    wire N__49319;
    wire N__49316;
    wire N__49311;
    wire N__49308;
    wire N__49307;
    wire N__49304;
    wire N__49301;
    wire N__49296;
    wire N__49293;
    wire N__49290;
    wire N__49287;
    wire N__49286;
    wire N__49283;
    wire N__49280;
    wire N__49277;
    wire N__49274;
    wire N__49269;
    wire N__49266;
    wire N__49263;
    wire N__49260;
    wire N__49257;
    wire N__49256;
    wire N__49253;
    wire N__49250;
    wire N__49249;
    wire N__49246;
    wire N__49243;
    wire N__49240;
    wire N__49233;
    wire N__49232;
    wire N__49229;
    wire N__49226;
    wire N__49225;
    wire N__49222;
    wire N__49217;
    wire N__49212;
    wire N__49209;
    wire N__49208;
    wire N__49205;
    wire N__49202;
    wire N__49197;
    wire N__49194;
    wire N__49191;
    wire N__49188;
    wire N__49185;
    wire N__49184;
    wire N__49181;
    wire N__49178;
    wire N__49177;
    wire N__49174;
    wire N__49171;
    wire N__49168;
    wire N__49161;
    wire N__49158;
    wire N__49155;
    wire N__49152;
    wire N__49149;
    wire N__49146;
    wire N__49143;
    wire N__49140;
    wire N__49139;
    wire N__49138;
    wire N__49135;
    wire N__49132;
    wire N__49129;
    wire N__49126;
    wire N__49121;
    wire N__49118;
    wire N__49113;
    wire N__49110;
    wire N__49107;
    wire N__49104;
    wire N__49101;
    wire N__49098;
    wire N__49095;
    wire N__49092;
    wire N__49089;
    wire N__49086;
    wire N__49083;
    wire N__49080;
    wire N__49079;
    wire N__49076;
    wire N__49075;
    wire N__49072;
    wire N__49069;
    wire N__49064;
    wire N__49059;
    wire N__49056;
    wire N__49053;
    wire N__49050;
    wire N__49047;
    wire N__49044;
    wire N__49041;
    wire N__49038;
    wire N__49035;
    wire N__49032;
    wire N__49029;
    wire N__49026;
    wire N__49023;
    wire N__49020;
    wire N__49017;
    wire N__49014;
    wire N__49011;
    wire N__49008;
    wire N__49007;
    wire N__49004;
    wire N__49001;
    wire N__49000;
    wire N__48999;
    wire N__48998;
    wire N__48997;
    wire N__48994;
    wire N__48993;
    wire N__48992;
    wire N__48991;
    wire N__48988;
    wire N__48987;
    wire N__48984;
    wire N__48981;
    wire N__48980;
    wire N__48977;
    wire N__48976;
    wire N__48973;
    wire N__48972;
    wire N__48969;
    wire N__48966;
    wire N__48961;
    wire N__48958;
    wire N__48941;
    wire N__48930;
    wire N__48927;
    wire N__48926;
    wire N__48923;
    wire N__48920;
    wire N__48917;
    wire N__48914;
    wire N__48913;
    wire N__48908;
    wire N__48905;
    wire N__48900;
    wire N__48897;
    wire N__48894;
    wire N__48893;
    wire N__48890;
    wire N__48887;
    wire N__48886;
    wire N__48885;
    wire N__48884;
    wire N__48881;
    wire N__48878;
    wire N__48877;
    wire N__48876;
    wire N__48875;
    wire N__48874;
    wire N__48871;
    wire N__48870;
    wire N__48867;
    wire N__48866;
    wire N__48863;
    wire N__48862;
    wire N__48861;
    wire N__48860;
    wire N__48857;
    wire N__48854;
    wire N__48851;
    wire N__48844;
    wire N__48839;
    wire N__48834;
    wire N__48825;
    wire N__48810;
    wire N__48809;
    wire N__48806;
    wire N__48803;
    wire N__48800;
    wire N__48797;
    wire N__48792;
    wire N__48789;
    wire N__48788;
    wire N__48787;
    wire N__48784;
    wire N__48781;
    wire N__48778;
    wire N__48775;
    wire N__48770;
    wire N__48767;
    wire N__48764;
    wire N__48759;
    wire N__48756;
    wire N__48753;
    wire N__48750;
    wire N__48749;
    wire N__48746;
    wire N__48743;
    wire N__48742;
    wire N__48739;
    wire N__48736;
    wire N__48733;
    wire N__48726;
    wire N__48723;
    wire N__48720;
    wire N__48717;
    wire N__48714;
    wire N__48711;
    wire N__48708;
    wire N__48705;
    wire N__48702;
    wire N__48699;
    wire N__48696;
    wire N__48695;
    wire N__48694;
    wire N__48693;
    wire N__48690;
    wire N__48687;
    wire N__48684;
    wire N__48681;
    wire N__48672;
    wire N__48671;
    wire N__48668;
    wire N__48665;
    wire N__48660;
    wire N__48659;
    wire N__48656;
    wire N__48653;
    wire N__48648;
    wire N__48647;
    wire N__48644;
    wire N__48641;
    wire N__48638;
    wire N__48633;
    wire N__48632;
    wire N__48629;
    wire N__48626;
    wire N__48621;
    wire N__48620;
    wire N__48617;
    wire N__48614;
    wire N__48609;
    wire N__48608;
    wire N__48605;
    wire N__48602;
    wire N__48597;
    wire N__48594;
    wire N__48593;
    wire N__48590;
    wire N__48587;
    wire N__48582;
    wire N__48579;
    wire N__48578;
    wire N__48577;
    wire N__48574;
    wire N__48571;
    wire N__48568;
    wire N__48565;
    wire N__48558;
    wire N__48555;
    wire N__48554;
    wire N__48551;
    wire N__48550;
    wire N__48547;
    wire N__48544;
    wire N__48541;
    wire N__48536;
    wire N__48531;
    wire N__48528;
    wire N__48527;
    wire N__48526;
    wire N__48523;
    wire N__48520;
    wire N__48517;
    wire N__48514;
    wire N__48507;
    wire N__48504;
    wire N__48501;
    wire N__48500;
    wire N__48499;
    wire N__48496;
    wire N__48493;
    wire N__48490;
    wire N__48487;
    wire N__48480;
    wire N__48477;
    wire N__48476;
    wire N__48475;
    wire N__48472;
    wire N__48469;
    wire N__48464;
    wire N__48463;
    wire N__48462;
    wire N__48459;
    wire N__48456;
    wire N__48453;
    wire N__48450;
    wire N__48447;
    wire N__48444;
    wire N__48435;
    wire N__48432;
    wire N__48429;
    wire N__48428;
    wire N__48427;
    wire N__48424;
    wire N__48421;
    wire N__48418;
    wire N__48415;
    wire N__48408;
    wire N__48405;
    wire N__48402;
    wire N__48399;
    wire N__48396;
    wire N__48395;
    wire N__48394;
    wire N__48393;
    wire N__48388;
    wire N__48385;
    wire N__48382;
    wire N__48379;
    wire N__48372;
    wire N__48369;
    wire N__48368;
    wire N__48367;
    wire N__48364;
    wire N__48361;
    wire N__48358;
    wire N__48355;
    wire N__48348;
    wire N__48345;
    wire N__48344;
    wire N__48341;
    wire N__48340;
    wire N__48337;
    wire N__48334;
    wire N__48331;
    wire N__48328;
    wire N__48321;
    wire N__48318;
    wire N__48315;
    wire N__48314;
    wire N__48313;
    wire N__48310;
    wire N__48307;
    wire N__48304;
    wire N__48301;
    wire N__48294;
    wire N__48291;
    wire N__48290;
    wire N__48289;
    wire N__48286;
    wire N__48283;
    wire N__48280;
    wire N__48273;
    wire N__48270;
    wire N__48267;
    wire N__48266;
    wire N__48265;
    wire N__48262;
    wire N__48259;
    wire N__48256;
    wire N__48251;
    wire N__48246;
    wire N__48243;
    wire N__48242;
    wire N__48239;
    wire N__48236;
    wire N__48235;
    wire N__48232;
    wire N__48229;
    wire N__48226;
    wire N__48221;
    wire N__48216;
    wire N__48213;
    wire N__48212;
    wire N__48211;
    wire N__48210;
    wire N__48203;
    wire N__48202;
    wire N__48199;
    wire N__48196;
    wire N__48193;
    wire N__48190;
    wire N__48187;
    wire N__48180;
    wire N__48177;
    wire N__48174;
    wire N__48173;
    wire N__48170;
    wire N__48167;
    wire N__48164;
    wire N__48159;
    wire N__48156;
    wire N__48155;
    wire N__48152;
    wire N__48149;
    wire N__48146;
    wire N__48141;
    wire N__48138;
    wire N__48137;
    wire N__48134;
    wire N__48131;
    wire N__48128;
    wire N__48123;
    wire N__48120;
    wire N__48119;
    wire N__48118;
    wire N__48115;
    wire N__48110;
    wire N__48105;
    wire N__48102;
    wire N__48099;
    wire N__48098;
    wire N__48095;
    wire N__48092;
    wire N__48089;
    wire N__48084;
    wire N__48081;
    wire N__48080;
    wire N__48079;
    wire N__48076;
    wire N__48073;
    wire N__48070;
    wire N__48067;
    wire N__48060;
    wire N__48057;
    wire N__48056;
    wire N__48053;
    wire N__48050;
    wire N__48049;
    wire N__48048;
    wire N__48045;
    wire N__48042;
    wire N__48039;
    wire N__48036;
    wire N__48033;
    wire N__48030;
    wire N__48021;
    wire N__48018;
    wire N__48017;
    wire N__48014;
    wire N__48011;
    wire N__48010;
    wire N__48009;
    wire N__48006;
    wire N__48003;
    wire N__48000;
    wire N__47997;
    wire N__47994;
    wire N__47991;
    wire N__47982;
    wire N__47979;
    wire N__47978;
    wire N__47977;
    wire N__47974;
    wire N__47971;
    wire N__47968;
    wire N__47967;
    wire N__47964;
    wire N__47961;
    wire N__47958;
    wire N__47955;
    wire N__47950;
    wire N__47943;
    wire N__47940;
    wire N__47937;
    wire N__47934;
    wire N__47931;
    wire N__47928;
    wire N__47925;
    wire N__47922;
    wire N__47919;
    wire N__47916;
    wire N__47913;
    wire N__47910;
    wire N__47907;
    wire N__47904;
    wire N__47901;
    wire N__47898;
    wire N__47895;
    wire N__47892;
    wire N__47889;
    wire N__47886;
    wire N__47883;
    wire N__47880;
    wire N__47877;
    wire N__47874;
    wire N__47873;
    wire N__47870;
    wire N__47867;
    wire N__47864;
    wire N__47861;
    wire N__47858;
    wire N__47855;
    wire N__47850;
    wire N__47847;
    wire N__47844;
    wire N__47841;
    wire N__47838;
    wire N__47837;
    wire N__47832;
    wire N__47829;
    wire N__47826;
    wire N__47823;
    wire N__47820;
    wire N__47817;
    wire N__47814;
    wire N__47811;
    wire N__47808;
    wire N__47805;
    wire N__47802;
    wire N__47799;
    wire N__47796;
    wire N__47793;
    wire N__47790;
    wire N__47789;
    wire N__47786;
    wire N__47783;
    wire N__47778;
    wire N__47775;
    wire N__47772;
    wire N__47769;
    wire N__47766;
    wire N__47763;
    wire N__47760;
    wire N__47757;
    wire N__47754;
    wire N__47751;
    wire N__47748;
    wire N__47745;
    wire N__47742;
    wire N__47739;
    wire N__47738;
    wire N__47735;
    wire N__47732;
    wire N__47727;
    wire N__47724;
    wire N__47721;
    wire N__47718;
    wire N__47715;
    wire N__47712;
    wire N__47711;
    wire N__47708;
    wire N__47707;
    wire N__47704;
    wire N__47701;
    wire N__47698;
    wire N__47695;
    wire N__47692;
    wire N__47689;
    wire N__47682;
    wire N__47681;
    wire N__47678;
    wire N__47675;
    wire N__47672;
    wire N__47669;
    wire N__47664;
    wire N__47661;
    wire N__47658;
    wire N__47655;
    wire N__47652;
    wire N__47649;
    wire N__47648;
    wire N__47647;
    wire N__47644;
    wire N__47641;
    wire N__47638;
    wire N__47631;
    wire N__47628;
    wire N__47625;
    wire N__47622;
    wire N__47619;
    wire N__47616;
    wire N__47615;
    wire N__47612;
    wire N__47611;
    wire N__47608;
    wire N__47605;
    wire N__47602;
    wire N__47595;
    wire N__47592;
    wire N__47589;
    wire N__47586;
    wire N__47583;
    wire N__47580;
    wire N__47579;
    wire N__47576;
    wire N__47573;
    wire N__47572;
    wire N__47569;
    wire N__47566;
    wire N__47563;
    wire N__47556;
    wire N__47553;
    wire N__47550;
    wire N__47547;
    wire N__47544;
    wire N__47543;
    wire N__47540;
    wire N__47537;
    wire N__47536;
    wire N__47533;
    wire N__47530;
    wire N__47527;
    wire N__47520;
    wire N__47517;
    wire N__47514;
    wire N__47511;
    wire N__47508;
    wire N__47505;
    wire N__47502;
    wire N__47499;
    wire N__47496;
    wire N__47493;
    wire N__47490;
    wire N__47489;
    wire N__47486;
    wire N__47483;
    wire N__47478;
    wire N__47475;
    wire N__47472;
    wire N__47469;
    wire N__47466;
    wire N__47463;
    wire N__47460;
    wire N__47457;
    wire N__47454;
    wire N__47451;
    wire N__47448;
    wire N__47445;
    wire N__47442;
    wire N__47439;
    wire N__47436;
    wire N__47433;
    wire N__47430;
    wire N__47427;
    wire N__47424;
    wire N__47421;
    wire N__47418;
    wire N__47415;
    wire N__47412;
    wire N__47409;
    wire N__47406;
    wire N__47405;
    wire N__47402;
    wire N__47401;
    wire N__47398;
    wire N__47395;
    wire N__47392;
    wire N__47385;
    wire N__47382;
    wire N__47379;
    wire N__47376;
    wire N__47373;
    wire N__47370;
    wire N__47369;
    wire N__47366;
    wire N__47365;
    wire N__47362;
    wire N__47359;
    wire N__47356;
    wire N__47353;
    wire N__47350;
    wire N__47347;
    wire N__47340;
    wire N__47337;
    wire N__47336;
    wire N__47335;
    wire N__47332;
    wire N__47327;
    wire N__47322;
    wire N__47321;
    wire N__47318;
    wire N__47315;
    wire N__47312;
    wire N__47309;
    wire N__47306;
    wire N__47301;
    wire N__47298;
    wire N__47295;
    wire N__47292;
    wire N__47289;
    wire N__47286;
    wire N__47283;
    wire N__47280;
    wire N__47277;
    wire N__47276;
    wire N__47273;
    wire N__47270;
    wire N__47267;
    wire N__47264;
    wire N__47259;
    wire N__47256;
    wire N__47253;
    wire N__47250;
    wire N__47247;
    wire N__47246;
    wire N__47245;
    wire N__47242;
    wire N__47239;
    wire N__47236;
    wire N__47229;
    wire N__47226;
    wire N__47223;
    wire N__47220;
    wire N__47217;
    wire N__47214;
    wire N__47211;
    wire N__47208;
    wire N__47207;
    wire N__47204;
    wire N__47201;
    wire N__47200;
    wire N__47197;
    wire N__47194;
    wire N__47191;
    wire N__47184;
    wire N__47181;
    wire N__47180;
    wire N__47177;
    wire N__47174;
    wire N__47173;
    wire N__47170;
    wire N__47167;
    wire N__47164;
    wire N__47157;
    wire N__47154;
    wire N__47151;
    wire N__47148;
    wire N__47145;
    wire N__47144;
    wire N__47141;
    wire N__47138;
    wire N__47135;
    wire N__47132;
    wire N__47129;
    wire N__47126;
    wire N__47123;
    wire N__47118;
    wire N__47117;
    wire N__47112;
    wire N__47109;
    wire N__47106;
    wire N__47103;
    wire N__47100;
    wire N__47097;
    wire N__47094;
    wire N__47091;
    wire N__47088;
    wire N__47085;
    wire N__47082;
    wire N__47081;
    wire N__47078;
    wire N__47075;
    wire N__47072;
    wire N__47069;
    wire N__47064;
    wire N__47063;
    wire N__47060;
    wire N__47057;
    wire N__47056;
    wire N__47053;
    wire N__47050;
    wire N__47047;
    wire N__47040;
    wire N__47037;
    wire N__47034;
    wire N__47031;
    wire N__47028;
    wire N__47025;
    wire N__47022;
    wire N__47019;
    wire N__47016;
    wire N__47013;
    wire N__47010;
    wire N__47007;
    wire N__47006;
    wire N__47005;
    wire N__47004;
    wire N__47001;
    wire N__47000;
    wire N__46997;
    wire N__46992;
    wire N__46989;
    wire N__46988;
    wire N__46985;
    wire N__46980;
    wire N__46977;
    wire N__46974;
    wire N__46971;
    wire N__46968;
    wire N__46959;
    wire N__46958;
    wire N__46957;
    wire N__46956;
    wire N__46955;
    wire N__46952;
    wire N__46949;
    wire N__46944;
    wire N__46941;
    wire N__46934;
    wire N__46931;
    wire N__46928;
    wire N__46927;
    wire N__46924;
    wire N__46921;
    wire N__46918;
    wire N__46915;
    wire N__46912;
    wire N__46905;
    wire N__46904;
    wire N__46903;
    wire N__46900;
    wire N__46899;
    wire N__46896;
    wire N__46893;
    wire N__46892;
    wire N__46887;
    wire N__46884;
    wire N__46881;
    wire N__46878;
    wire N__46875;
    wire N__46870;
    wire N__46867;
    wire N__46866;
    wire N__46863;
    wire N__46858;
    wire N__46855;
    wire N__46850;
    wire N__46845;
    wire N__46842;
    wire N__46839;
    wire N__46836;
    wire N__46833;
    wire N__46830;
    wire N__46829;
    wire N__46826;
    wire N__46823;
    wire N__46818;
    wire N__46815;
    wire N__46812;
    wire N__46809;
    wire N__46806;
    wire N__46805;
    wire N__46802;
    wire N__46799;
    wire N__46796;
    wire N__46793;
    wire N__46788;
    wire N__46785;
    wire N__46784;
    wire N__46781;
    wire N__46778;
    wire N__46775;
    wire N__46770;
    wire N__46767;
    wire N__46766;
    wire N__46765;
    wire N__46760;
    wire N__46757;
    wire N__46752;
    wire N__46749;
    wire N__46748;
    wire N__46745;
    wire N__46742;
    wire N__46737;
    wire N__46734;
    wire N__46731;
    wire N__46728;
    wire N__46725;
    wire N__46722;
    wire N__46721;
    wire N__46720;
    wire N__46719;
    wire N__46718;
    wire N__46715;
    wire N__46712;
    wire N__46711;
    wire N__46710;
    wire N__46699;
    wire N__46694;
    wire N__46693;
    wire N__46692;
    wire N__46687;
    wire N__46682;
    wire N__46677;
    wire N__46674;
    wire N__46671;
    wire N__46668;
    wire N__46665;
    wire N__46664;
    wire N__46661;
    wire N__46660;
    wire N__46659;
    wire N__46658;
    wire N__46655;
    wire N__46652;
    wire N__46649;
    wire N__46644;
    wire N__46641;
    wire N__46638;
    wire N__46633;
    wire N__46630;
    wire N__46623;
    wire N__46622;
    wire N__46617;
    wire N__46616;
    wire N__46615;
    wire N__46614;
    wire N__46611;
    wire N__46608;
    wire N__46605;
    wire N__46602;
    wire N__46601;
    wire N__46598;
    wire N__46591;
    wire N__46588;
    wire N__46583;
    wire N__46578;
    wire N__46575;
    wire N__46572;
    wire N__46571;
    wire N__46568;
    wire N__46565;
    wire N__46562;
    wire N__46559;
    wire N__46556;
    wire N__46553;
    wire N__46548;
    wire N__46547;
    wire N__46544;
    wire N__46541;
    wire N__46540;
    wire N__46535;
    wire N__46532;
    wire N__46527;
    wire N__46526;
    wire N__46523;
    wire N__46520;
    wire N__46517;
    wire N__46512;
    wire N__46509;
    wire N__46506;
    wire N__46503;
    wire N__46500;
    wire N__46499;
    wire N__46496;
    wire N__46493;
    wire N__46490;
    wire N__46485;
    wire N__46482;
    wire N__46479;
    wire N__46476;
    wire N__46475;
    wire N__46470;
    wire N__46467;
    wire N__46464;
    wire N__46461;
    wire N__46458;
    wire N__46457;
    wire N__46456;
    wire N__46453;
    wire N__46450;
    wire N__46447;
    wire N__46442;
    wire N__46439;
    wire N__46434;
    wire N__46431;
    wire N__46428;
    wire N__46425;
    wire N__46424;
    wire N__46421;
    wire N__46418;
    wire N__46417;
    wire N__46412;
    wire N__46409;
    wire N__46406;
    wire N__46401;
    wire N__46400;
    wire N__46397;
    wire N__46396;
    wire N__46395;
    wire N__46394;
    wire N__46393;
    wire N__46390;
    wire N__46387;
    wire N__46380;
    wire N__46377;
    wire N__46372;
    wire N__46369;
    wire N__46366;
    wire N__46361;
    wire N__46356;
    wire N__46353;
    wire N__46350;
    wire N__46347;
    wire N__46344;
    wire N__46341;
    wire N__46340;
    wire N__46337;
    wire N__46334;
    wire N__46333;
    wire N__46332;
    wire N__46327;
    wire N__46322;
    wire N__46319;
    wire N__46316;
    wire N__46313;
    wire N__46308;
    wire N__46307;
    wire N__46306;
    wire N__46303;
    wire N__46300;
    wire N__46297;
    wire N__46294;
    wire N__46291;
    wire N__46288;
    wire N__46281;
    wire N__46278;
    wire N__46277;
    wire N__46274;
    wire N__46271;
    wire N__46270;
    wire N__46269;
    wire N__46266;
    wire N__46263;
    wire N__46260;
    wire N__46257;
    wire N__46254;
    wire N__46251;
    wire N__46248;
    wire N__46239;
    wire N__46236;
    wire N__46233;
    wire N__46230;
    wire N__46227;
    wire N__46224;
    wire N__46221;
    wire N__46218;
    wire N__46215;
    wire N__46212;
    wire N__46209;
    wire N__46208;
    wire N__46205;
    wire N__46202;
    wire N__46197;
    wire N__46196;
    wire N__46191;
    wire N__46188;
    wire N__46185;
    wire N__46184;
    wire N__46179;
    wire N__46176;
    wire N__46173;
    wire N__46170;
    wire N__46167;
    wire N__46164;
    wire N__46161;
    wire N__46158;
    wire N__46155;
    wire N__46152;
    wire N__46149;
    wire N__46146;
    wire N__46143;
    wire N__46142;
    wire N__46139;
    wire N__46136;
    wire N__46131;
    wire N__46128;
    wire N__46125;
    wire N__46122;
    wire N__46119;
    wire N__46116;
    wire N__46113;
    wire N__46110;
    wire N__46107;
    wire N__46104;
    wire N__46101;
    wire N__46100;
    wire N__46097;
    wire N__46096;
    wire N__46093;
    wire N__46090;
    wire N__46087;
    wire N__46080;
    wire N__46077;
    wire N__46074;
    wire N__46071;
    wire N__46068;
    wire N__46065;
    wire N__46064;
    wire N__46061;
    wire N__46058;
    wire N__46055;
    wire N__46050;
    wire N__46047;
    wire N__46044;
    wire N__46041;
    wire N__46038;
    wire N__46037;
    wire N__46036;
    wire N__46033;
    wire N__46028;
    wire N__46023;
    wire N__46020;
    wire N__46017;
    wire N__46014;
    wire N__46013;
    wire N__46012;
    wire N__46009;
    wire N__46008;
    wire N__46005;
    wire N__46004;
    wire N__46003;
    wire N__46002;
    wire N__45999;
    wire N__45996;
    wire N__45993;
    wire N__45984;
    wire N__45975;
    wire N__45972;
    wire N__45969;
    wire N__45968;
    wire N__45965;
    wire N__45962;
    wire N__45957;
    wire N__45954;
    wire N__45951;
    wire N__45948;
    wire N__45945;
    wire N__45942;
    wire N__45939;
    wire N__45936;
    wire N__45933;
    wire N__45930;
    wire N__45927;
    wire N__45924;
    wire N__45923;
    wire N__45920;
    wire N__45917;
    wire N__45912;
    wire N__45909;
    wire N__45906;
    wire N__45903;
    wire N__45900;
    wire N__45899;
    wire N__45896;
    wire N__45893;
    wire N__45888;
    wire N__45885;
    wire N__45882;
    wire N__45879;
    wire N__45876;
    wire N__45875;
    wire N__45872;
    wire N__45869;
    wire N__45864;
    wire N__45861;
    wire N__45858;
    wire N__45855;
    wire N__45854;
    wire N__45851;
    wire N__45850;
    wire N__45847;
    wire N__45844;
    wire N__45841;
    wire N__45834;
    wire N__45831;
    wire N__45828;
    wire N__45825;
    wire N__45822;
    wire N__45819;
    wire N__45816;
    wire N__45813;
    wire N__45810;
    wire N__45807;
    wire N__45804;
    wire N__45801;
    wire N__45800;
    wire N__45799;
    wire N__45796;
    wire N__45793;
    wire N__45790;
    wire N__45787;
    wire N__45784;
    wire N__45781;
    wire N__45776;
    wire N__45771;
    wire N__45768;
    wire N__45765;
    wire N__45762;
    wire N__45759;
    wire N__45758;
    wire N__45757;
    wire N__45754;
    wire N__45751;
    wire N__45748;
    wire N__45743;
    wire N__45740;
    wire N__45737;
    wire N__45732;
    wire N__45729;
    wire N__45726;
    wire N__45723;
    wire N__45720;
    wire N__45717;
    wire N__45714;
    wire N__45711;
    wire N__45708;
    wire N__45705;
    wire N__45702;
    wire N__45701;
    wire N__45698;
    wire N__45695;
    wire N__45692;
    wire N__45689;
    wire N__45684;
    wire N__45681;
    wire N__45678;
    wire N__45677;
    wire N__45674;
    wire N__45671;
    wire N__45670;
    wire N__45667;
    wire N__45664;
    wire N__45661;
    wire N__45654;
    wire N__45651;
    wire N__45648;
    wire N__45645;
    wire N__45642;
    wire N__45639;
    wire N__45636;
    wire N__45633;
    wire N__45630;
    wire N__45627;
    wire N__45624;
    wire N__45621;
    wire N__45618;
    wire N__45617;
    wire N__45616;
    wire N__45615;
    wire N__45614;
    wire N__45613;
    wire N__45610;
    wire N__45609;
    wire N__45608;
    wire N__45605;
    wire N__45604;
    wire N__45603;
    wire N__45602;
    wire N__45599;
    wire N__45598;
    wire N__45597;
    wire N__45594;
    wire N__45591;
    wire N__45588;
    wire N__45587;
    wire N__45586;
    wire N__45583;
    wire N__45578;
    wire N__45575;
    wire N__45564;
    wire N__45559;
    wire N__45550;
    wire N__45537;
    wire N__45534;
    wire N__45533;
    wire N__45530;
    wire N__45527;
    wire N__45526;
    wire N__45523;
    wire N__45520;
    wire N__45517;
    wire N__45510;
    wire N__45507;
    wire N__45506;
    wire N__45503;
    wire N__45502;
    wire N__45501;
    wire N__45500;
    wire N__45499;
    wire N__45496;
    wire N__45493;
    wire N__45490;
    wire N__45487;
    wire N__45486;
    wire N__45485;
    wire N__45484;
    wire N__45481;
    wire N__45480;
    wire N__45477;
    wire N__45476;
    wire N__45473;
    wire N__45468;
    wire N__45465;
    wire N__45462;
    wire N__45461;
    wire N__45458;
    wire N__45457;
    wire N__45456;
    wire N__45455;
    wire N__45454;
    wire N__45451;
    wire N__45448;
    wire N__45445;
    wire N__45440;
    wire N__45433;
    wire N__45422;
    wire N__45417;
    wire N__45410;
    wire N__45399;
    wire N__45396;
    wire N__45393;
    wire N__45390;
    wire N__45389;
    wire N__45386;
    wire N__45383;
    wire N__45380;
    wire N__45377;
    wire N__45372;
    wire N__45371;
    wire N__45368;
    wire N__45365;
    wire N__45364;
    wire N__45361;
    wire N__45358;
    wire N__45355;
    wire N__45348;
    wire N__45345;
    wire N__45342;
    wire N__45341;
    wire N__45338;
    wire N__45335;
    wire N__45332;
    wire N__45329;
    wire N__45324;
    wire N__45321;
    wire N__45318;
    wire N__45315;
    wire N__45314;
    wire N__45311;
    wire N__45310;
    wire N__45307;
    wire N__45304;
    wire N__45301;
    wire N__45294;
    wire N__45291;
    wire N__45288;
    wire N__45285;
    wire N__45282;
    wire N__45279;
    wire N__45278;
    wire N__45277;
    wire N__45274;
    wire N__45269;
    wire N__45264;
    wire N__45261;
    wire N__45258;
    wire N__45255;
    wire N__45252;
    wire N__45249;
    wire N__45246;
    wire N__45245;
    wire N__45242;
    wire N__45239;
    wire N__45236;
    wire N__45235;
    wire N__45232;
    wire N__45229;
    wire N__45226;
    wire N__45219;
    wire N__45216;
    wire N__45213;
    wire N__45210;
    wire N__45209;
    wire N__45206;
    wire N__45203;
    wire N__45200;
    wire N__45197;
    wire N__45196;
    wire N__45193;
    wire N__45190;
    wire N__45187;
    wire N__45180;
    wire N__45177;
    wire N__45174;
    wire N__45171;
    wire N__45168;
    wire N__45167;
    wire N__45164;
    wire N__45161;
    wire N__45156;
    wire N__45155;
    wire N__45152;
    wire N__45149;
    wire N__45146;
    wire N__45141;
    wire N__45138;
    wire N__45135;
    wire N__45132;
    wire N__45129;
    wire N__45126;
    wire N__45123;
    wire N__45120;
    wire N__45117;
    wire N__45114;
    wire N__45111;
    wire N__45108;
    wire N__45105;
    wire N__45102;
    wire N__45099;
    wire N__45096;
    wire N__45093;
    wire N__45090;
    wire N__45087;
    wire N__45084;
    wire N__45081;
    wire N__45078;
    wire N__45077;
    wire N__45072;
    wire N__45069;
    wire N__45066;
    wire N__45063;
    wire N__45060;
    wire N__45059;
    wire N__45054;
    wire N__45051;
    wire N__45050;
    wire N__45049;
    wire N__45046;
    wire N__45039;
    wire N__45036;
    wire N__45033;
    wire N__45030;
    wire N__45027;
    wire N__45024;
    wire N__45021;
    wire N__45020;
    wire N__45015;
    wire N__45012;
    wire N__45009;
    wire N__45006;
    wire N__45005;
    wire N__45000;
    wire N__44997;
    wire N__44994;
    wire N__44991;
    wire N__44988;
    wire N__44985;
    wire N__44982;
    wire N__44979;
    wire N__44976;
    wire N__44973;
    wire N__44970;
    wire N__44967;
    wire N__44964;
    wire N__44961;
    wire N__44958;
    wire N__44955;
    wire N__44954;
    wire N__44951;
    wire N__44948;
    wire N__44943;
    wire N__44940;
    wire N__44937;
    wire N__44934;
    wire N__44931;
    wire N__44928;
    wire N__44925;
    wire N__44922;
    wire N__44919;
    wire N__44916;
    wire N__44913;
    wire N__44910;
    wire N__44907;
    wire N__44904;
    wire N__44901;
    wire N__44898;
    wire N__44895;
    wire N__44892;
    wire N__44889;
    wire N__44886;
    wire N__44883;
    wire N__44880;
    wire N__44879;
    wire N__44878;
    wire N__44875;
    wire N__44870;
    wire N__44865;
    wire N__44862;
    wire N__44859;
    wire N__44856;
    wire N__44853;
    wire N__44850;
    wire N__44847;
    wire N__44844;
    wire N__44841;
    wire N__44838;
    wire N__44835;
    wire N__44832;
    wire N__44829;
    wire N__44826;
    wire N__44823;
    wire N__44820;
    wire N__44819;
    wire N__44816;
    wire N__44813;
    wire N__44808;
    wire N__44807;
    wire N__44802;
    wire N__44799;
    wire N__44796;
    wire N__44793;
    wire N__44790;
    wire N__44789;
    wire N__44788;
    wire N__44785;
    wire N__44782;
    wire N__44779;
    wire N__44774;
    wire N__44769;
    wire N__44766;
    wire N__44765;
    wire N__44760;
    wire N__44757;
    wire N__44754;
    wire N__44751;
    wire N__44748;
    wire N__44747;
    wire N__44744;
    wire N__44741;
    wire N__44738;
    wire N__44733;
    wire N__44732;
    wire N__44729;
    wire N__44726;
    wire N__44721;
    wire N__44718;
    wire N__44715;
    wire N__44712;
    wire N__44711;
    wire N__44708;
    wire N__44705;
    wire N__44700;
    wire N__44697;
    wire N__44696;
    wire N__44691;
    wire N__44688;
    wire N__44685;
    wire N__44682;
    wire N__44679;
    wire N__44678;
    wire N__44677;
    wire N__44674;
    wire N__44669;
    wire N__44664;
    wire N__44661;
    wire N__44658;
    wire N__44655;
    wire N__44652;
    wire N__44649;
    wire N__44646;
    wire N__44643;
    wire N__44640;
    wire N__44639;
    wire N__44636;
    wire N__44633;
    wire N__44628;
    wire N__44625;
    wire N__44622;
    wire N__44619;
    wire N__44618;
    wire N__44613;
    wire N__44610;
    wire N__44607;
    wire N__44604;
    wire N__44601;
    wire N__44598;
    wire N__44595;
    wire N__44592;
    wire N__44591;
    wire N__44588;
    wire N__44585;
    wire N__44580;
    wire N__44577;
    wire N__44574;
    wire N__44571;
    wire N__44570;
    wire N__44567;
    wire N__44564;
    wire N__44559;
    wire N__44556;
    wire N__44553;
    wire N__44550;
    wire N__44547;
    wire N__44544;
    wire N__44543;
    wire N__44540;
    wire N__44537;
    wire N__44532;
    wire N__44529;
    wire N__44526;
    wire N__44523;
    wire N__44520;
    wire N__44517;
    wire N__44514;
    wire N__44511;
    wire N__44508;
    wire N__44505;
    wire N__44502;
    wire N__44501;
    wire N__44498;
    wire N__44495;
    wire N__44490;
    wire N__44487;
    wire N__44484;
    wire N__44483;
    wire N__44478;
    wire N__44475;
    wire N__44472;
    wire N__44469;
    wire N__44466;
    wire N__44463;
    wire N__44460;
    wire N__44457;
    wire N__44454;
    wire N__44451;
    wire N__44450;
    wire N__44447;
    wire N__44444;
    wire N__44439;
    wire N__44436;
    wire N__44433;
    wire N__44430;
    wire N__44427;
    wire N__44424;
    wire N__44421;
    wire N__44418;
    wire N__44415;
    wire N__44412;
    wire N__44409;
    wire N__44406;
    wire N__44403;
    wire N__44400;
    wire N__44397;
    wire N__44394;
    wire N__44391;
    wire N__44388;
    wire N__44385;
    wire N__44382;
    wire N__44379;
    wire N__44376;
    wire N__44373;
    wire N__44370;
    wire N__44367;
    wire N__44364;
    wire N__44361;
    wire N__44358;
    wire N__44355;
    wire N__44352;
    wire N__44349;
    wire N__44346;
    wire N__44343;
    wire N__44340;
    wire N__44337;
    wire N__44334;
    wire N__44333;
    wire N__44330;
    wire N__44327;
    wire N__44322;
    wire N__44319;
    wire N__44316;
    wire N__44313;
    wire N__44310;
    wire N__44309;
    wire N__44306;
    wire N__44303;
    wire N__44300;
    wire N__44297;
    wire N__44294;
    wire N__44291;
    wire N__44288;
    wire N__44283;
    wire N__44280;
    wire N__44277;
    wire N__44274;
    wire N__44271;
    wire N__44270;
    wire N__44267;
    wire N__44264;
    wire N__44261;
    wire N__44258;
    wire N__44255;
    wire N__44252;
    wire N__44247;
    wire N__44244;
    wire N__44241;
    wire N__44238;
    wire N__44235;
    wire N__44232;
    wire N__44231;
    wire N__44228;
    wire N__44225;
    wire N__44222;
    wire N__44219;
    wire N__44214;
    wire N__44211;
    wire N__44208;
    wire N__44205;
    wire N__44202;
    wire N__44201;
    wire N__44198;
    wire N__44195;
    wire N__44192;
    wire N__44189;
    wire N__44186;
    wire N__44181;
    wire N__44178;
    wire N__44175;
    wire N__44172;
    wire N__44169;
    wire N__44166;
    wire N__44163;
    wire N__44160;
    wire N__44157;
    wire N__44154;
    wire N__44151;
    wire N__44150;
    wire N__44147;
    wire N__44144;
    wire N__44139;
    wire N__44136;
    wire N__44133;
    wire N__44130;
    wire N__44127;
    wire N__44124;
    wire N__44121;
    wire N__44120;
    wire N__44117;
    wire N__44114;
    wire N__44111;
    wire N__44108;
    wire N__44105;
    wire N__44100;
    wire N__44097;
    wire N__44094;
    wire N__44093;
    wire N__44092;
    wire N__44091;
    wire N__44090;
    wire N__44089;
    wire N__44086;
    wire N__44083;
    wire N__44076;
    wire N__44073;
    wire N__44064;
    wire N__44063;
    wire N__44060;
    wire N__44057;
    wire N__44054;
    wire N__44051;
    wire N__44046;
    wire N__44043;
    wire N__44040;
    wire N__44037;
    wire N__44034;
    wire N__44031;
    wire N__44028;
    wire N__44025;
    wire N__44022;
    wire N__44019;
    wire N__44016;
    wire N__44013;
    wire N__44010;
    wire N__44007;
    wire N__44004;
    wire N__44001;
    wire N__43998;
    wire N__43995;
    wire N__43992;
    wire N__43991;
    wire N__43988;
    wire N__43985;
    wire N__43980;
    wire N__43977;
    wire N__43974;
    wire N__43971;
    wire N__43968;
    wire N__43965;
    wire N__43962;
    wire N__43959;
    wire N__43958;
    wire N__43955;
    wire N__43952;
    wire N__43947;
    wire N__43944;
    wire N__43941;
    wire N__43938;
    wire N__43935;
    wire N__43932;
    wire N__43929;
    wire N__43926;
    wire N__43923;
    wire N__43920;
    wire N__43917;
    wire N__43916;
    wire N__43913;
    wire N__43910;
    wire N__43909;
    wire N__43906;
    wire N__43903;
    wire N__43900;
    wire N__43897;
    wire N__43894;
    wire N__43887;
    wire N__43884;
    wire N__43881;
    wire N__43878;
    wire N__43875;
    wire N__43874;
    wire N__43871;
    wire N__43868;
    wire N__43863;
    wire N__43860;
    wire N__43857;
    wire N__43854;
    wire N__43851;
    wire N__43848;
    wire N__43845;
    wire N__43842;
    wire N__43839;
    wire N__43838;
    wire N__43837;
    wire N__43834;
    wire N__43831;
    wire N__43828;
    wire N__43825;
    wire N__43822;
    wire N__43817;
    wire N__43814;
    wire N__43809;
    wire N__43808;
    wire N__43805;
    wire N__43802;
    wire N__43801;
    wire N__43798;
    wire N__43795;
    wire N__43792;
    wire N__43787;
    wire N__43784;
    wire N__43779;
    wire N__43776;
    wire N__43773;
    wire N__43770;
    wire N__43767;
    wire N__43764;
    wire N__43761;
    wire N__43758;
    wire N__43755;
    wire N__43752;
    wire N__43749;
    wire N__43748;
    wire N__43745;
    wire N__43742;
    wire N__43739;
    wire N__43736;
    wire N__43735;
    wire N__43730;
    wire N__43727;
    wire N__43724;
    wire N__43719;
    wire N__43716;
    wire N__43713;
    wire N__43710;
    wire N__43707;
    wire N__43704;
    wire N__43701;
    wire N__43698;
    wire N__43695;
    wire N__43692;
    wire N__43689;
    wire N__43688;
    wire N__43687;
    wire N__43684;
    wire N__43681;
    wire N__43678;
    wire N__43671;
    wire N__43668;
    wire N__43665;
    wire N__43662;
    wire N__43659;
    wire N__43656;
    wire N__43655;
    wire N__43652;
    wire N__43649;
    wire N__43648;
    wire N__43645;
    wire N__43642;
    wire N__43639;
    wire N__43634;
    wire N__43631;
    wire N__43626;
    wire N__43623;
    wire N__43620;
    wire N__43619;
    wire N__43616;
    wire N__43613;
    wire N__43610;
    wire N__43607;
    wire N__43604;
    wire N__43599;
    wire N__43596;
    wire N__43593;
    wire N__43592;
    wire N__43589;
    wire N__43586;
    wire N__43585;
    wire N__43582;
    wire N__43579;
    wire N__43576;
    wire N__43571;
    wire N__43566;
    wire N__43563;
    wire N__43560;
    wire N__43557;
    wire N__43554;
    wire N__43553;
    wire N__43550;
    wire N__43547;
    wire N__43544;
    wire N__43539;
    wire N__43536;
    wire N__43533;
    wire N__43530;
    wire N__43527;
    wire N__43524;
    wire N__43521;
    wire N__43518;
    wire N__43515;
    wire N__43512;
    wire N__43509;
    wire N__43506;
    wire N__43503;
    wire N__43500;
    wire N__43497;
    wire N__43494;
    wire N__43491;
    wire N__43488;
    wire N__43487;
    wire N__43484;
    wire N__43483;
    wire N__43480;
    wire N__43477;
    wire N__43474;
    wire N__43467;
    wire N__43464;
    wire N__43461;
    wire N__43458;
    wire N__43455;
    wire N__43452;
    wire N__43449;
    wire N__43448;
    wire N__43445;
    wire N__43442;
    wire N__43437;
    wire N__43434;
    wire N__43431;
    wire N__43428;
    wire N__43425;
    wire N__43422;
    wire N__43419;
    wire N__43418;
    wire N__43415;
    wire N__43412;
    wire N__43407;
    wire N__43404;
    wire N__43401;
    wire N__43398;
    wire N__43395;
    wire N__43392;
    wire N__43391;
    wire N__43390;
    wire N__43387;
    wire N__43384;
    wire N__43381;
    wire N__43376;
    wire N__43373;
    wire N__43368;
    wire N__43365;
    wire N__43362;
    wire N__43359;
    wire N__43356;
    wire N__43353;
    wire N__43350;
    wire N__43347;
    wire N__43344;
    wire N__43341;
    wire N__43338;
    wire N__43335;
    wire N__43332;
    wire N__43329;
    wire N__43326;
    wire N__43323;
    wire N__43320;
    wire N__43317;
    wire N__43314;
    wire N__43311;
    wire N__43310;
    wire N__43307;
    wire N__43304;
    wire N__43303;
    wire N__43300;
    wire N__43297;
    wire N__43294;
    wire N__43287;
    wire N__43284;
    wire N__43281;
    wire N__43278;
    wire N__43275;
    wire N__43272;
    wire N__43271;
    wire N__43268;
    wire N__43265;
    wire N__43262;
    wire N__43259;
    wire N__43254;
    wire N__43251;
    wire N__43248;
    wire N__43245;
    wire N__43242;
    wire N__43239;
    wire N__43236;
    wire N__43233;
    wire N__43230;
    wire N__43227;
    wire N__43224;
    wire N__43221;
    wire N__43218;
    wire N__43215;
    wire N__43212;
    wire N__43209;
    wire N__43206;
    wire N__43203;
    wire N__43200;
    wire N__43197;
    wire N__43194;
    wire N__43193;
    wire N__43190;
    wire N__43187;
    wire N__43186;
    wire N__43183;
    wire N__43180;
    wire N__43177;
    wire N__43170;
    wire N__43169;
    wire N__43166;
    wire N__43163;
    wire N__43162;
    wire N__43159;
    wire N__43156;
    wire N__43153;
    wire N__43146;
    wire N__43143;
    wire N__43142;
    wire N__43139;
    wire N__43136;
    wire N__43135;
    wire N__43132;
    wire N__43129;
    wire N__43126;
    wire N__43119;
    wire N__43116;
    wire N__43113;
    wire N__43112;
    wire N__43111;
    wire N__43108;
    wire N__43105;
    wire N__43102;
    wire N__43099;
    wire N__43096;
    wire N__43093;
    wire N__43086;
    wire N__43083;
    wire N__43082;
    wire N__43079;
    wire N__43076;
    wire N__43075;
    wire N__43072;
    wire N__43069;
    wire N__43066;
    wire N__43059;
    wire N__43058;
    wire N__43057;
    wire N__43054;
    wire N__43051;
    wire N__43046;
    wire N__43043;
    wire N__43040;
    wire N__43035;
    wire N__43032;
    wire N__43031;
    wire N__43028;
    wire N__43027;
    wire N__43024;
    wire N__43021;
    wire N__43018;
    wire N__43015;
    wire N__43010;
    wire N__43005;
    wire N__43002;
    wire N__42999;
    wire N__42996;
    wire N__42993;
    wire N__42990;
    wire N__42987;
    wire N__42984;
    wire N__42981;
    wire N__42980;
    wire N__42979;
    wire N__42972;
    wire N__42969;
    wire N__42966;
    wire N__42965;
    wire N__42964;
    wire N__42961;
    wire N__42958;
    wire N__42955;
    wire N__42952;
    wire N__42947;
    wire N__42942;
    wire N__42939;
    wire N__42936;
    wire N__42933;
    wire N__42930;
    wire N__42929;
    wire N__42926;
    wire N__42923;
    wire N__42920;
    wire N__42917;
    wire N__42914;
    wire N__42911;
    wire N__42906;
    wire N__42903;
    wire N__42900;
    wire N__42897;
    wire N__42896;
    wire N__42891;
    wire N__42888;
    wire N__42885;
    wire N__42882;
    wire N__42879;
    wire N__42878;
    wire N__42875;
    wire N__42872;
    wire N__42869;
    wire N__42866;
    wire N__42861;
    wire N__42858;
    wire N__42855;
    wire N__42852;
    wire N__42849;
    wire N__42848;
    wire N__42845;
    wire N__42842;
    wire N__42841;
    wire N__42838;
    wire N__42835;
    wire N__42832;
    wire N__42825;
    wire N__42822;
    wire N__42819;
    wire N__42816;
    wire N__42815;
    wire N__42810;
    wire N__42807;
    wire N__42804;
    wire N__42803;
    wire N__42800;
    wire N__42797;
    wire N__42794;
    wire N__42789;
    wire N__42786;
    wire N__42783;
    wire N__42780;
    wire N__42779;
    wire N__42774;
    wire N__42771;
    wire N__42768;
    wire N__42765;
    wire N__42762;
    wire N__42759;
    wire N__42756;
    wire N__42753;
    wire N__42750;
    wire N__42747;
    wire N__42744;
    wire N__42741;
    wire N__42738;
    wire N__42735;
    wire N__42732;
    wire N__42729;
    wire N__42726;
    wire N__42723;
    wire N__42720;
    wire N__42717;
    wire N__42714;
    wire N__42711;
    wire N__42708;
    wire N__42705;
    wire N__42704;
    wire N__42703;
    wire N__42696;
    wire N__42693;
    wire N__42690;
    wire N__42687;
    wire N__42684;
    wire N__42681;
    wire N__42678;
    wire N__42675;
    wire N__42672;
    wire N__42669;
    wire N__42666;
    wire N__42663;
    wire N__42660;
    wire N__42657;
    wire N__42654;
    wire N__42651;
    wire N__42648;
    wire N__42645;
    wire N__42642;
    wire N__42639;
    wire N__42636;
    wire N__42633;
    wire N__42630;
    wire N__42627;
    wire N__42624;
    wire N__42621;
    wire N__42618;
    wire N__42615;
    wire N__42612;
    wire N__42609;
    wire N__42606;
    wire N__42603;
    wire N__42600;
    wire N__42597;
    wire N__42594;
    wire N__42591;
    wire N__42588;
    wire N__42585;
    wire N__42582;
    wire N__42579;
    wire N__42576;
    wire N__42573;
    wire N__42570;
    wire N__42567;
    wire N__42564;
    wire N__42561;
    wire N__42558;
    wire N__42555;
    wire N__42552;
    wire N__42549;
    wire N__42546;
    wire N__42543;
    wire N__42540;
    wire N__42537;
    wire N__42534;
    wire N__42531;
    wire N__42528;
    wire N__42525;
    wire N__42522;
    wire N__42519;
    wire N__42516;
    wire N__42513;
    wire N__42510;
    wire N__42507;
    wire N__42504;
    wire N__42501;
    wire N__42498;
    wire N__42495;
    wire N__42492;
    wire N__42489;
    wire N__42486;
    wire N__42483;
    wire N__42480;
    wire N__42477;
    wire N__42474;
    wire N__42471;
    wire N__42468;
    wire N__42465;
    wire N__42462;
    wire N__42459;
    wire N__42456;
    wire N__42453;
    wire N__42450;
    wire N__42447;
    wire N__42444;
    wire N__42441;
    wire N__42438;
    wire N__42435;
    wire N__42432;
    wire N__42429;
    wire N__42428;
    wire N__42427;
    wire N__42424;
    wire N__42421;
    wire N__42418;
    wire N__42415;
    wire N__42410;
    wire N__42407;
    wire N__42404;
    wire N__42399;
    wire N__42396;
    wire N__42393;
    wire N__42390;
    wire N__42387;
    wire N__42384;
    wire N__42381;
    wire N__42378;
    wire N__42377;
    wire N__42374;
    wire N__42371;
    wire N__42366;
    wire N__42363;
    wire N__42360;
    wire N__42357;
    wire N__42354;
    wire N__42351;
    wire N__42348;
    wire N__42347;
    wire N__42344;
    wire N__42341;
    wire N__42340;
    wire N__42337;
    wire N__42334;
    wire N__42331;
    wire N__42326;
    wire N__42323;
    wire N__42318;
    wire N__42317;
    wire N__42316;
    wire N__42313;
    wire N__42310;
    wire N__42307;
    wire N__42304;
    wire N__42301;
    wire N__42298;
    wire N__42295;
    wire N__42292;
    wire N__42289;
    wire N__42282;
    wire N__42281;
    wire N__42278;
    wire N__42275;
    wire N__42272;
    wire N__42269;
    wire N__42264;
    wire N__42263;
    wire N__42260;
    wire N__42257;
    wire N__42256;
    wire N__42253;
    wire N__42250;
    wire N__42247;
    wire N__42244;
    wire N__42241;
    wire N__42238;
    wire N__42231;
    wire N__42228;
    wire N__42225;
    wire N__42222;
    wire N__42221;
    wire N__42220;
    wire N__42219;
    wire N__42212;
    wire N__42209;
    wire N__42204;
    wire N__42201;
    wire N__42198;
    wire N__42195;
    wire N__42194;
    wire N__42193;
    wire N__42190;
    wire N__42189;
    wire N__42188;
    wire N__42185;
    wire N__42182;
    wire N__42175;
    wire N__42168;
    wire N__42165;
    wire N__42162;
    wire N__42159;
    wire N__42156;
    wire N__42155;
    wire N__42152;
    wire N__42151;
    wire N__42148;
    wire N__42145;
    wire N__42142;
    wire N__42135;
    wire N__42132;
    wire N__42129;
    wire N__42126;
    wire N__42125;
    wire N__42122;
    wire N__42119;
    wire N__42118;
    wire N__42115;
    wire N__42112;
    wire N__42109;
    wire N__42106;
    wire N__42099;
    wire N__42096;
    wire N__42093;
    wire N__42090;
    wire N__42087;
    wire N__42084;
    wire N__42081;
    wire N__42078;
    wire N__42075;
    wire N__42074;
    wire N__42073;
    wire N__42070;
    wire N__42067;
    wire N__42064;
    wire N__42063;
    wire N__42060;
    wire N__42057;
    wire N__42054;
    wire N__42051;
    wire N__42048;
    wire N__42045;
    wire N__42036;
    wire N__42033;
    wire N__42030;
    wire N__42027;
    wire N__42024;
    wire N__42021;
    wire N__42020;
    wire N__42019;
    wire N__42016;
    wire N__42013;
    wire N__42010;
    wire N__42007;
    wire N__42004;
    wire N__42003;
    wire N__42000;
    wire N__41995;
    wire N__41992;
    wire N__41985;
    wire N__41982;
    wire N__41979;
    wire N__41976;
    wire N__41973;
    wire N__41970;
    wire N__41967;
    wire N__41964;
    wire N__41961;
    wire N__41958;
    wire N__41955;
    wire N__41954;
    wire N__41951;
    wire N__41950;
    wire N__41949;
    wire N__41946;
    wire N__41943;
    wire N__41940;
    wire N__41937;
    wire N__41928;
    wire N__41925;
    wire N__41922;
    wire N__41919;
    wire N__41918;
    wire N__41917;
    wire N__41914;
    wire N__41909;
    wire N__41904;
    wire N__41901;
    wire N__41898;
    wire N__41895;
    wire N__41892;
    wire N__41889;
    wire N__41886;
    wire N__41883;
    wire N__41880;
    wire N__41877;
    wire N__41874;
    wire N__41871;
    wire N__41868;
    wire N__41865;
    wire N__41862;
    wire N__41859;
    wire N__41856;
    wire N__41853;
    wire N__41850;
    wire N__41847;
    wire N__41846;
    wire N__41843;
    wire N__41840;
    wire N__41835;
    wire N__41832;
    wire N__41829;
    wire N__41828;
    wire N__41825;
    wire N__41822;
    wire N__41821;
    wire N__41818;
    wire N__41817;
    wire N__41814;
    wire N__41811;
    wire N__41808;
    wire N__41805;
    wire N__41796;
    wire N__41793;
    wire N__41790;
    wire N__41787;
    wire N__41786;
    wire N__41785;
    wire N__41784;
    wire N__41781;
    wire N__41778;
    wire N__41775;
    wire N__41772;
    wire N__41767;
    wire N__41760;
    wire N__41757;
    wire N__41754;
    wire N__41751;
    wire N__41748;
    wire N__41745;
    wire N__41744;
    wire N__41741;
    wire N__41738;
    wire N__41735;
    wire N__41732;
    wire N__41729;
    wire N__41726;
    wire N__41725;
    wire N__41720;
    wire N__41717;
    wire N__41712;
    wire N__41709;
    wire N__41706;
    wire N__41703;
    wire N__41702;
    wire N__41699;
    wire N__41696;
    wire N__41693;
    wire N__41690;
    wire N__41687;
    wire N__41684;
    wire N__41683;
    wire N__41680;
    wire N__41677;
    wire N__41674;
    wire N__41667;
    wire N__41666;
    wire N__41665;
    wire N__41662;
    wire N__41657;
    wire N__41654;
    wire N__41649;
    wire N__41646;
    wire N__41643;
    wire N__41640;
    wire N__41637;
    wire N__41636;
    wire N__41633;
    wire N__41630;
    wire N__41627;
    wire N__41624;
    wire N__41621;
    wire N__41618;
    wire N__41613;
    wire N__41610;
    wire N__41607;
    wire N__41604;
    wire N__41601;
    wire N__41600;
    wire N__41597;
    wire N__41596;
    wire N__41593;
    wire N__41590;
    wire N__41587;
    wire N__41584;
    wire N__41581;
    wire N__41578;
    wire N__41571;
    wire N__41570;
    wire N__41567;
    wire N__41564;
    wire N__41563;
    wire N__41560;
    wire N__41557;
    wire N__41554;
    wire N__41551;
    wire N__41546;
    wire N__41541;
    wire N__41538;
    wire N__41535;
    wire N__41532;
    wire N__41529;
    wire N__41526;
    wire N__41523;
    wire N__41520;
    wire N__41519;
    wire N__41516;
    wire N__41515;
    wire N__41514;
    wire N__41513;
    wire N__41512;
    wire N__41509;
    wire N__41506;
    wire N__41505;
    wire N__41504;
    wire N__41503;
    wire N__41502;
    wire N__41501;
    wire N__41498;
    wire N__41497;
    wire N__41496;
    wire N__41495;
    wire N__41494;
    wire N__41491;
    wire N__41490;
    wire N__41489;
    wire N__41486;
    wire N__41483;
    wire N__41482;
    wire N__41477;
    wire N__41472;
    wire N__41465;
    wire N__41462;
    wire N__41455;
    wire N__41446;
    wire N__41439;
    wire N__41432;
    wire N__41421;
    wire N__41420;
    wire N__41417;
    wire N__41414;
    wire N__41411;
    wire N__41408;
    wire N__41405;
    wire N__41402;
    wire N__41397;
    wire N__41394;
    wire N__41391;
    wire N__41388;
    wire N__41385;
    wire N__41382;
    wire N__41379;
    wire N__41378;
    wire N__41375;
    wire N__41374;
    wire N__41371;
    wire N__41370;
    wire N__41369;
    wire N__41368;
    wire N__41367;
    wire N__41366;
    wire N__41363;
    wire N__41360;
    wire N__41359;
    wire N__41358;
    wire N__41357;
    wire N__41356;
    wire N__41353;
    wire N__41350;
    wire N__41347;
    wire N__41344;
    wire N__41343;
    wire N__41342;
    wire N__41341;
    wire N__41340;
    wire N__41337;
    wire N__41334;
    wire N__41333;
    wire N__41332;
    wire N__41327;
    wire N__41324;
    wire N__41317;
    wire N__41314;
    wire N__41311;
    wire N__41298;
    wire N__41289;
    wire N__41274;
    wire N__41273;
    wire N__41272;
    wire N__41269;
    wire N__41266;
    wire N__41263;
    wire N__41260;
    wire N__41257;
    wire N__41254;
    wire N__41251;
    wire N__41248;
    wire N__41245;
    wire N__41240;
    wire N__41237;
    wire N__41234;
    wire N__41229;
    wire N__41228;
    wire N__41227;
    wire N__41224;
    wire N__41221;
    wire N__41218;
    wire N__41215;
    wire N__41212;
    wire N__41209;
    wire N__41206;
    wire N__41203;
    wire N__41200;
    wire N__41193;
    wire N__41190;
    wire N__41187;
    wire N__41184;
    wire N__41181;
    wire N__41178;
    wire N__41175;
    wire N__41172;
    wire N__41169;
    wire N__41166;
    wire N__41163;
    wire N__41160;
    wire N__41157;
    wire N__41154;
    wire N__41151;
    wire N__41148;
    wire N__41145;
    wire N__41142;
    wire N__41139;
    wire N__41136;
    wire N__41133;
    wire N__41132;
    wire N__41129;
    wire N__41126;
    wire N__41123;
    wire N__41120;
    wire N__41117;
    wire N__41114;
    wire N__41111;
    wire N__41106;
    wire N__41103;
    wire N__41100;
    wire N__41097;
    wire N__41094;
    wire N__41091;
    wire N__41088;
    wire N__41087;
    wire N__41084;
    wire N__41081;
    wire N__41078;
    wire N__41075;
    wire N__41070;
    wire N__41067;
    wire N__41064;
    wire N__41061;
    wire N__41058;
    wire N__41055;
    wire N__41052;
    wire N__41049;
    wire N__41046;
    wire N__41043;
    wire N__41040;
    wire N__41037;
    wire N__41034;
    wire N__41031;
    wire N__41028;
    wire N__41025;
    wire N__41022;
    wire N__41019;
    wire N__41016;
    wire N__41013;
    wire N__41010;
    wire N__41007;
    wire N__41004;
    wire N__41001;
    wire N__40998;
    wire N__40995;
    wire N__40992;
    wire N__40991;
    wire N__40990;
    wire N__40985;
    wire N__40982;
    wire N__40977;
    wire N__40974;
    wire N__40971;
    wire N__40970;
    wire N__40967;
    wire N__40964;
    wire N__40959;
    wire N__40956;
    wire N__40953;
    wire N__40950;
    wire N__40949;
    wire N__40948;
    wire N__40945;
    wire N__40942;
    wire N__40939;
    wire N__40934;
    wire N__40931;
    wire N__40928;
    wire N__40925;
    wire N__40920;
    wire N__40917;
    wire N__40914;
    wire N__40911;
    wire N__40910;
    wire N__40907;
    wire N__40904;
    wire N__40901;
    wire N__40898;
    wire N__40893;
    wire N__40890;
    wire N__40887;
    wire N__40884;
    wire N__40883;
    wire N__40880;
    wire N__40879;
    wire N__40876;
    wire N__40873;
    wire N__40870;
    wire N__40863;
    wire N__40860;
    wire N__40857;
    wire N__40854;
    wire N__40851;
    wire N__40848;
    wire N__40847;
    wire N__40844;
    wire N__40841;
    wire N__40836;
    wire N__40833;
    wire N__40830;
    wire N__40827;
    wire N__40824;
    wire N__40821;
    wire N__40818;
    wire N__40815;
    wire N__40812;
    wire N__40809;
    wire N__40806;
    wire N__40803;
    wire N__40800;
    wire N__40797;
    wire N__40794;
    wire N__40791;
    wire N__40788;
    wire N__40785;
    wire N__40784;
    wire N__40781;
    wire N__40780;
    wire N__40775;
    wire N__40772;
    wire N__40767;
    wire N__40764;
    wire N__40763;
    wire N__40762;
    wire N__40757;
    wire N__40754;
    wire N__40749;
    wire N__40746;
    wire N__40743;
    wire N__40742;
    wire N__40741;
    wire N__40736;
    wire N__40733;
    wire N__40728;
    wire N__40725;
    wire N__40722;
    wire N__40719;
    wire N__40716;
    wire N__40713;
    wire N__40710;
    wire N__40707;
    wire N__40704;
    wire N__40701;
    wire N__40698;
    wire N__40695;
    wire N__40692;
    wire N__40689;
    wire N__40686;
    wire N__40683;
    wire N__40680;
    wire N__40677;
    wire N__40674;
    wire N__40671;
    wire N__40668;
    wire N__40665;
    wire N__40662;
    wire N__40659;
    wire N__40656;
    wire N__40653;
    wire N__40650;
    wire N__40647;
    wire N__40644;
    wire N__40641;
    wire N__40638;
    wire N__40635;
    wire N__40632;
    wire N__40629;
    wire N__40626;
    wire N__40623;
    wire N__40620;
    wire N__40617;
    wire N__40614;
    wire N__40611;
    wire N__40608;
    wire N__40605;
    wire N__40602;
    wire N__40599;
    wire N__40596;
    wire N__40593;
    wire N__40590;
    wire N__40587;
    wire N__40584;
    wire N__40581;
    wire N__40578;
    wire N__40575;
    wire N__40572;
    wire N__40569;
    wire N__40566;
    wire N__40563;
    wire N__40562;
    wire N__40559;
    wire N__40556;
    wire N__40551;
    wire N__40548;
    wire N__40545;
    wire N__40542;
    wire N__40541;
    wire N__40538;
    wire N__40535;
    wire N__40532;
    wire N__40527;
    wire N__40526;
    wire N__40525;
    wire N__40524;
    wire N__40523;
    wire N__40522;
    wire N__40521;
    wire N__40520;
    wire N__40519;
    wire N__40518;
    wire N__40517;
    wire N__40516;
    wire N__40515;
    wire N__40514;
    wire N__40513;
    wire N__40512;
    wire N__40509;
    wire N__40508;
    wire N__40505;
    wire N__40504;
    wire N__40501;
    wire N__40500;
    wire N__40497;
    wire N__40496;
    wire N__40493;
    wire N__40492;
    wire N__40489;
    wire N__40488;
    wire N__40485;
    wire N__40484;
    wire N__40481;
    wire N__40480;
    wire N__40477;
    wire N__40476;
    wire N__40473;
    wire N__40472;
    wire N__40469;
    wire N__40468;
    wire N__40467;
    wire N__40464;
    wire N__40463;
    wire N__40460;
    wire N__40459;
    wire N__40456;
    wire N__40455;
    wire N__40438;
    wire N__40421;
    wire N__40404;
    wire N__40389;
    wire N__40386;
    wire N__40379;
    wire N__40374;
    wire N__40371;
    wire N__40368;
    wire N__40365;
    wire N__40362;
    wire N__40359;
    wire N__40356;
    wire N__40353;
    wire N__40350;
    wire N__40347;
    wire N__40344;
    wire N__40341;
    wire N__40338;
    wire N__40335;
    wire N__40332;
    wire N__40329;
    wire N__40326;
    wire N__40323;
    wire N__40320;
    wire N__40317;
    wire N__40314;
    wire N__40311;
    wire N__40308;
    wire N__40305;
    wire N__40304;
    wire N__40303;
    wire N__40302;
    wire N__40299;
    wire N__40296;
    wire N__40293;
    wire N__40290;
    wire N__40287;
    wire N__40284;
    wire N__40281;
    wire N__40278;
    wire N__40275;
    wire N__40272;
    wire N__40267;
    wire N__40260;
    wire N__40257;
    wire N__40254;
    wire N__40251;
    wire N__40248;
    wire N__40245;
    wire N__40242;
    wire N__40239;
    wire N__40236;
    wire N__40233;
    wire N__40232;
    wire N__40231;
    wire N__40230;
    wire N__40229;
    wire N__40228;
    wire N__40227;
    wire N__40226;
    wire N__40225;
    wire N__40224;
    wire N__40223;
    wire N__40222;
    wire N__40221;
    wire N__40220;
    wire N__40217;
    wire N__40214;
    wire N__40211;
    wire N__40210;
    wire N__40207;
    wire N__40206;
    wire N__40203;
    wire N__40200;
    wire N__40197;
    wire N__40194;
    wire N__40191;
    wire N__40188;
    wire N__40185;
    wire N__40182;
    wire N__40179;
    wire N__40176;
    wire N__40175;
    wire N__40174;
    wire N__40173;
    wire N__40172;
    wire N__40171;
    wire N__40170;
    wire N__40169;
    wire N__40164;
    wire N__40151;
    wire N__40142;
    wire N__40133;
    wire N__40130;
    wire N__40127;
    wire N__40124;
    wire N__40121;
    wire N__40118;
    wire N__40115;
    wire N__40112;
    wire N__40111;
    wire N__40102;
    wire N__40095;
    wire N__40084;
    wire N__40083;
    wire N__40080;
    wire N__40075;
    wire N__40072;
    wire N__40065;
    wire N__40062;
    wire N__40059;
    wire N__40056;
    wire N__40053;
    wire N__40050;
    wire N__40047;
    wire N__40044;
    wire N__40041;
    wire N__40038;
    wire N__40035;
    wire N__40032;
    wire N__40029;
    wire N__40026;
    wire N__40023;
    wire N__40020;
    wire N__40017;
    wire N__40014;
    wire N__40011;
    wire N__40008;
    wire N__40005;
    wire N__40002;
    wire N__40001;
    wire N__40000;
    wire N__39997;
    wire N__39994;
    wire N__39991;
    wire N__39988;
    wire N__39981;
    wire N__39978;
    wire N__39975;
    wire N__39972;
    wire N__39971;
    wire N__39970;
    wire N__39967;
    wire N__39964;
    wire N__39961;
    wire N__39958;
    wire N__39955;
    wire N__39952;
    wire N__39949;
    wire N__39946;
    wire N__39939;
    wire N__39936;
    wire N__39933;
    wire N__39930;
    wire N__39929;
    wire N__39928;
    wire N__39925;
    wire N__39922;
    wire N__39919;
    wire N__39916;
    wire N__39909;
    wire N__39906;
    wire N__39903;
    wire N__39900;
    wire N__39897;
    wire N__39894;
    wire N__39891;
    wire N__39888;
    wire N__39885;
    wire N__39882;
    wire N__39879;
    wire N__39876;
    wire N__39873;
    wire N__39870;
    wire N__39867;
    wire N__39864;
    wire N__39861;
    wire N__39858;
    wire N__39855;
    wire N__39852;
    wire N__39849;
    wire N__39846;
    wire N__39843;
    wire N__39840;
    wire N__39837;
    wire N__39834;
    wire N__39831;
    wire N__39828;
    wire N__39827;
    wire N__39826;
    wire N__39823;
    wire N__39818;
    wire N__39813;
    wire N__39810;
    wire N__39807;
    wire N__39804;
    wire N__39801;
    wire N__39800;
    wire N__39799;
    wire N__39796;
    wire N__39793;
    wire N__39790;
    wire N__39787;
    wire N__39780;
    wire N__39777;
    wire N__39774;
    wire N__39771;
    wire N__39768;
    wire N__39765;
    wire N__39764;
    wire N__39761;
    wire N__39760;
    wire N__39757;
    wire N__39754;
    wire N__39751;
    wire N__39748;
    wire N__39743;
    wire N__39738;
    wire N__39735;
    wire N__39732;
    wire N__39731;
    wire N__39728;
    wire N__39727;
    wire N__39724;
    wire N__39721;
    wire N__39718;
    wire N__39715;
    wire N__39712;
    wire N__39709;
    wire N__39702;
    wire N__39699;
    wire N__39696;
    wire N__39695;
    wire N__39692;
    wire N__39691;
    wire N__39688;
    wire N__39685;
    wire N__39682;
    wire N__39675;
    wire N__39672;
    wire N__39671;
    wire N__39668;
    wire N__39665;
    wire N__39664;
    wire N__39661;
    wire N__39658;
    wire N__39655;
    wire N__39648;
    wire N__39645;
    wire N__39642;
    wire N__39639;
    wire N__39636;
    wire N__39633;
    wire N__39632;
    wire N__39631;
    wire N__39628;
    wire N__39625;
    wire N__39622;
    wire N__39615;
    wire N__39612;
    wire N__39609;
    wire N__39608;
    wire N__39605;
    wire N__39602;
    wire N__39601;
    wire N__39598;
    wire N__39595;
    wire N__39592;
    wire N__39585;
    wire N__39582;
    wire N__39579;
    wire N__39578;
    wire N__39575;
    wire N__39572;
    wire N__39571;
    wire N__39568;
    wire N__39565;
    wire N__39562;
    wire N__39555;
    wire N__39552;
    wire N__39549;
    wire N__39546;
    wire N__39543;
    wire N__39540;
    wire N__39537;
    wire N__39536;
    wire N__39535;
    wire N__39532;
    wire N__39529;
    wire N__39526;
    wire N__39521;
    wire N__39518;
    wire N__39513;
    wire N__39510;
    wire N__39507;
    wire N__39506;
    wire N__39505;
    wire N__39502;
    wire N__39499;
    wire N__39496;
    wire N__39493;
    wire N__39490;
    wire N__39483;
    wire N__39480;
    wire N__39477;
    wire N__39474;
    wire N__39473;
    wire N__39470;
    wire N__39469;
    wire N__39466;
    wire N__39463;
    wire N__39460;
    wire N__39453;
    wire N__39450;
    wire N__39447;
    wire N__39444;
    wire N__39441;
    wire N__39440;
    wire N__39439;
    wire N__39436;
    wire N__39433;
    wire N__39430;
    wire N__39427;
    wire N__39424;
    wire N__39417;
    wire N__39414;
    wire N__39413;
    wire N__39410;
    wire N__39407;
    wire N__39404;
    wire N__39403;
    wire N__39400;
    wire N__39397;
    wire N__39394;
    wire N__39387;
    wire N__39384;
    wire N__39381;
    wire N__39380;
    wire N__39379;
    wire N__39376;
    wire N__39373;
    wire N__39370;
    wire N__39367;
    wire N__39364;
    wire N__39357;
    wire N__39354;
    wire N__39353;
    wire N__39350;
    wire N__39349;
    wire N__39346;
    wire N__39343;
    wire N__39340;
    wire N__39337;
    wire N__39334;
    wire N__39331;
    wire N__39328;
    wire N__39321;
    wire N__39320;
    wire N__39317;
    wire N__39314;
    wire N__39313;
    wire N__39310;
    wire N__39307;
    wire N__39304;
    wire N__39301;
    wire N__39298;
    wire N__39295;
    wire N__39292;
    wire N__39285;
    wire N__39282;
    wire N__39281;
    wire N__39280;
    wire N__39277;
    wire N__39274;
    wire N__39271;
    wire N__39268;
    wire N__39265;
    wire N__39262;
    wire N__39255;
    wire N__39252;
    wire N__39249;
    wire N__39246;
    wire N__39243;
    wire N__39242;
    wire N__39239;
    wire N__39236;
    wire N__39233;
    wire N__39230;
    wire N__39225;
    wire N__39224;
    wire N__39221;
    wire N__39218;
    wire N__39215;
    wire N__39214;
    wire N__39211;
    wire N__39208;
    wire N__39205;
    wire N__39198;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39188;
    wire N__39187;
    wire N__39186;
    wire N__39185;
    wire N__39184;
    wire N__39183;
    wire N__39182;
    wire N__39181;
    wire N__39176;
    wire N__39165;
    wire N__39160;
    wire N__39157;
    wire N__39150;
    wire N__39147;
    wire N__39144;
    wire N__39141;
    wire N__39138;
    wire N__39135;
    wire N__39132;
    wire N__39129;
    wire N__39126;
    wire N__39123;
    wire N__39122;
    wire N__39119;
    wire N__39118;
    wire N__39115;
    wire N__39112;
    wire N__39109;
    wire N__39106;
    wire N__39103;
    wire N__39100;
    wire N__39097;
    wire N__39090;
    wire N__39087;
    wire N__39084;
    wire N__39081;
    wire N__39078;
    wire N__39077;
    wire N__39074;
    wire N__39071;
    wire N__39070;
    wire N__39067;
    wire N__39064;
    wire N__39061;
    wire N__39054;
    wire N__39053;
    wire N__39052;
    wire N__39049;
    wire N__39046;
    wire N__39043;
    wire N__39040;
    wire N__39037;
    wire N__39030;
    wire N__39027;
    wire N__39026;
    wire N__39025;
    wire N__39022;
    wire N__39017;
    wire N__39012;
    wire N__39009;
    wire N__39006;
    wire N__39003;
    wire N__39002;
    wire N__39001;
    wire N__38998;
    wire N__38995;
    wire N__38992;
    wire N__38985;
    wire N__38982;
    wire N__38979;
    wire N__38976;
    wire N__38975;
    wire N__38974;
    wire N__38971;
    wire N__38966;
    wire N__38961;
    wire N__38958;
    wire N__38955;
    wire N__38954;
    wire N__38951;
    wire N__38950;
    wire N__38947;
    wire N__38942;
    wire N__38937;
    wire N__38934;
    wire N__38931;
    wire N__38928;
    wire N__38927;
    wire N__38924;
    wire N__38923;
    wire N__38920;
    wire N__38917;
    wire N__38914;
    wire N__38907;
    wire N__38904;
    wire N__38901;
    wire N__38898;
    wire N__38895;
    wire N__38892;
    wire N__38889;
    wire N__38886;
    wire N__38885;
    wire N__38882;
    wire N__38879;
    wire N__38874;
    wire N__38871;
    wire N__38870;
    wire N__38867;
    wire N__38864;
    wire N__38861;
    wire N__38858;
    wire N__38857;
    wire N__38854;
    wire N__38851;
    wire N__38848;
    wire N__38841;
    wire N__38838;
    wire N__38835;
    wire N__38832;
    wire N__38829;
    wire N__38826;
    wire N__38823;
    wire N__38820;
    wire N__38817;
    wire N__38814;
    wire N__38811;
    wire N__38808;
    wire N__38805;
    wire N__38802;
    wire N__38801;
    wire N__38800;
    wire N__38799;
    wire N__38796;
    wire N__38795;
    wire N__38792;
    wire N__38791;
    wire N__38788;
    wire N__38787;
    wire N__38772;
    wire N__38769;
    wire N__38766;
    wire N__38763;
    wire N__38760;
    wire N__38757;
    wire N__38754;
    wire N__38751;
    wire N__38748;
    wire N__38745;
    wire N__38742;
    wire N__38739;
    wire N__38736;
    wire N__38733;
    wire N__38730;
    wire N__38727;
    wire N__38724;
    wire N__38721;
    wire N__38718;
    wire N__38715;
    wire N__38712;
    wire N__38709;
    wire N__38706;
    wire N__38703;
    wire N__38700;
    wire N__38697;
    wire N__38694;
    wire N__38691;
    wire N__38688;
    wire N__38685;
    wire N__38682;
    wire N__38679;
    wire N__38676;
    wire N__38673;
    wire N__38670;
    wire N__38667;
    wire N__38664;
    wire N__38661;
    wire N__38658;
    wire N__38655;
    wire N__38652;
    wire N__38649;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38634;
    wire N__38631;
    wire N__38628;
    wire N__38625;
    wire N__38622;
    wire N__38619;
    wire N__38616;
    wire N__38613;
    wire N__38610;
    wire N__38607;
    wire N__38604;
    wire N__38601;
    wire N__38598;
    wire N__38595;
    wire N__38592;
    wire N__38589;
    wire N__38586;
    wire N__38583;
    wire N__38580;
    wire N__38577;
    wire N__38574;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38562;
    wire N__38559;
    wire N__38556;
    wire N__38553;
    wire N__38550;
    wire N__38547;
    wire N__38544;
    wire N__38541;
    wire N__38538;
    wire N__38535;
    wire N__38532;
    wire N__38529;
    wire N__38526;
    wire N__38523;
    wire N__38520;
    wire N__38517;
    wire N__38514;
    wire N__38511;
    wire N__38508;
    wire N__38505;
    wire N__38502;
    wire N__38499;
    wire N__38496;
    wire N__38493;
    wire N__38490;
    wire N__38487;
    wire N__38484;
    wire N__38481;
    wire N__38478;
    wire N__38475;
    wire N__38472;
    wire N__38469;
    wire N__38466;
    wire N__38463;
    wire N__38460;
    wire N__38457;
    wire N__38454;
    wire N__38451;
    wire N__38448;
    wire N__38445;
    wire N__38442;
    wire N__38439;
    wire N__38436;
    wire N__38433;
    wire N__38430;
    wire N__38427;
    wire N__38424;
    wire N__38421;
    wire N__38418;
    wire N__38415;
    wire N__38412;
    wire N__38409;
    wire N__38406;
    wire N__38403;
    wire N__38400;
    wire N__38397;
    wire N__38394;
    wire N__38391;
    wire N__38388;
    wire N__38385;
    wire N__38382;
    wire N__38379;
    wire N__38376;
    wire N__38373;
    wire N__38370;
    wire N__38367;
    wire N__38364;
    wire N__38361;
    wire N__38358;
    wire N__38355;
    wire N__38352;
    wire N__38349;
    wire N__38346;
    wire N__38345;
    wire N__38344;
    wire N__38341;
    wire N__38338;
    wire N__38335;
    wire N__38330;
    wire N__38327;
    wire N__38324;
    wire N__38321;
    wire N__38318;
    wire N__38313;
    wire N__38310;
    wire N__38307;
    wire N__38304;
    wire N__38301;
    wire N__38298;
    wire N__38295;
    wire N__38292;
    wire N__38289;
    wire N__38286;
    wire N__38283;
    wire N__38280;
    wire N__38277;
    wire N__38274;
    wire N__38271;
    wire N__38268;
    wire N__38265;
    wire N__38262;
    wire N__38259;
    wire N__38256;
    wire N__38253;
    wire N__38250;
    wire N__38247;
    wire N__38244;
    wire N__38241;
    wire N__38238;
    wire N__38235;
    wire N__38232;
    wire N__38229;
    wire N__38226;
    wire N__38223;
    wire N__38220;
    wire N__38217;
    wire N__38214;
    wire N__38211;
    wire N__38210;
    wire N__38207;
    wire N__38206;
    wire N__38203;
    wire N__38200;
    wire N__38197;
    wire N__38194;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38182;
    wire N__38179;
    wire N__38176;
    wire N__38169;
    wire N__38166;
    wire N__38163;
    wire N__38160;
    wire N__38159;
    wire N__38158;
    wire N__38153;
    wire N__38150;
    wire N__38147;
    wire N__38142;
    wire N__38139;
    wire N__38138;
    wire N__38137;
    wire N__38134;
    wire N__38131;
    wire N__38128;
    wire N__38123;
    wire N__38118;
    wire N__38117;
    wire N__38114;
    wire N__38111;
    wire N__38108;
    wire N__38107;
    wire N__38102;
    wire N__38099;
    wire N__38096;
    wire N__38093;
    wire N__38088;
    wire N__38087;
    wire N__38084;
    wire N__38081;
    wire N__38080;
    wire N__38075;
    wire N__38072;
    wire N__38067;
    wire N__38064;
    wire N__38061;
    wire N__38058;
    wire N__38055;
    wire N__38052;
    wire N__38049;
    wire N__38046;
    wire N__38043;
    wire N__38040;
    wire N__38037;
    wire N__38034;
    wire N__38031;
    wire N__38028;
    wire N__38027;
    wire N__38024;
    wire N__38021;
    wire N__38016;
    wire N__38013;
    wire N__38010;
    wire N__38007;
    wire N__38004;
    wire N__38001;
    wire N__37998;
    wire N__37995;
    wire N__37992;
    wire N__37989;
    wire N__37986;
    wire N__37983;
    wire N__37980;
    wire N__37977;
    wire N__37974;
    wire N__37971;
    wire N__37968;
    wire N__37965;
    wire N__37962;
    wire N__37959;
    wire N__37956;
    wire N__37953;
    wire N__37952;
    wire N__37949;
    wire N__37946;
    wire N__37943;
    wire N__37940;
    wire N__37937;
    wire N__37932;
    wire N__37929;
    wire N__37926;
    wire N__37925;
    wire N__37920;
    wire N__37917;
    wire N__37914;
    wire N__37911;
    wire N__37908;
    wire N__37907;
    wire N__37906;
    wire N__37903;
    wire N__37900;
    wire N__37897;
    wire N__37894;
    wire N__37891;
    wire N__37888;
    wire N__37881;
    wire N__37878;
    wire N__37875;
    wire N__37872;
    wire N__37869;
    wire N__37866;
    wire N__37863;
    wire N__37860;
    wire N__37857;
    wire N__37854;
    wire N__37851;
    wire N__37848;
    wire N__37845;
    wire N__37842;
    wire N__37839;
    wire N__37836;
    wire N__37833;
    wire N__37830;
    wire N__37827;
    wire N__37824;
    wire N__37821;
    wire N__37818;
    wire N__37815;
    wire N__37812;
    wire N__37809;
    wire N__37806;
    wire N__37803;
    wire N__37800;
    wire N__37797;
    wire N__37794;
    wire N__37791;
    wire N__37788;
    wire N__37785;
    wire N__37782;
    wire N__37779;
    wire N__37776;
    wire N__37773;
    wire N__37770;
    wire N__37767;
    wire N__37764;
    wire N__37761;
    wire N__37758;
    wire N__37755;
    wire N__37754;
    wire N__37753;
    wire N__37750;
    wire N__37747;
    wire N__37744;
    wire N__37741;
    wire N__37736;
    wire N__37731;
    wire N__37728;
    wire N__37725;
    wire N__37722;
    wire N__37719;
    wire N__37716;
    wire N__37715;
    wire N__37714;
    wire N__37711;
    wire N__37708;
    wire N__37705;
    wire N__37702;
    wire N__37699;
    wire N__37694;
    wire N__37689;
    wire N__37686;
    wire N__37683;
    wire N__37680;
    wire N__37677;
    wire N__37674;
    wire N__37673;
    wire N__37672;
    wire N__37669;
    wire N__37664;
    wire N__37659;
    wire N__37656;
    wire N__37653;
    wire N__37650;
    wire N__37647;
    wire N__37644;
    wire N__37641;
    wire N__37640;
    wire N__37639;
    wire N__37636;
    wire N__37633;
    wire N__37630;
    wire N__37627;
    wire N__37624;
    wire N__37621;
    wire N__37614;
    wire N__37611;
    wire N__37608;
    wire N__37605;
    wire N__37602;
    wire N__37599;
    wire N__37598;
    wire N__37595;
    wire N__37594;
    wire N__37591;
    wire N__37588;
    wire N__37585;
    wire N__37582;
    wire N__37579;
    wire N__37576;
    wire N__37573;
    wire N__37566;
    wire N__37563;
    wire N__37560;
    wire N__37557;
    wire N__37554;
    wire N__37551;
    wire N__37550;
    wire N__37549;
    wire N__37546;
    wire N__37543;
    wire N__37540;
    wire N__37535;
    wire N__37532;
    wire N__37529;
    wire N__37524;
    wire N__37521;
    wire N__37518;
    wire N__37515;
    wire N__37512;
    wire N__37509;
    wire N__37506;
    wire N__37503;
    wire N__37500;
    wire N__37497;
    wire N__37494;
    wire N__37491;
    wire N__37488;
    wire N__37485;
    wire N__37482;
    wire N__37479;
    wire N__37476;
    wire N__37473;
    wire N__37472;
    wire N__37471;
    wire N__37468;
    wire N__37465;
    wire N__37462;
    wire N__37459;
    wire N__37456;
    wire N__37449;
    wire N__37446;
    wire N__37443;
    wire N__37440;
    wire N__37437;
    wire N__37436;
    wire N__37433;
    wire N__37432;
    wire N__37429;
    wire N__37426;
    wire N__37423;
    wire N__37416;
    wire N__37413;
    wire N__37410;
    wire N__37407;
    wire N__37404;
    wire N__37403;
    wire N__37400;
    wire N__37399;
    wire N__37396;
    wire N__37393;
    wire N__37390;
    wire N__37383;
    wire N__37380;
    wire N__37377;
    wire N__37374;
    wire N__37373;
    wire N__37370;
    wire N__37367;
    wire N__37366;
    wire N__37361;
    wire N__37358;
    wire N__37353;
    wire N__37350;
    wire N__37347;
    wire N__37344;
    wire N__37341;
    wire N__37340;
    wire N__37337;
    wire N__37334;
    wire N__37333;
    wire N__37328;
    wire N__37325;
    wire N__37320;
    wire N__37317;
    wire N__37314;
    wire N__37311;
    wire N__37308;
    wire N__37307;
    wire N__37304;
    wire N__37301;
    wire N__37298;
    wire N__37293;
    wire N__37290;
    wire N__37287;
    wire N__37284;
    wire N__37281;
    wire N__37278;
    wire N__37277;
    wire N__37274;
    wire N__37273;
    wire N__37270;
    wire N__37267;
    wire N__37264;
    wire N__37257;
    wire N__37254;
    wire N__37251;
    wire N__37248;
    wire N__37247;
    wire N__37246;
    wire N__37243;
    wire N__37240;
    wire N__37237;
    wire N__37234;
    wire N__37231;
    wire N__37224;
    wire N__37221;
    wire N__37218;
    wire N__37215;
    wire N__37212;
    wire N__37211;
    wire N__37208;
    wire N__37207;
    wire N__37204;
    wire N__37201;
    wire N__37198;
    wire N__37195;
    wire N__37192;
    wire N__37185;
    wire N__37182;
    wire N__37179;
    wire N__37176;
    wire N__37173;
    wire N__37172;
    wire N__37169;
    wire N__37166;
    wire N__37165;
    wire N__37162;
    wire N__37157;
    wire N__37152;
    wire N__37149;
    wire N__37146;
    wire N__37143;
    wire N__37140;
    wire N__37139;
    wire N__37136;
    wire N__37133;
    wire N__37130;
    wire N__37129;
    wire N__37126;
    wire N__37123;
    wire N__37120;
    wire N__37113;
    wire N__37110;
    wire N__37107;
    wire N__37104;
    wire N__37101;
    wire N__37098;
    wire N__37095;
    wire N__37094;
    wire N__37091;
    wire N__37090;
    wire N__37087;
    wire N__37084;
    wire N__37081;
    wire N__37074;
    wire N__37071;
    wire N__37068;
    wire N__37065;
    wire N__37062;
    wire N__37059;
    wire N__37058;
    wire N__37055;
    wire N__37052;
    wire N__37049;
    wire N__37048;
    wire N__37045;
    wire N__37042;
    wire N__37039;
    wire N__37032;
    wire N__37029;
    wire N__37026;
    wire N__37023;
    wire N__37020;
    wire N__37019;
    wire N__37016;
    wire N__37015;
    wire N__37012;
    wire N__37009;
    wire N__37006;
    wire N__36999;
    wire N__36996;
    wire N__36993;
    wire N__36990;
    wire N__36987;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36976;
    wire N__36973;
    wire N__36970;
    wire N__36967;
    wire N__36960;
    wire N__36957;
    wire N__36954;
    wire N__36951;
    wire N__36948;
    wire N__36945;
    wire N__36942;
    wire N__36939;
    wire N__36936;
    wire N__36933;
    wire N__36932;
    wire N__36929;
    wire N__36926;
    wire N__36923;
    wire N__36918;
    wire N__36915;
    wire N__36912;
    wire N__36909;
    wire N__36906;
    wire N__36903;
    wire N__36900;
    wire N__36899;
    wire N__36896;
    wire N__36895;
    wire N__36892;
    wire N__36889;
    wire N__36886;
    wire N__36879;
    wire N__36876;
    wire N__36873;
    wire N__36870;
    wire N__36867;
    wire N__36866;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36856;
    wire N__36853;
    wire N__36846;
    wire N__36843;
    wire N__36840;
    wire N__36837;
    wire N__36834;
    wire N__36833;
    wire N__36832;
    wire N__36829;
    wire N__36826;
    wire N__36823;
    wire N__36820;
    wire N__36813;
    wire N__36810;
    wire N__36807;
    wire N__36804;
    wire N__36801;
    wire N__36800;
    wire N__36797;
    wire N__36794;
    wire N__36793;
    wire N__36790;
    wire N__36787;
    wire N__36784;
    wire N__36779;
    wire N__36774;
    wire N__36771;
    wire N__36768;
    wire N__36765;
    wire N__36762;
    wire N__36759;
    wire N__36758;
    wire N__36755;
    wire N__36752;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36738;
    wire N__36735;
    wire N__36732;
    wire N__36729;
    wire N__36726;
    wire N__36723;
    wire N__36720;
    wire N__36717;
    wire N__36716;
    wire N__36713;
    wire N__36712;
    wire N__36709;
    wire N__36706;
    wire N__36703;
    wire N__36696;
    wire N__36693;
    wire N__36690;
    wire N__36687;
    wire N__36684;
    wire N__36681;
    wire N__36678;
    wire N__36677;
    wire N__36674;
    wire N__36671;
    wire N__36668;
    wire N__36663;
    wire N__36660;
    wire N__36657;
    wire N__36654;
    wire N__36651;
    wire N__36648;
    wire N__36645;
    wire N__36642;
    wire N__36641;
    wire N__36638;
    wire N__36635;
    wire N__36632;
    wire N__36627;
    wire N__36624;
    wire N__36621;
    wire N__36618;
    wire N__36617;
    wire N__36614;
    wire N__36611;
    wire N__36608;
    wire N__36605;
    wire N__36602;
    wire N__36599;
    wire N__36594;
    wire N__36593;
    wire N__36592;
    wire N__36589;
    wire N__36586;
    wire N__36583;
    wire N__36576;
    wire N__36573;
    wire N__36570;
    wire N__36567;
    wire N__36564;
    wire N__36561;
    wire N__36558;
    wire N__36557;
    wire N__36554;
    wire N__36551;
    wire N__36548;
    wire N__36545;
    wire N__36540;
    wire N__36537;
    wire N__36534;
    wire N__36531;
    wire N__36528;
    wire N__36525;
    wire N__36522;
    wire N__36519;
    wire N__36516;
    wire N__36513;
    wire N__36510;
    wire N__36507;
    wire N__36504;
    wire N__36501;
    wire N__36498;
    wire N__36495;
    wire N__36492;
    wire N__36491;
    wire N__36488;
    wire N__36485;
    wire N__36482;
    wire N__36479;
    wire N__36476;
    wire N__36473;
    wire N__36468;
    wire N__36465;
    wire N__36462;
    wire N__36459;
    wire N__36458;
    wire N__36457;
    wire N__36456;
    wire N__36455;
    wire N__36454;
    wire N__36453;
    wire N__36450;
    wire N__36447;
    wire N__36446;
    wire N__36445;
    wire N__36442;
    wire N__36439;
    wire N__36438;
    wire N__36437;
    wire N__36434;
    wire N__36431;
    wire N__36430;
    wire N__36429;
    wire N__36428;
    wire N__36427;
    wire N__36426;
    wire N__36425;
    wire N__36424;
    wire N__36423;
    wire N__36422;
    wire N__36419;
    wire N__36418;
    wire N__36417;
    wire N__36412;
    wire N__36411;
    wire N__36410;
    wire N__36409;
    wire N__36408;
    wire N__36405;
    wire N__36402;
    wire N__36393;
    wire N__36380;
    wire N__36375;
    wire N__36370;
    wire N__36363;
    wire N__36360;
    wire N__36357;
    wire N__36354;
    wire N__36349;
    wire N__36342;
    wire N__36335;
    wire N__36330;
    wire N__36327;
    wire N__36312;
    wire N__36309;
    wire N__36306;
    wire N__36303;
    wire N__36300;
    wire N__36297;
    wire N__36296;
    wire N__36295;
    wire N__36294;
    wire N__36293;
    wire N__36292;
    wire N__36289;
    wire N__36286;
    wire N__36283;
    wire N__36282;
    wire N__36281;
    wire N__36280;
    wire N__36279;
    wire N__36278;
    wire N__36277;
    wire N__36276;
    wire N__36275;
    wire N__36272;
    wire N__36269;
    wire N__36268;
    wire N__36267;
    wire N__36266;
    wire N__36263;
    wire N__36262;
    wire N__36259;
    wire N__36258;
    wire N__36255;
    wire N__36252;
    wire N__36249;
    wire N__36246;
    wire N__36245;
    wire N__36242;
    wire N__36241;
    wire N__36240;
    wire N__36239;
    wire N__36236;
    wire N__36235;
    wire N__36234;
    wire N__36231;
    wire N__36228;
    wire N__36225;
    wire N__36224;
    wire N__36217;
    wire N__36212;
    wire N__36205;
    wire N__36202;
    wire N__36199;
    wire N__36194;
    wire N__36189;
    wire N__36184;
    wire N__36179;
    wire N__36170;
    wire N__36161;
    wire N__36154;
    wire N__36135;
    wire N__36132;
    wire N__36129;
    wire N__36126;
    wire N__36123;
    wire N__36120;
    wire N__36117;
    wire N__36114;
    wire N__36113;
    wire N__36110;
    wire N__36107;
    wire N__36102;
    wire N__36101;
    wire N__36100;
    wire N__36099;
    wire N__36098;
    wire N__36097;
    wire N__36096;
    wire N__36095;
    wire N__36094;
    wire N__36091;
    wire N__36090;
    wire N__36087;
    wire N__36086;
    wire N__36085;
    wire N__36082;
    wire N__36077;
    wire N__36074;
    wire N__36071;
    wire N__36070;
    wire N__36069;
    wire N__36068;
    wire N__36065;
    wire N__36058;
    wire N__36057;
    wire N__36054;
    wire N__36051;
    wire N__36050;
    wire N__36049;
    wire N__36048;
    wire N__36045;
    wire N__36044;
    wire N__36041;
    wire N__36038;
    wire N__36035;
    wire N__36032;
    wire N__36031;
    wire N__36030;
    wire N__36027;
    wire N__36024;
    wire N__36023;
    wire N__36020;
    wire N__36015;
    wire N__36012;
    wire N__36011;
    wire N__36008;
    wire N__35995;
    wire N__35986;
    wire N__35975;
    wire N__35968;
    wire N__35965;
    wire N__35952;
    wire N__35949;
    wire N__35948;
    wire N__35945;
    wire N__35942;
    wire N__35939;
    wire N__35936;
    wire N__35933;
    wire N__35930;
    wire N__35927;
    wire N__35924;
    wire N__35921;
    wire N__35918;
    wire N__35913;
    wire N__35912;
    wire N__35911;
    wire N__35908;
    wire N__35905;
    wire N__35904;
    wire N__35903;
    wire N__35902;
    wire N__35901;
    wire N__35900;
    wire N__35899;
    wire N__35898;
    wire N__35897;
    wire N__35896;
    wire N__35893;
    wire N__35890;
    wire N__35881;
    wire N__35878;
    wire N__35875;
    wire N__35874;
    wire N__35871;
    wire N__35870;
    wire N__35869;
    wire N__35868;
    wire N__35867;
    wire N__35866;
    wire N__35863;
    wire N__35862;
    wire N__35861;
    wire N__35860;
    wire N__35857;
    wire N__35856;
    wire N__35855;
    wire N__35852;
    wire N__35847;
    wire N__35844;
    wire N__35839;
    wire N__35832;
    wire N__35829;
    wire N__35822;
    wire N__35813;
    wire N__35806;
    wire N__35801;
    wire N__35796;
    wire N__35781;
    wire N__35778;
    wire N__35775;
    wire N__35772;
    wire N__35769;
    wire N__35766;
    wire N__35765;
    wire N__35762;
    wire N__35759;
    wire N__35754;
    wire N__35751;
    wire N__35748;
    wire N__35747;
    wire N__35746;
    wire N__35745;
    wire N__35744;
    wire N__35743;
    wire N__35742;
    wire N__35741;
    wire N__35740;
    wire N__35739;
    wire N__35738;
    wire N__35735;
    wire N__35730;
    wire N__35727;
    wire N__35724;
    wire N__35723;
    wire N__35722;
    wire N__35719;
    wire N__35718;
    wire N__35717;
    wire N__35716;
    wire N__35713;
    wire N__35710;
    wire N__35709;
    wire N__35708;
    wire N__35705;
    wire N__35704;
    wire N__35703;
    wire N__35702;
    wire N__35699;
    wire N__35696;
    wire N__35695;
    wire N__35690;
    wire N__35687;
    wire N__35684;
    wire N__35675;
    wire N__35670;
    wire N__35663;
    wire N__35656;
    wire N__35645;
    wire N__35628;
    wire N__35625;
    wire N__35622;
    wire N__35619;
    wire N__35616;
    wire N__35613;
    wire N__35612;
    wire N__35609;
    wire N__35606;
    wire N__35601;
    wire N__35598;
    wire N__35597;
    wire N__35596;
    wire N__35595;
    wire N__35594;
    wire N__35591;
    wire N__35590;
    wire N__35589;
    wire N__35588;
    wire N__35587;
    wire N__35584;
    wire N__35581;
    wire N__35578;
    wire N__35575;
    wire N__35574;
    wire N__35573;
    wire N__35570;
    wire N__35567;
    wire N__35566;
    wire N__35563;
    wire N__35562;
    wire N__35561;
    wire N__35558;
    wire N__35555;
    wire N__35554;
    wire N__35551;
    wire N__35542;
    wire N__35541;
    wire N__35540;
    wire N__35539;
    wire N__35538;
    wire N__35537;
    wire N__35534;
    wire N__35533;
    wire N__35530;
    wire N__35525;
    wire N__35518;
    wire N__35511;
    wire N__35506;
    wire N__35501;
    wire N__35490;
    wire N__35475;
    wire N__35472;
    wire N__35469;
    wire N__35466;
    wire N__35463;
    wire N__35462;
    wire N__35459;
    wire N__35456;
    wire N__35451;
    wire N__35448;
    wire N__35447;
    wire N__35446;
    wire N__35445;
    wire N__35444;
    wire N__35443;
    wire N__35442;
    wire N__35441;
    wire N__35438;
    wire N__35437;
    wire N__35436;
    wire N__35433;
    wire N__35430;
    wire N__35427;
    wire N__35424;
    wire N__35421;
    wire N__35420;
    wire N__35419;
    wire N__35418;
    wire N__35417;
    wire N__35416;
    wire N__35413;
    wire N__35410;
    wire N__35409;
    wire N__35408;
    wire N__35405;
    wire N__35400;
    wire N__35399;
    wire N__35396;
    wire N__35391;
    wire N__35380;
    wire N__35379;
    wire N__35378;
    wire N__35373;
    wire N__35364;
    wire N__35359;
    wire N__35356;
    wire N__35353;
    wire N__35348;
    wire N__35343;
    wire N__35328;
    wire N__35325;
    wire N__35322;
    wire N__35319;
    wire N__35316;
    wire N__35315;
    wire N__35312;
    wire N__35309;
    wire N__35304;
    wire N__35303;
    wire N__35302;
    wire N__35299;
    wire N__35298;
    wire N__35297;
    wire N__35296;
    wire N__35293;
    wire N__35292;
    wire N__35289;
    wire N__35288;
    wire N__35285;
    wire N__35282;
    wire N__35281;
    wire N__35280;
    wire N__35279;
    wire N__35278;
    wire N__35277;
    wire N__35276;
    wire N__35271;
    wire N__35266;
    wire N__35263;
    wire N__35262;
    wire N__35259;
    wire N__35258;
    wire N__35257;
    wire N__35254;
    wire N__35251;
    wire N__35248;
    wire N__35245;
    wire N__35244;
    wire N__35243;
    wire N__35240;
    wire N__35233;
    wire N__35230;
    wire N__35225;
    wire N__35218;
    wire N__35215;
    wire N__35210;
    wire N__35203;
    wire N__35200;
    wire N__35181;
    wire N__35178;
    wire N__35177;
    wire N__35176;
    wire N__35173;
    wire N__35170;
    wire N__35167;
    wire N__35164;
    wire N__35161;
    wire N__35158;
    wire N__35153;
    wire N__35148;
    wire N__35145;
    wire N__35142;
    wire N__35141;
    wire N__35138;
    wire N__35137;
    wire N__35134;
    wire N__35131;
    wire N__35128;
    wire N__35125;
    wire N__35118;
    wire N__35115;
    wire N__35112;
    wire N__35109;
    wire N__35106;
    wire N__35103;
    wire N__35100;
    wire N__35099;
    wire N__35096;
    wire N__35095;
    wire N__35094;
    wire N__35093;
    wire N__35092;
    wire N__35091;
    wire N__35090;
    wire N__35089;
    wire N__35088;
    wire N__35087;
    wire N__35084;
    wire N__35081;
    wire N__35080;
    wire N__35079;
    wire N__35078;
    wire N__35077;
    wire N__35076;
    wire N__35073;
    wire N__35072;
    wire N__35069;
    wire N__35068;
    wire N__35067;
    wire N__35066;
    wire N__35063;
    wire N__35058;
    wire N__35057;
    wire N__35054;
    wire N__35051;
    wire N__35050;
    wire N__35049;
    wire N__35046;
    wire N__35045;
    wire N__35042;
    wire N__35041;
    wire N__35040;
    wire N__35039;
    wire N__35038;
    wire N__35037;
    wire N__35036;
    wire N__35035;
    wire N__35032;
    wire N__35029;
    wire N__35016;
    wire N__35003;
    wire N__35000;
    wire N__34987;
    wire N__34980;
    wire N__34967;
    wire N__34950;
    wire N__34947;
    wire N__34944;
    wire N__34941;
    wire N__34940;
    wire N__34937;
    wire N__34934;
    wire N__34931;
    wire N__34928;
    wire N__34923;
    wire N__34922;
    wire N__34919;
    wire N__34918;
    wire N__34917;
    wire N__34916;
    wire N__34915;
    wire N__34912;
    wire N__34911;
    wire N__34910;
    wire N__34909;
    wire N__34908;
    wire N__34907;
    wire N__34906;
    wire N__34901;
    wire N__34898;
    wire N__34895;
    wire N__34892;
    wire N__34891;
    wire N__34890;
    wire N__34889;
    wire N__34888;
    wire N__34885;
    wire N__34882;
    wire N__34881;
    wire N__34880;
    wire N__34877;
    wire N__34876;
    wire N__34875;
    wire N__34874;
    wire N__34871;
    wire N__34870;
    wire N__34867;
    wire N__34866;
    wire N__34863;
    wire N__34862;
    wire N__34859;
    wire N__34858;
    wire N__34855;
    wire N__34852;
    wire N__34843;
    wire N__34840;
    wire N__34839;
    wire N__34836;
    wire N__34835;
    wire N__34832;
    wire N__34829;
    wire N__34826;
    wire N__34825;
    wire N__34824;
    wire N__34823;
    wire N__34814;
    wire N__34807;
    wire N__34802;
    wire N__34793;
    wire N__34790;
    wire N__34783;
    wire N__34776;
    wire N__34771;
    wire N__34762;
    wire N__34743;
    wire N__34740;
    wire N__34739;
    wire N__34736;
    wire N__34733;
    wire N__34730;
    wire N__34727;
    wire N__34724;
    wire N__34721;
    wire N__34716;
    wire N__34715;
    wire N__34714;
    wire N__34711;
    wire N__34710;
    wire N__34709;
    wire N__34708;
    wire N__34705;
    wire N__34704;
    wire N__34703;
    wire N__34700;
    wire N__34699;
    wire N__34698;
    wire N__34697;
    wire N__34696;
    wire N__34695;
    wire N__34690;
    wire N__34687;
    wire N__34686;
    wire N__34683;
    wire N__34682;
    wire N__34681;
    wire N__34678;
    wire N__34673;
    wire N__34666;
    wire N__34665;
    wire N__34664;
    wire N__34661;
    wire N__34660;
    wire N__34659;
    wire N__34658;
    wire N__34657;
    wire N__34654;
    wire N__34653;
    wire N__34650;
    wire N__34649;
    wire N__34646;
    wire N__34635;
    wire N__34632;
    wire N__34627;
    wire N__34620;
    wire N__34617;
    wire N__34614;
    wire N__34613;
    wire N__34612;
    wire N__34611;
    wire N__34608;
    wire N__34605;
    wire N__34604;
    wire N__34603;
    wire N__34594;
    wire N__34589;
    wire N__34582;
    wire N__34579;
    wire N__34576;
    wire N__34563;
    wire N__34560;
    wire N__34555;
    wire N__34542;
    wire N__34539;
    wire N__34536;
    wire N__34533;
    wire N__34532;
    wire N__34529;
    wire N__34526;
    wire N__34523;
    wire N__34520;
    wire N__34515;
    wire N__34514;
    wire N__34513;
    wire N__34512;
    wire N__34511;
    wire N__34510;
    wire N__34509;
    wire N__34506;
    wire N__34505;
    wire N__34504;
    wire N__34503;
    wire N__34502;
    wire N__34499;
    wire N__34494;
    wire N__34493;
    wire N__34490;
    wire N__34487;
    wire N__34484;
    wire N__34483;
    wire N__34480;
    wire N__34479;
    wire N__34476;
    wire N__34475;
    wire N__34474;
    wire N__34473;
    wire N__34472;
    wire N__34469;
    wire N__34468;
    wire N__34467;
    wire N__34466;
    wire N__34463;
    wire N__34462;
    wire N__34461;
    wire N__34460;
    wire N__34459;
    wire N__34458;
    wire N__34455;
    wire N__34454;
    wire N__34453;
    wire N__34450;
    wire N__34447;
    wire N__34436;
    wire N__34433;
    wire N__34430;
    wire N__34427;
    wire N__34420;
    wire N__34413;
    wire N__34406;
    wire N__34403;
    wire N__34398;
    wire N__34387;
    wire N__34380;
    wire N__34359;
    wire N__34356;
    wire N__34353;
    wire N__34352;
    wire N__34349;
    wire N__34346;
    wire N__34341;
    wire N__34338;
    wire N__34335;
    wire N__34334;
    wire N__34333;
    wire N__34332;
    wire N__34329;
    wire N__34328;
    wire N__34325;
    wire N__34324;
    wire N__34323;
    wire N__34322;
    wire N__34321;
    wire N__34320;
    wire N__34317;
    wire N__34316;
    wire N__34315;
    wire N__34314;
    wire N__34311;
    wire N__34306;
    wire N__34303;
    wire N__34302;
    wire N__34301;
    wire N__34298;
    wire N__34297;
    wire N__34294;
    wire N__34293;
    wire N__34292;
    wire N__34291;
    wire N__34290;
    wire N__34289;
    wire N__34286;
    wire N__34283;
    wire N__34282;
    wire N__34279;
    wire N__34278;
    wire N__34277;
    wire N__34272;
    wire N__34271;
    wire N__34268;
    wire N__34267;
    wire N__34264;
    wire N__34263;
    wire N__34260;
    wire N__34257;
    wire N__34254;
    wire N__34249;
    wire N__34244;
    wire N__34239;
    wire N__34230;
    wire N__34227;
    wire N__34222;
    wire N__34215;
    wire N__34212;
    wire N__34201;
    wire N__34196;
    wire N__34173;
    wire N__34170;
    wire N__34167;
    wire N__34166;
    wire N__34165;
    wire N__34162;
    wire N__34159;
    wire N__34156;
    wire N__34151;
    wire N__34148;
    wire N__34145;
    wire N__34142;
    wire N__34139;
    wire N__34134;
    wire N__34131;
    wire N__34128;
    wire N__34125;
    wire N__34122;
    wire N__34119;
    wire N__34118;
    wire N__34115;
    wire N__34112;
    wire N__34109;
    wire N__34106;
    wire N__34103;
    wire N__34102;
    wire N__34099;
    wire N__34096;
    wire N__34093;
    wire N__34086;
    wire N__34083;
    wire N__34082;
    wire N__34079;
    wire N__34076;
    wire N__34075;
    wire N__34072;
    wire N__34069;
    wire N__34066;
    wire N__34061;
    wire N__34058;
    wire N__34053;
    wire N__34050;
    wire N__34047;
    wire N__34044;
    wire N__34043;
    wire N__34040;
    wire N__34037;
    wire N__34034;
    wire N__34031;
    wire N__34030;
    wire N__34027;
    wire N__34024;
    wire N__34021;
    wire N__34014;
    wire N__34011;
    wire N__34010;
    wire N__34007;
    wire N__34004;
    wire N__34001;
    wire N__33998;
    wire N__33997;
    wire N__33992;
    wire N__33989;
    wire N__33984;
    wire N__33983;
    wire N__33980;
    wire N__33977;
    wire N__33974;
    wire N__33969;
    wire N__33968;
    wire N__33965;
    wire N__33962;
    wire N__33957;
    wire N__33954;
    wire N__33951;
    wire N__33948;
    wire N__33945;
    wire N__33944;
    wire N__33941;
    wire N__33938;
    wire N__33933;
    wire N__33930;
    wire N__33927;
    wire N__33924;
    wire N__33921;
    wire N__33918;
    wire N__33917;
    wire N__33914;
    wire N__33911;
    wire N__33908;
    wire N__33907;
    wire N__33904;
    wire N__33901;
    wire N__33898;
    wire N__33891;
    wire N__33888;
    wire N__33885;
    wire N__33882;
    wire N__33879;
    wire N__33878;
    wire N__33875;
    wire N__33872;
    wire N__33871;
    wire N__33868;
    wire N__33865;
    wire N__33862;
    wire N__33859;
    wire N__33856;
    wire N__33853;
    wire N__33850;
    wire N__33845;
    wire N__33840;
    wire N__33839;
    wire N__33836;
    wire N__33833;
    wire N__33832;
    wire N__33829;
    wire N__33826;
    wire N__33823;
    wire N__33816;
    wire N__33813;
    wire N__33810;
    wire N__33807;
    wire N__33806;
    wire N__33805;
    wire N__33802;
    wire N__33799;
    wire N__33796;
    wire N__33793;
    wire N__33790;
    wire N__33787;
    wire N__33780;
    wire N__33777;
    wire N__33776;
    wire N__33775;
    wire N__33772;
    wire N__33769;
    wire N__33766;
    wire N__33763;
    wire N__33760;
    wire N__33757;
    wire N__33750;
    wire N__33747;
    wire N__33744;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33732;
    wire N__33731;
    wire N__33728;
    wire N__33725;
    wire N__33722;
    wire N__33721;
    wire N__33718;
    wire N__33715;
    wire N__33712;
    wire N__33705;
    wire N__33704;
    wire N__33701;
    wire N__33698;
    wire N__33695;
    wire N__33692;
    wire N__33687;
    wire N__33684;
    wire N__33681;
    wire N__33678;
    wire N__33677;
    wire N__33674;
    wire N__33671;
    wire N__33668;
    wire N__33665;
    wire N__33662;
    wire N__33661;
    wire N__33658;
    wire N__33655;
    wire N__33652;
    wire N__33645;
    wire N__33642;
    wire N__33639;
    wire N__33636;
    wire N__33633;
    wire N__33632;
    wire N__33629;
    wire N__33626;
    wire N__33621;
    wire N__33620;
    wire N__33617;
    wire N__33614;
    wire N__33609;
    wire N__33606;
    wire N__33605;
    wire N__33602;
    wire N__33601;
    wire N__33598;
    wire N__33595;
    wire N__33592;
    wire N__33589;
    wire N__33582;
    wire N__33581;
    wire N__33578;
    wire N__33577;
    wire N__33574;
    wire N__33571;
    wire N__33568;
    wire N__33565;
    wire N__33562;
    wire N__33559;
    wire N__33556;
    wire N__33553;
    wire N__33548;
    wire N__33545;
    wire N__33540;
    wire N__33539;
    wire N__33536;
    wire N__33533;
    wire N__33530;
    wire N__33527;
    wire N__33524;
    wire N__33523;
    wire N__33520;
    wire N__33517;
    wire N__33514;
    wire N__33509;
    wire N__33506;
    wire N__33501;
    wire N__33500;
    wire N__33497;
    wire N__33496;
    wire N__33493;
    wire N__33490;
    wire N__33487;
    wire N__33484;
    wire N__33481;
    wire N__33478;
    wire N__33473;
    wire N__33470;
    wire N__33465;
    wire N__33464;
    wire N__33461;
    wire N__33458;
    wire N__33455;
    wire N__33452;
    wire N__33447;
    wire N__33444;
    wire N__33443;
    wire N__33440;
    wire N__33437;
    wire N__33436;
    wire N__33433;
    wire N__33430;
    wire N__33427;
    wire N__33420;
    wire N__33419;
    wire N__33416;
    wire N__33413;
    wire N__33412;
    wire N__33409;
    wire N__33406;
    wire N__33403;
    wire N__33396;
    wire N__33393;
    wire N__33392;
    wire N__33389;
    wire N__33386;
    wire N__33385;
    wire N__33382;
    wire N__33379;
    wire N__33376;
    wire N__33369;
    wire N__33368;
    wire N__33365;
    wire N__33362;
    wire N__33359;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33345;
    wire N__33342;
    wire N__33341;
    wire N__33338;
    wire N__33335;
    wire N__33334;
    wire N__33331;
    wire N__33328;
    wire N__33325;
    wire N__33318;
    wire N__33315;
    wire N__33314;
    wire N__33311;
    wire N__33308;
    wire N__33307;
    wire N__33304;
    wire N__33301;
    wire N__33298;
    wire N__33291;
    wire N__33288;
    wire N__33287;
    wire N__33286;
    wire N__33283;
    wire N__33280;
    wire N__33277;
    wire N__33270;
    wire N__33269;
    wire N__33268;
    wire N__33265;
    wire N__33262;
    wire N__33259;
    wire N__33256;
    wire N__33253;
    wire N__33250;
    wire N__33243;
    wire N__33240;
    wire N__33237;
    wire N__33234;
    wire N__33231;
    wire N__33228;
    wire N__33227;
    wire N__33224;
    wire N__33221;
    wire N__33220;
    wire N__33217;
    wire N__33214;
    wire N__33211;
    wire N__33208;
    wire N__33205;
    wire N__33202;
    wire N__33195;
    wire N__33192;
    wire N__33189;
    wire N__33186;
    wire N__33183;
    wire N__33180;
    wire N__33177;
    wire N__33176;
    wire N__33175;
    wire N__33172;
    wire N__33167;
    wire N__33162;
    wire N__33159;
    wire N__33156;
    wire N__33153;
    wire N__33150;
    wire N__33147;
    wire N__33144;
    wire N__33141;
    wire N__33140;
    wire N__33137;
    wire N__33134;
    wire N__33131;
    wire N__33128;
    wire N__33123;
    wire N__33120;
    wire N__33117;
    wire N__33114;
    wire N__33111;
    wire N__33110;
    wire N__33107;
    wire N__33104;
    wire N__33103;
    wire N__33098;
    wire N__33095;
    wire N__33092;
    wire N__33089;
    wire N__33084;
    wire N__33083;
    wire N__33080;
    wire N__33077;
    wire N__33074;
    wire N__33071;
    wire N__33066;
    wire N__33063;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33051;
    wire N__33048;
    wire N__33045;
    wire N__33042;
    wire N__33039;
    wire N__33036;
    wire N__33033;
    wire N__33030;
    wire N__33027;
    wire N__33024;
    wire N__33021;
    wire N__33018;
    wire N__33015;
    wire N__33012;
    wire N__33009;
    wire N__33006;
    wire N__33003;
    wire N__33000;
    wire N__32997;
    wire N__32994;
    wire N__32991;
    wire N__32988;
    wire N__32985;
    wire N__32982;
    wire N__32979;
    wire N__32976;
    wire N__32973;
    wire N__32970;
    wire N__32967;
    wire N__32964;
    wire N__32961;
    wire N__32958;
    wire N__32957;
    wire N__32954;
    wire N__32951;
    wire N__32946;
    wire N__32943;
    wire N__32940;
    wire N__32937;
    wire N__32934;
    wire N__32931;
    wire N__32928;
    wire N__32925;
    wire N__32922;
    wire N__32919;
    wire N__32916;
    wire N__32915;
    wire N__32912;
    wire N__32909;
    wire N__32906;
    wire N__32905;
    wire N__32902;
    wire N__32899;
    wire N__32896;
    wire N__32889;
    wire N__32886;
    wire N__32883;
    wire N__32880;
    wire N__32877;
    wire N__32874;
    wire N__32871;
    wire N__32868;
    wire N__32865;
    wire N__32862;
    wire N__32859;
    wire N__32858;
    wire N__32855;
    wire N__32852;
    wire N__32849;
    wire N__32844;
    wire N__32841;
    wire N__32838;
    wire N__32835;
    wire N__32832;
    wire N__32829;
    wire N__32826;
    wire N__32823;
    wire N__32822;
    wire N__32819;
    wire N__32818;
    wire N__32815;
    wire N__32812;
    wire N__32809;
    wire N__32802;
    wire N__32799;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32781;
    wire N__32780;
    wire N__32777;
    wire N__32774;
    wire N__32769;
    wire N__32766;
    wire N__32763;
    wire N__32760;
    wire N__32757;
    wire N__32754;
    wire N__32751;
    wire N__32750;
    wire N__32747;
    wire N__32744;
    wire N__32739;
    wire N__32736;
    wire N__32733;
    wire N__32732;
    wire N__32729;
    wire N__32726;
    wire N__32723;
    wire N__32722;
    wire N__32717;
    wire N__32714;
    wire N__32709;
    wire N__32706;
    wire N__32703;
    wire N__32702;
    wire N__32699;
    wire N__32696;
    wire N__32695;
    wire N__32692;
    wire N__32689;
    wire N__32686;
    wire N__32679;
    wire N__32676;
    wire N__32673;
    wire N__32670;
    wire N__32667;
    wire N__32664;
    wire N__32661;
    wire N__32658;
    wire N__32657;
    wire N__32654;
    wire N__32651;
    wire N__32648;
    wire N__32645;
    wire N__32642;
    wire N__32637;
    wire N__32634;
    wire N__32631;
    wire N__32628;
    wire N__32625;
    wire N__32624;
    wire N__32621;
    wire N__32618;
    wire N__32617;
    wire N__32614;
    wire N__32611;
    wire N__32608;
    wire N__32605;
    wire N__32600;
    wire N__32595;
    wire N__32592;
    wire N__32591;
    wire N__32588;
    wire N__32585;
    wire N__32580;
    wire N__32579;
    wire N__32576;
    wire N__32573;
    wire N__32568;
    wire N__32565;
    wire N__32562;
    wire N__32559;
    wire N__32556;
    wire N__32555;
    wire N__32552;
    wire N__32549;
    wire N__32548;
    wire N__32545;
    wire N__32542;
    wire N__32539;
    wire N__32536;
    wire N__32531;
    wire N__32526;
    wire N__32523;
    wire N__32520;
    wire N__32517;
    wire N__32514;
    wire N__32513;
    wire N__32510;
    wire N__32507;
    wire N__32504;
    wire N__32499;
    wire N__32496;
    wire N__32493;
    wire N__32490;
    wire N__32487;
    wire N__32484;
    wire N__32481;
    wire N__32478;
    wire N__32475;
    wire N__32472;
    wire N__32469;
    wire N__32466;
    wire N__32463;
    wire N__32460;
    wire N__32457;
    wire N__32454;
    wire N__32451;
    wire N__32450;
    wire N__32447;
    wire N__32446;
    wire N__32443;
    wire N__32440;
    wire N__32437;
    wire N__32430;
    wire N__32427;
    wire N__32424;
    wire N__32421;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32409;
    wire N__32408;
    wire N__32405;
    wire N__32404;
    wire N__32401;
    wire N__32398;
    wire N__32395;
    wire N__32388;
    wire N__32385;
    wire N__32382;
    wire N__32379;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32358;
    wire N__32355;
    wire N__32352;
    wire N__32349;
    wire N__32348;
    wire N__32345;
    wire N__32342;
    wire N__32339;
    wire N__32336;
    wire N__32331;
    wire N__32330;
    wire N__32327;
    wire N__32324;
    wire N__32319;
    wire N__32316;
    wire N__32313;
    wire N__32310;
    wire N__32307;
    wire N__32306;
    wire N__32305;
    wire N__32302;
    wire N__32299;
    wire N__32296;
    wire N__32293;
    wire N__32288;
    wire N__32283;
    wire N__32280;
    wire N__32277;
    wire N__32274;
    wire N__32271;
    wire N__32270;
    wire N__32267;
    wire N__32264;
    wire N__32261;
    wire N__32258;
    wire N__32253;
    wire N__32250;
    wire N__32247;
    wire N__32244;
    wire N__32241;
    wire N__32240;
    wire N__32237;
    wire N__32234;
    wire N__32233;
    wire N__32230;
    wire N__32227;
    wire N__32224;
    wire N__32217;
    wire N__32214;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32199;
    wire N__32196;
    wire N__32193;
    wire N__32190;
    wire N__32189;
    wire N__32186;
    wire N__32183;
    wire N__32178;
    wire N__32175;
    wire N__32172;
    wire N__32169;
    wire N__32166;
    wire N__32163;
    wire N__32160;
    wire N__32157;
    wire N__32156;
    wire N__32153;
    wire N__32150;
    wire N__32145;
    wire N__32142;
    wire N__32139;
    wire N__32136;
    wire N__32133;
    wire N__32130;
    wire N__32127;
    wire N__32124;
    wire N__32121;
    wire N__32120;
    wire N__32117;
    wire N__32114;
    wire N__32109;
    wire N__32106;
    wire N__32103;
    wire N__32100;
    wire N__32097;
    wire N__32094;
    wire N__32091;
    wire N__32090;
    wire N__32087;
    wire N__32084;
    wire N__32081;
    wire N__32078;
    wire N__32075;
    wire N__32070;
    wire N__32067;
    wire N__32064;
    wire N__32061;
    wire N__32058;
    wire N__32055;
    wire N__32054;
    wire N__32053;
    wire N__32050;
    wire N__32047;
    wire N__32042;
    wire N__32037;
    wire N__32034;
    wire N__32031;
    wire N__32028;
    wire N__32025;
    wire N__32022;
    wire N__32019;
    wire N__32016;
    wire N__32015;
    wire N__32012;
    wire N__32009;
    wire N__32008;
    wire N__32003;
    wire N__32000;
    wire N__31995;
    wire N__31992;
    wire N__31989;
    wire N__31986;
    wire N__31983;
    wire N__31980;
    wire N__31979;
    wire N__31976;
    wire N__31973;
    wire N__31972;
    wire N__31969;
    wire N__31966;
    wire N__31963;
    wire N__31956;
    wire N__31953;
    wire N__31950;
    wire N__31947;
    wire N__31944;
    wire N__31941;
    wire N__31940;
    wire N__31937;
    wire N__31934;
    wire N__31929;
    wire N__31926;
    wire N__31923;
    wire N__31920;
    wire N__31917;
    wire N__31916;
    wire N__31913;
    wire N__31910;
    wire N__31909;
    wire N__31906;
    wire N__31903;
    wire N__31900;
    wire N__31893;
    wire N__31890;
    wire N__31887;
    wire N__31884;
    wire N__31881;
    wire N__31878;
    wire N__31875;
    wire N__31872;
    wire N__31869;
    wire N__31866;
    wire N__31865;
    wire N__31862;
    wire N__31859;
    wire N__31856;
    wire N__31851;
    wire N__31848;
    wire N__31845;
    wire N__31842;
    wire N__31839;
    wire N__31836;
    wire N__31835;
    wire N__31834;
    wire N__31831;
    wire N__31826;
    wire N__31821;
    wire N__31818;
    wire N__31815;
    wire N__31812;
    wire N__31809;
    wire N__31808;
    wire N__31805;
    wire N__31802;
    wire N__31799;
    wire N__31798;
    wire N__31793;
    wire N__31790;
    wire N__31785;
    wire N__31782;
    wire N__31779;
    wire N__31776;
    wire N__31773;
    wire N__31770;
    wire N__31767;
    wire N__31764;
    wire N__31761;
    wire N__31760;
    wire N__31757;
    wire N__31754;
    wire N__31753;
    wire N__31750;
    wire N__31747;
    wire N__31744;
    wire N__31737;
    wire N__31734;
    wire N__31731;
    wire N__31728;
    wire N__31727;
    wire N__31724;
    wire N__31721;
    wire N__31718;
    wire N__31715;
    wire N__31710;
    wire N__31707;
    wire N__31704;
    wire N__31701;
    wire N__31698;
    wire N__31695;
    wire N__31692;
    wire N__31691;
    wire N__31688;
    wire N__31685;
    wire N__31680;
    wire N__31677;
    wire N__31674;
    wire N__31671;
    wire N__31668;
    wire N__31667;
    wire N__31666;
    wire N__31663;
    wire N__31660;
    wire N__31657;
    wire N__31650;
    wire N__31647;
    wire N__31644;
    wire N__31641;
    wire N__31640;
    wire N__31637;
    wire N__31634;
    wire N__31631;
    wire N__31628;
    wire N__31623;
    wire N__31620;
    wire N__31617;
    wire N__31614;
    wire N__31611;
    wire N__31610;
    wire N__31607;
    wire N__31606;
    wire N__31603;
    wire N__31600;
    wire N__31597;
    wire N__31594;
    wire N__31587;
    wire N__31584;
    wire N__31581;
    wire N__31578;
    wire N__31575;
    wire N__31572;
    wire N__31571;
    wire N__31568;
    wire N__31565;
    wire N__31562;
    wire N__31559;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31538;
    wire N__31535;
    wire N__31532;
    wire N__31531;
    wire N__31528;
    wire N__31525;
    wire N__31522;
    wire N__31515;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31503;
    wire N__31502;
    wire N__31499;
    wire N__31498;
    wire N__31495;
    wire N__31492;
    wire N__31489;
    wire N__31482;
    wire N__31479;
    wire N__31476;
    wire N__31473;
    wire N__31470;
    wire N__31467;
    wire N__31464;
    wire N__31463;
    wire N__31460;
    wire N__31457;
    wire N__31452;
    wire N__31449;
    wire N__31446;
    wire N__31443;
    wire N__31440;
    wire N__31437;
    wire N__31434;
    wire N__31431;
    wire N__31430;
    wire N__31427;
    wire N__31424;
    wire N__31421;
    wire N__31420;
    wire N__31417;
    wire N__31414;
    wire N__31411;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31395;
    wire N__31392;
    wire N__31389;
    wire N__31386;
    wire N__31383;
    wire N__31380;
    wire N__31377;
    wire N__31376;
    wire N__31371;
    wire N__31368;
    wire N__31365;
    wire N__31362;
    wire N__31359;
    wire N__31356;
    wire N__31355;
    wire N__31352;
    wire N__31349;
    wire N__31346;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31336;
    wire N__31333;
    wire N__31330;
    wire N__31323;
    wire N__31320;
    wire N__31317;
    wire N__31314;
    wire N__31313;
    wire N__31312;
    wire N__31309;
    wire N__31306;
    wire N__31303;
    wire N__31300;
    wire N__31297;
    wire N__31294;
    wire N__31291;
    wire N__31288;
    wire N__31285;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31269;
    wire N__31266;
    wire N__31263;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31251;
    wire N__31248;
    wire N__31245;
    wire N__31242;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31230;
    wire N__31227;
    wire N__31224;
    wire N__31221;
    wire N__31218;
    wire N__31217;
    wire N__31214;
    wire N__31211;
    wire N__31206;
    wire N__31203;
    wire N__31200;
    wire N__31199;
    wire N__31196;
    wire N__31193;
    wire N__31190;
    wire N__31187;
    wire N__31182;
    wire N__31181;
    wire N__31178;
    wire N__31175;
    wire N__31170;
    wire N__31167;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31155;
    wire N__31152;
    wire N__31149;
    wire N__31146;
    wire N__31143;
    wire N__31140;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31125;
    wire N__31122;
    wire N__31119;
    wire N__31116;
    wire N__31113;
    wire N__31110;
    wire N__31107;
    wire N__31104;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31089;
    wire N__31086;
    wire N__31083;
    wire N__31080;
    wire N__31077;
    wire N__31074;
    wire N__31071;
    wire N__31068;
    wire N__31065;
    wire N__31064;
    wire N__31063;
    wire N__31060;
    wire N__31057;
    wire N__31054;
    wire N__31047;
    wire N__31044;
    wire N__31041;
    wire N__31038;
    wire N__31035;
    wire N__31032;
    wire N__31029;
    wire N__31028;
    wire N__31027;
    wire N__31024;
    wire N__31021;
    wire N__31018;
    wire N__31011;
    wire N__31008;
    wire N__31005;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30992;
    wire N__30989;
    wire N__30986;
    wire N__30985;
    wire N__30982;
    wire N__30979;
    wire N__30976;
    wire N__30973;
    wire N__30968;
    wire N__30963;
    wire N__30962;
    wire N__30959;
    wire N__30956;
    wire N__30953;
    wire N__30952;
    wire N__30949;
    wire N__30946;
    wire N__30943;
    wire N__30936;
    wire N__30933;
    wire N__30930;
    wire N__30927;
    wire N__30924;
    wire N__30921;
    wire N__30918;
    wire N__30915;
    wire N__30912;
    wire N__30909;
    wire N__30906;
    wire N__30903;
    wire N__30900;
    wire N__30897;
    wire N__30894;
    wire N__30891;
    wire N__30890;
    wire N__30887;
    wire N__30884;
    wire N__30883;
    wire N__30878;
    wire N__30875;
    wire N__30870;
    wire N__30867;
    wire N__30864;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30852;
    wire N__30851;
    wire N__30848;
    wire N__30847;
    wire N__30844;
    wire N__30841;
    wire N__30838;
    wire N__30831;
    wire N__30828;
    wire N__30825;
    wire N__30822;
    wire N__30819;
    wire N__30816;
    wire N__30813;
    wire N__30812;
    wire N__30811;
    wire N__30808;
    wire N__30805;
    wire N__30802;
    wire N__30799;
    wire N__30796;
    wire N__30793;
    wire N__30786;
    wire N__30783;
    wire N__30780;
    wire N__30777;
    wire N__30774;
    wire N__30771;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30753;
    wire N__30750;
    wire N__30747;
    wire N__30744;
    wire N__30741;
    wire N__30738;
    wire N__30737;
    wire N__30734;
    wire N__30731;
    wire N__30730;
    wire N__30727;
    wire N__30724;
    wire N__30721;
    wire N__30716;
    wire N__30711;
    wire N__30708;
    wire N__30705;
    wire N__30702;
    wire N__30699;
    wire N__30696;
    wire N__30693;
    wire N__30692;
    wire N__30689;
    wire N__30686;
    wire N__30681;
    wire N__30678;
    wire N__30675;
    wire N__30672;
    wire N__30669;
    wire N__30666;
    wire N__30665;
    wire N__30662;
    wire N__30659;
    wire N__30658;
    wire N__30653;
    wire N__30650;
    wire N__30645;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30627;
    wire N__30624;
    wire N__30623;
    wire N__30620;
    wire N__30617;
    wire N__30614;
    wire N__30609;
    wire N__30608;
    wire N__30605;
    wire N__30602;
    wire N__30597;
    wire N__30594;
    wire N__30591;
    wire N__30588;
    wire N__30587;
    wire N__30584;
    wire N__30581;
    wire N__30580;
    wire N__30577;
    wire N__30574;
    wire N__30571;
    wire N__30564;
    wire N__30561;
    wire N__30560;
    wire N__30557;
    wire N__30554;
    wire N__30551;
    wire N__30548;
    wire N__30545;
    wire N__30544;
    wire N__30541;
    wire N__30538;
    wire N__30535;
    wire N__30528;
    wire N__30525;
    wire N__30522;
    wire N__30519;
    wire N__30516;
    wire N__30513;
    wire N__30510;
    wire N__30507;
    wire N__30506;
    wire N__30503;
    wire N__30500;
    wire N__30497;
    wire N__30492;
    wire N__30489;
    wire N__30488;
    wire N__30485;
    wire N__30484;
    wire N__30481;
    wire N__30478;
    wire N__30475;
    wire N__30468;
    wire N__30465;
    wire N__30462;
    wire N__30459;
    wire N__30456;
    wire N__30453;
    wire N__30450;
    wire N__30447;
    wire N__30444;
    wire N__30441;
    wire N__30438;
    wire N__30435;
    wire N__30432;
    wire N__30431;
    wire N__30428;
    wire N__30425;
    wire N__30422;
    wire N__30421;
    wire N__30418;
    wire N__30415;
    wire N__30412;
    wire N__30405;
    wire N__30402;
    wire N__30399;
    wire N__30396;
    wire N__30393;
    wire N__30390;
    wire N__30389;
    wire N__30386;
    wire N__30385;
    wire N__30382;
    wire N__30379;
    wire N__30376;
    wire N__30369;
    wire N__30368;
    wire N__30365;
    wire N__30362;
    wire N__30359;
    wire N__30356;
    wire N__30355;
    wire N__30352;
    wire N__30349;
    wire N__30346;
    wire N__30339;
    wire N__30336;
    wire N__30333;
    wire N__30330;
    wire N__30327;
    wire N__30324;
    wire N__30323;
    wire N__30320;
    wire N__30317;
    wire N__30314;
    wire N__30311;
    wire N__30310;
    wire N__30307;
    wire N__30304;
    wire N__30301;
    wire N__30294;
    wire N__30291;
    wire N__30290;
    wire N__30287;
    wire N__30286;
    wire N__30283;
    wire N__30280;
    wire N__30277;
    wire N__30270;
    wire N__30267;
    wire N__30264;
    wire N__30261;
    wire N__30258;
    wire N__30255;
    wire N__30252;
    wire N__30251;
    wire N__30248;
    wire N__30245;
    wire N__30242;
    wire N__30239;
    wire N__30238;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30222;
    wire N__30221;
    wire N__30220;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30203;
    wire N__30198;
    wire N__30195;
    wire N__30192;
    wire N__30189;
    wire N__30186;
    wire N__30183;
    wire N__30180;
    wire N__30179;
    wire N__30176;
    wire N__30173;
    wire N__30172;
    wire N__30169;
    wire N__30166;
    wire N__30163;
    wire N__30156;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30144;
    wire N__30141;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30130;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30118;
    wire N__30111;
    wire N__30108;
    wire N__30105;
    wire N__30102;
    wire N__30099;
    wire N__30096;
    wire N__30095;
    wire N__30092;
    wire N__30089;
    wire N__30086;
    wire N__30081;
    wire N__30078;
    wire N__30077;
    wire N__30074;
    wire N__30073;
    wire N__30070;
    wire N__30067;
    wire N__30064;
    wire N__30057;
    wire N__30054;
    wire N__30051;
    wire N__30048;
    wire N__30045;
    wire N__30042;
    wire N__30039;
    wire N__30038;
    wire N__30035;
    wire N__30032;
    wire N__30027;
    wire N__30024;
    wire N__30021;
    wire N__30018;
    wire N__30015;
    wire N__30012;
    wire N__30009;
    wire N__30008;
    wire N__30007;
    wire N__30004;
    wire N__30001;
    wire N__29998;
    wire N__29995;
    wire N__29992;
    wire N__29989;
    wire N__29984;
    wire N__29979;
    wire N__29978;
    wire N__29975;
    wire N__29972;
    wire N__29969;
    wire N__29966;
    wire N__29963;
    wire N__29958;
    wire N__29955;
    wire N__29954;
    wire N__29951;
    wire N__29948;
    wire N__29947;
    wire N__29944;
    wire N__29941;
    wire N__29938;
    wire N__29931;
    wire N__29928;
    wire N__29927;
    wire N__29926;
    wire N__29923;
    wire N__29920;
    wire N__29917;
    wire N__29914;
    wire N__29907;
    wire N__29904;
    wire N__29901;
    wire N__29898;
    wire N__29895;
    wire N__29892;
    wire N__29889;
    wire N__29888;
    wire N__29885;
    wire N__29884;
    wire N__29881;
    wire N__29878;
    wire N__29875;
    wire N__29872;
    wire N__29869;
    wire N__29866;
    wire N__29863;
    wire N__29856;
    wire N__29853;
    wire N__29852;
    wire N__29849;
    wire N__29848;
    wire N__29845;
    wire N__29842;
    wire N__29839;
    wire N__29832;
    wire N__29831;
    wire N__29828;
    wire N__29827;
    wire N__29824;
    wire N__29821;
    wire N__29818;
    wire N__29815;
    wire N__29810;
    wire N__29805;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29790;
    wire N__29787;
    wire N__29784;
    wire N__29781;
    wire N__29778;
    wire N__29775;
    wire N__29774;
    wire N__29771;
    wire N__29768;
    wire N__29767;
    wire N__29762;
    wire N__29759;
    wire N__29756;
    wire N__29751;
    wire N__29748;
    wire N__29745;
    wire N__29742;
    wire N__29739;
    wire N__29736;
    wire N__29733;
    wire N__29732;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29720;
    wire N__29715;
    wire N__29712;
    wire N__29709;
    wire N__29708;
    wire N__29705;
    wire N__29702;
    wire N__29701;
    wire N__29696;
    wire N__29693;
    wire N__29688;
    wire N__29685;
    wire N__29684;
    wire N__29683;
    wire N__29680;
    wire N__29677;
    wire N__29674;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29662;
    wire N__29659;
    wire N__29656;
    wire N__29649;
    wire N__29648;
    wire N__29645;
    wire N__29642;
    wire N__29639;
    wire N__29636;
    wire N__29635;
    wire N__29632;
    wire N__29629;
    wire N__29626;
    wire N__29623;
    wire N__29616;
    wire N__29613;
    wire N__29610;
    wire N__29607;
    wire N__29604;
    wire N__29601;
    wire N__29598;
    wire N__29595;
    wire N__29592;
    wire N__29591;
    wire N__29590;
    wire N__29587;
    wire N__29582;
    wire N__29579;
    wire N__29574;
    wire N__29571;
    wire N__29568;
    wire N__29565;
    wire N__29562;
    wire N__29561;
    wire N__29558;
    wire N__29555;
    wire N__29552;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29540;
    wire N__29537;
    wire N__29534;
    wire N__29533;
    wire N__29530;
    wire N__29527;
    wire N__29524;
    wire N__29521;
    wire N__29516;
    wire N__29511;
    wire N__29508;
    wire N__29505;
    wire N__29502;
    wire N__29501;
    wire N__29500;
    wire N__29497;
    wire N__29494;
    wire N__29491;
    wire N__29488;
    wire N__29483;
    wire N__29480;
    wire N__29475;
    wire N__29472;
    wire N__29469;
    wire N__29466;
    wire N__29463;
    wire N__29460;
    wire N__29457;
    wire N__29454;
    wire N__29453;
    wire N__29450;
    wire N__29447;
    wire N__29444;
    wire N__29439;
    wire N__29438;
    wire N__29435;
    wire N__29434;
    wire N__29431;
    wire N__29428;
    wire N__29425;
    wire N__29422;
    wire N__29419;
    wire N__29416;
    wire N__29413;
    wire N__29410;
    wire N__29407;
    wire N__29404;
    wire N__29401;
    wire N__29394;
    wire N__29391;
    wire N__29388;
    wire N__29387;
    wire N__29384;
    wire N__29383;
    wire N__29380;
    wire N__29377;
    wire N__29374;
    wire N__29371;
    wire N__29368;
    wire N__29365;
    wire N__29362;
    wire N__29357;
    wire N__29352;
    wire N__29349;
    wire N__29346;
    wire N__29343;
    wire N__29340;
    wire N__29337;
    wire N__29336;
    wire N__29333;
    wire N__29330;
    wire N__29329;
    wire N__29326;
    wire N__29323;
    wire N__29320;
    wire N__29313;
    wire N__29310;
    wire N__29307;
    wire N__29304;
    wire N__29301;
    wire N__29300;
    wire N__29297;
    wire N__29294;
    wire N__29291;
    wire N__29288;
    wire N__29283;
    wire N__29280;
    wire N__29277;
    wire N__29274;
    wire N__29271;
    wire N__29268;
    wire N__29265;
    wire N__29262;
    wire N__29259;
    wire N__29256;
    wire N__29253;
    wire N__29252;
    wire N__29249;
    wire N__29246;
    wire N__29243;
    wire N__29240;
    wire N__29239;
    wire N__29236;
    wire N__29233;
    wire N__29230;
    wire N__29227;
    wire N__29220;
    wire N__29217;
    wire N__29214;
    wire N__29211;
    wire N__29208;
    wire N__29205;
    wire N__29202;
    wire N__29199;
    wire N__29196;
    wire N__29195;
    wire N__29192;
    wire N__29189;
    wire N__29186;
    wire N__29183;
    wire N__29182;
    wire N__29179;
    wire N__29176;
    wire N__29173;
    wire N__29170;
    wire N__29163;
    wire N__29160;
    wire N__29157;
    wire N__29154;
    wire N__29151;
    wire N__29148;
    wire N__29145;
    wire N__29142;
    wire N__29139;
    wire N__29136;
    wire N__29133;
    wire N__29130;
    wire N__29127;
    wire N__29124;
    wire N__29123;
    wire N__29120;
    wire N__29117;
    wire N__29114;
    wire N__29111;
    wire N__29108;
    wire N__29105;
    wire N__29104;
    wire N__29101;
    wire N__29098;
    wire N__29095;
    wire N__29088;
    wire N__29085;
    wire N__29082;
    wire N__29079;
    wire N__29076;
    wire N__29073;
    wire N__29070;
    wire N__29069;
    wire N__29066;
    wire N__29063;
    wire N__29060;
    wire N__29059;
    wire N__29056;
    wire N__29053;
    wire N__29050;
    wire N__29045;
    wire N__29040;
    wire N__29037;
    wire N__29034;
    wire N__29031;
    wire N__29028;
    wire N__29025;
    wire N__29024;
    wire N__29021;
    wire N__29018;
    wire N__29017;
    wire N__29014;
    wire N__29011;
    wire N__29008;
    wire N__29005;
    wire N__29002;
    wire N__28999;
    wire N__28992;
    wire N__28989;
    wire N__28986;
    wire N__28983;
    wire N__28980;
    wire N__28979;
    wire N__28976;
    wire N__28973;
    wire N__28972;
    wire N__28969;
    wire N__28966;
    wire N__28963;
    wire N__28960;
    wire N__28957;
    wire N__28954;
    wire N__28947;
    wire N__28944;
    wire N__28941;
    wire N__28938;
    wire N__28935;
    wire N__28932;
    wire N__28929;
    wire N__28926;
    wire N__28923;
    wire N__28922;
    wire N__28919;
    wire N__28916;
    wire N__28913;
    wire N__28910;
    wire N__28907;
    wire N__28904;
    wire N__28899;
    wire N__28896;
    wire N__28895;
    wire N__28892;
    wire N__28891;
    wire N__28888;
    wire N__28885;
    wire N__28882;
    wire N__28879;
    wire N__28872;
    wire N__28869;
    wire N__28866;
    wire N__28863;
    wire N__28860;
    wire N__28859;
    wire N__28856;
    wire N__28853;
    wire N__28850;
    wire N__28849;
    wire N__28846;
    wire N__28843;
    wire N__28840;
    wire N__28833;
    wire N__28832;
    wire N__28831;
    wire N__28828;
    wire N__28825;
    wire N__28822;
    wire N__28819;
    wire N__28816;
    wire N__28813;
    wire N__28808;
    wire N__28803;
    wire N__28800;
    wire N__28797;
    wire N__28794;
    wire N__28791;
    wire N__28790;
    wire N__28787;
    wire N__28784;
    wire N__28781;
    wire N__28778;
    wire N__28775;
    wire N__28774;
    wire N__28769;
    wire N__28766;
    wire N__28761;
    wire N__28758;
    wire N__28755;
    wire N__28752;
    wire N__28749;
    wire N__28746;
    wire N__28743;
    wire N__28740;
    wire N__28737;
    wire N__28736;
    wire N__28733;
    wire N__28730;
    wire N__28727;
    wire N__28724;
    wire N__28721;
    wire N__28720;
    wire N__28717;
    wire N__28714;
    wire N__28711;
    wire N__28704;
    wire N__28701;
    wire N__28698;
    wire N__28695;
    wire N__28692;
    wire N__28689;
    wire N__28688;
    wire N__28685;
    wire N__28682;
    wire N__28681;
    wire N__28678;
    wire N__28675;
    wire N__28672;
    wire N__28669;
    wire N__28664;
    wire N__28659;
    wire N__28656;
    wire N__28653;
    wire N__28650;
    wire N__28647;
    wire N__28644;
    wire N__28641;
    wire N__28638;
    wire N__28637;
    wire N__28634;
    wire N__28631;
    wire N__28628;
    wire N__28625;
    wire N__28622;
    wire N__28619;
    wire N__28614;
    wire N__28611;
    wire N__28608;
    wire N__28607;
    wire N__28604;
    wire N__28601;
    wire N__28600;
    wire N__28597;
    wire N__28594;
    wire N__28591;
    wire N__28584;
    wire N__28581;
    wire N__28578;
    wire N__28575;
    wire N__28574;
    wire N__28573;
    wire N__28570;
    wire N__28567;
    wire N__28564;
    wire N__28561;
    wire N__28558;
    wire N__28555;
    wire N__28548;
    wire N__28545;
    wire N__28542;
    wire N__28539;
    wire N__28536;
    wire N__28535;
    wire N__28532;
    wire N__28531;
    wire N__28528;
    wire N__28525;
    wire N__28522;
    wire N__28519;
    wire N__28516;
    wire N__28513;
    wire N__28506;
    wire N__28503;
    wire N__28500;
    wire N__28499;
    wire N__28496;
    wire N__28493;
    wire N__28488;
    wire N__28485;
    wire N__28484;
    wire N__28483;
    wire N__28480;
    wire N__28477;
    wire N__28474;
    wire N__28471;
    wire N__28468;
    wire N__28461;
    wire N__28458;
    wire N__28455;
    wire N__28452;
    wire N__28451;
    wire N__28450;
    wire N__28447;
    wire N__28444;
    wire N__28441;
    wire N__28438;
    wire N__28435;
    wire N__28432;
    wire N__28425;
    wire N__28422;
    wire N__28421;
    wire N__28420;
    wire N__28417;
    wire N__28412;
    wire N__28407;
    wire N__28404;
    wire N__28401;
    wire N__28398;
    wire N__28395;
    wire N__28392;
    wire N__28389;
    wire N__28386;
    wire N__28385;
    wire N__28384;
    wire N__28381;
    wire N__28376;
    wire N__28373;
    wire N__28370;
    wire N__28367;
    wire N__28364;
    wire N__28361;
    wire N__28356;
    wire N__28353;
    wire N__28350;
    wire N__28347;
    wire N__28344;
    wire N__28341;
    wire N__28340;
    wire N__28337;
    wire N__28336;
    wire N__28333;
    wire N__28330;
    wire N__28327;
    wire N__28324;
    wire N__28319;
    wire N__28314;
    wire N__28311;
    wire N__28308;
    wire N__28305;
    wire N__28304;
    wire N__28301;
    wire N__28298;
    wire N__28295;
    wire N__28292;
    wire N__28289;
    wire N__28288;
    wire N__28285;
    wire N__28282;
    wire N__28279;
    wire N__28272;
    wire N__28269;
    wire N__28266;
    wire N__28263;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28251;
    wire N__28248;
    wire N__28247;
    wire N__28246;
    wire N__28243;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28224;
    wire N__28223;
    wire N__28220;
    wire N__28217;
    wire N__28214;
    wire N__28209;
    wire N__28208;
    wire N__28205;
    wire N__28202;
    wire N__28197;
    wire N__28196;
    wire N__28193;
    wire N__28190;
    wire N__28185;
    wire N__28182;
    wire N__28179;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28164;
    wire N__28161;
    wire N__28158;
    wire N__28155;
    wire N__28152;
    wire N__28151;
    wire N__28150;
    wire N__28147;
    wire N__28142;
    wire N__28137;
    wire N__28134;
    wire N__28131;
    wire N__28128;
    wire N__28127;
    wire N__28124;
    wire N__28121;
    wire N__28118;
    wire N__28115;
    wire N__28110;
    wire N__28107;
    wire N__28104;
    wire N__28101;
    wire N__28098;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28086;
    wire N__28083;
    wire N__28080;
    wire N__28077;
    wire N__28076;
    wire N__28075;
    wire N__28072;
    wire N__28069;
    wire N__28066;
    wire N__28059;
    wire N__28058;
    wire N__28057;
    wire N__28054;
    wire N__28051;
    wire N__28048;
    wire N__28041;
    wire N__28040;
    wire N__28037;
    wire N__28034;
    wire N__28031;
    wire N__28026;
    wire N__28023;
    wire N__28020;
    wire N__28017;
    wire N__28014;
    wire N__28011;
    wire N__28008;
    wire N__28007;
    wire N__28004;
    wire N__28001;
    wire N__27998;
    wire N__27995;
    wire N__27990;
    wire N__27987;
    wire N__27984;
    wire N__27981;
    wire N__27978;
    wire N__27975;
    wire N__27972;
    wire N__27969;
    wire N__27968;
    wire N__27967;
    wire N__27964;
    wire N__27961;
    wire N__27958;
    wire N__27955;
    wire N__27952;
    wire N__27949;
    wire N__27944;
    wire N__27939;
    wire N__27936;
    wire N__27933;
    wire N__27930;
    wire N__27927;
    wire N__27924;
    wire N__27921;
    wire N__27918;
    wire N__27915;
    wire N__27914;
    wire N__27913;
    wire N__27910;
    wire N__27907;
    wire N__27904;
    wire N__27897;
    wire N__27894;
    wire N__27891;
    wire N__27888;
    wire N__27885;
    wire N__27882;
    wire N__27881;
    wire N__27878;
    wire N__27877;
    wire N__27874;
    wire N__27871;
    wire N__27868;
    wire N__27863;
    wire N__27860;
    wire N__27857;
    wire N__27854;
    wire N__27849;
    wire N__27846;
    wire N__27843;
    wire N__27842;
    wire N__27839;
    wire N__27836;
    wire N__27831;
    wire N__27828;
    wire N__27825;
    wire N__27822;
    wire N__27819;
    wire N__27816;
    wire N__27813;
    wire N__27810;
    wire N__27809;
    wire N__27806;
    wire N__27803;
    wire N__27802;
    wire N__27799;
    wire N__27796;
    wire N__27793;
    wire N__27786;
    wire N__27783;
    wire N__27780;
    wire N__27777;
    wire N__27774;
    wire N__27771;
    wire N__27768;
    wire N__27765;
    wire N__27764;
    wire N__27761;
    wire N__27758;
    wire N__27755;
    wire N__27752;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27742;
    wire N__27735;
    wire N__27734;
    wire N__27733;
    wire N__27730;
    wire N__27727;
    wire N__27724;
    wire N__27721;
    wire N__27718;
    wire N__27715;
    wire N__27712;
    wire N__27705;
    wire N__27702;
    wire N__27699;
    wire N__27696;
    wire N__27693;
    wire N__27690;
    wire N__27687;
    wire N__27684;
    wire N__27683;
    wire N__27680;
    wire N__27677;
    wire N__27676;
    wire N__27671;
    wire N__27668;
    wire N__27663;
    wire N__27660;
    wire N__27657;
    wire N__27654;
    wire N__27651;
    wire N__27648;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27636;
    wire N__27633;
    wire N__27630;
    wire N__27627;
    wire N__27624;
    wire N__27621;
    wire N__27618;
    wire N__27615;
    wire N__27612;
    wire N__27609;
    wire N__27606;
    wire N__27603;
    wire N__27600;
    wire N__27597;
    wire N__27594;
    wire N__27591;
    wire N__27588;
    wire N__27587;
    wire N__27584;
    wire N__27581;
    wire N__27578;
    wire N__27575;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27565;
    wire N__27558;
    wire N__27555;
    wire N__27552;
    wire N__27551;
    wire N__27548;
    wire N__27545;
    wire N__27544;
    wire N__27541;
    wire N__27538;
    wire N__27535;
    wire N__27528;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27516;
    wire N__27513;
    wire N__27510;
    wire N__27507;
    wire N__27504;
    wire N__27501;
    wire N__27498;
    wire N__27495;
    wire N__27494;
    wire N__27491;
    wire N__27488;
    wire N__27487;
    wire N__27482;
    wire N__27479;
    wire N__27474;
    wire N__27471;
    wire N__27468;
    wire N__27465;
    wire N__27462;
    wire N__27461;
    wire N__27458;
    wire N__27457;
    wire N__27454;
    wire N__27451;
    wire N__27448;
    wire N__27445;
    wire N__27440;
    wire N__27435;
    wire N__27432;
    wire N__27431;
    wire N__27428;
    wire N__27425;
    wire N__27422;
    wire N__27419;
    wire N__27418;
    wire N__27413;
    wire N__27410;
    wire N__27405;
    wire N__27404;
    wire N__27401;
    wire N__27398;
    wire N__27395;
    wire N__27394;
    wire N__27391;
    wire N__27388;
    wire N__27385;
    wire N__27382;
    wire N__27377;
    wire N__27372;
    wire N__27369;
    wire N__27366;
    wire N__27365;
    wire N__27362;
    wire N__27359;
    wire N__27356;
    wire N__27353;
    wire N__27348;
    wire N__27347;
    wire N__27342;
    wire N__27341;
    wire N__27338;
    wire N__27335;
    wire N__27330;
    wire N__27327;
    wire N__27324;
    wire N__27323;
    wire N__27318;
    wire N__27315;
    wire N__27312;
    wire N__27311;
    wire N__27308;
    wire N__27305;
    wire N__27302;
    wire N__27299;
    wire N__27294;
    wire N__27291;
    wire N__27288;
    wire N__27285;
    wire N__27282;
    wire N__27279;
    wire N__27278;
    wire N__27277;
    wire N__27274;
    wire N__27271;
    wire N__27268;
    wire N__27263;
    wire N__27260;
    wire N__27257;
    wire N__27252;
    wire N__27249;
    wire N__27246;
    wire N__27243;
    wire N__27240;
    wire N__27239;
    wire N__27236;
    wire N__27235;
    wire N__27232;
    wire N__27229;
    wire N__27226;
    wire N__27223;
    wire N__27216;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27200;
    wire N__27197;
    wire N__27196;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27180;
    wire N__27177;
    wire N__27174;
    wire N__27171;
    wire N__27168;
    wire N__27167;
    wire N__27166;
    wire N__27163;
    wire N__27160;
    wire N__27157;
    wire N__27154;
    wire N__27151;
    wire N__27148;
    wire N__27145;
    wire N__27142;
    wire N__27139;
    wire N__27134;
    wire N__27129;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27119;
    wire N__27118;
    wire N__27115;
    wire N__27112;
    wire N__27109;
    wire N__27106;
    wire N__27103;
    wire N__27096;
    wire N__27093;
    wire N__27092;
    wire N__27091;
    wire N__27088;
    wire N__27083;
    wire N__27078;
    wire N__27075;
    wire N__27072;
    wire N__27071;
    wire N__27068;
    wire N__27065;
    wire N__27064;
    wire N__27059;
    wire N__27056;
    wire N__27053;
    wire N__27050;
    wire N__27045;
    wire N__27042;
    wire N__27041;
    wire N__27038;
    wire N__27035;
    wire N__27030;
    wire N__27027;
    wire N__27026;
    wire N__27023;
    wire N__27020;
    wire N__27017;
    wire N__27014;
    wire N__27011;
    wire N__27008;
    wire N__27003;
    wire N__27002;
    wire N__26999;
    wire N__26996;
    wire N__26993;
    wire N__26990;
    wire N__26987;
    wire N__26982;
    wire N__26979;
    wire N__26976;
    wire N__26973;
    wire N__26972;
    wire N__26971;
    wire N__26968;
    wire N__26965;
    wire N__26962;
    wire N__26957;
    wire N__26952;
    wire N__26949;
    wire N__26946;
    wire N__26943;
    wire N__26940;
    wire N__26937;
    wire N__26936;
    wire N__26935;
    wire N__26932;
    wire N__26927;
    wire N__26922;
    wire N__26919;
    wire N__26916;
    wire N__26913;
    wire N__26910;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26898;
    wire N__26895;
    wire N__26894;
    wire N__26893;
    wire N__26890;
    wire N__26885;
    wire N__26880;
    wire N__26877;
    wire N__26874;
    wire N__26871;
    wire N__26868;
    wire N__26865;
    wire N__26862;
    wire N__26859;
    wire N__26856;
    wire N__26853;
    wire N__26850;
    wire N__26847;
    wire N__26844;
    wire N__26843;
    wire N__26840;
    wire N__26837;
    wire N__26834;
    wire N__26833;
    wire N__26830;
    wire N__26827;
    wire N__26824;
    wire N__26817;
    wire N__26814;
    wire N__26813;
    wire N__26810;
    wire N__26807;
    wire N__26802;
    wire N__26799;
    wire N__26796;
    wire N__26795;
    wire N__26792;
    wire N__26789;
    wire N__26786;
    wire N__26781;
    wire N__26778;
    wire N__26775;
    wire N__26774;
    wire N__26773;
    wire N__26770;
    wire N__26767;
    wire N__26764;
    wire N__26757;
    wire N__26754;
    wire N__26751;
    wire N__26750;
    wire N__26747;
    wire N__26744;
    wire N__26741;
    wire N__26740;
    wire N__26737;
    wire N__26734;
    wire N__26731;
    wire N__26728;
    wire N__26723;
    wire N__26720;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26700;
    wire N__26699;
    wire N__26698;
    wire N__26695;
    wire N__26692;
    wire N__26689;
    wire N__26682;
    wire N__26679;
    wire N__26676;
    wire N__26675;
    wire N__26674;
    wire N__26671;
    wire N__26668;
    wire N__26665;
    wire N__26658;
    wire N__26655;
    wire N__26654;
    wire N__26653;
    wire N__26650;
    wire N__26647;
    wire N__26644;
    wire N__26637;
    wire N__26634;
    wire N__26631;
    wire N__26628;
    wire N__26625;
    wire N__26622;
    wire N__26619;
    wire N__26618;
    wire N__26615;
    wire N__26614;
    wire N__26611;
    wire N__26608;
    wire N__26605;
    wire N__26598;
    wire N__26595;
    wire N__26592;
    wire N__26589;
    wire N__26586;
    wire N__26583;
    wire N__26580;
    wire N__26577;
    wire N__26574;
    wire N__26573;
    wire N__26572;
    wire N__26569;
    wire N__26566;
    wire N__26563;
    wire N__26560;
    wire N__26557;
    wire N__26552;
    wire N__26549;
    wire N__26544;
    wire N__26541;
    wire N__26540;
    wire N__26537;
    wire N__26534;
    wire N__26533;
    wire N__26530;
    wire N__26525;
    wire N__26522;
    wire N__26517;
    wire N__26514;
    wire N__26511;
    wire N__26508;
    wire N__26505;
    wire N__26504;
    wire N__26501;
    wire N__26500;
    wire N__26497;
    wire N__26494;
    wire N__26491;
    wire N__26488;
    wire N__26485;
    wire N__26478;
    wire N__26475;
    wire N__26472;
    wire N__26471;
    wire N__26468;
    wire N__26465;
    wire N__26464;
    wire N__26461;
    wire N__26458;
    wire N__26455;
    wire N__26448;
    wire N__26447;
    wire N__26444;
    wire N__26441;
    wire N__26438;
    wire N__26435;
    wire N__26434;
    wire N__26429;
    wire N__26426;
    wire N__26421;
    wire N__26418;
    wire N__26415;
    wire N__26414;
    wire N__26411;
    wire N__26408;
    wire N__26403;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26395;
    wire N__26392;
    wire N__26389;
    wire N__26386;
    wire N__26383;
    wire N__26380;
    wire N__26377;
    wire N__26370;
    wire N__26367;
    wire N__26366;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26337;
    wire N__26334;
    wire N__26333;
    wire N__26332;
    wire N__26329;
    wire N__26324;
    wire N__26319;
    wire N__26316;
    wire N__26313;
    wire N__26310;
    wire N__26307;
    wire N__26304;
    wire N__26301;
    wire N__26298;
    wire N__26295;
    wire N__26292;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26281;
    wire N__26278;
    wire N__26275;
    wire N__26272;
    wire N__26265;
    wire N__26262;
    wire N__26261;
    wire N__26258;
    wire N__26255;
    wire N__26252;
    wire N__26247;
    wire N__26244;
    wire N__26241;
    wire N__26238;
    wire N__26235;
    wire N__26232;
    wire N__26231;
    wire N__26230;
    wire N__26227;
    wire N__26224;
    wire N__26221;
    wire N__26218;
    wire N__26215;
    wire N__26208;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26198;
    wire N__26195;
    wire N__26192;
    wire N__26191;
    wire N__26188;
    wire N__26185;
    wire N__26182;
    wire N__26175;
    wire N__26172;
    wire N__26169;
    wire N__26168;
    wire N__26165;
    wire N__26164;
    wire N__26161;
    wire N__26158;
    wire N__26155;
    wire N__26148;
    wire N__26145;
    wire N__26142;
    wire N__26139;
    wire N__26136;
    wire N__26135;
    wire N__26134;
    wire N__26131;
    wire N__26126;
    wire N__26123;
    wire N__26118;
    wire N__26115;
    wire N__26112;
    wire N__26109;
    wire N__26106;
    wire N__26103;
    wire N__26102;
    wire N__26099;
    wire N__26098;
    wire N__26095;
    wire N__26092;
    wire N__26089;
    wire N__26082;
    wire N__26079;
    wire N__26076;
    wire N__26073;
    wire N__26070;
    wire N__26067;
    wire N__26064;
    wire N__26061;
    wire N__26058;
    wire N__26055;
    wire N__26052;
    wire N__26049;
    wire N__26046;
    wire N__26043;
    wire N__26040;
    wire N__26037;
    wire N__26034;
    wire N__26033;
    wire N__26030;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26018;
    wire N__26017;
    wire N__26014;
    wire N__26011;
    wire N__26008;
    wire N__26003;
    wire N__25998;
    wire N__25997;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25985;
    wire N__25982;
    wire N__25979;
    wire N__25974;
    wire N__25971;
    wire N__25968;
    wire N__25965;
    wire N__25964;
    wire N__25963;
    wire N__25960;
    wire N__25957;
    wire N__25954;
    wire N__25951;
    wire N__25948;
    wire N__25945;
    wire N__25942;
    wire N__25935;
    wire N__25932;
    wire N__25929;
    wire N__25926;
    wire N__25923;
    wire N__25920;
    wire N__25917;
    wire N__25914;
    wire N__25911;
    wire N__25908;
    wire N__25905;
    wire N__25904;
    wire N__25901;
    wire N__25898;
    wire N__25895;
    wire N__25894;
    wire N__25891;
    wire N__25888;
    wire N__25885;
    wire N__25882;
    wire N__25875;
    wire N__25874;
    wire N__25871;
    wire N__25868;
    wire N__25865;
    wire N__25864;
    wire N__25861;
    wire N__25858;
    wire N__25855;
    wire N__25848;
    wire N__25845;
    wire N__25842;
    wire N__25839;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25827;
    wire N__25824;
    wire N__25821;
    wire N__25818;
    wire N__25815;
    wire N__25812;
    wire N__25809;
    wire N__25806;
    wire N__25805;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25788;
    wire N__25785;
    wire N__25782;
    wire N__25779;
    wire N__25778;
    wire N__25775;
    wire N__25774;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25758;
    wire N__25755;
    wire N__25752;
    wire N__25749;
    wire N__25746;
    wire N__25743;
    wire N__25740;
    wire N__25737;
    wire N__25734;
    wire N__25731;
    wire N__25728;
    wire N__25727;
    wire N__25724;
    wire N__25723;
    wire N__25720;
    wire N__25717;
    wire N__25714;
    wire N__25707;
    wire N__25704;
    wire N__25701;
    wire N__25698;
    wire N__25695;
    wire N__25692;
    wire N__25689;
    wire N__25688;
    wire N__25685;
    wire N__25682;
    wire N__25677;
    wire N__25674;
    wire N__25671;
    wire N__25668;
    wire N__25665;
    wire N__25662;
    wire N__25659;
    wire N__25656;
    wire N__25653;
    wire N__25652;
    wire N__25649;
    wire N__25646;
    wire N__25643;
    wire N__25640;
    wire N__25637;
    wire N__25636;
    wire N__25631;
    wire N__25628;
    wire N__25623;
    wire N__25622;
    wire N__25619;
    wire N__25618;
    wire N__25615;
    wire N__25612;
    wire N__25609;
    wire N__25602;
    wire N__25599;
    wire N__25596;
    wire N__25593;
    wire N__25590;
    wire N__25587;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25575;
    wire N__25574;
    wire N__25571;
    wire N__25568;
    wire N__25563;
    wire N__25560;
    wire N__25557;
    wire N__25554;
    wire N__25551;
    wire N__25548;
    wire N__25545;
    wire N__25542;
    wire N__25539;
    wire N__25536;
    wire N__25533;
    wire N__25530;
    wire N__25529;
    wire N__25526;
    wire N__25523;
    wire N__25518;
    wire N__25515;
    wire N__25512;
    wire N__25509;
    wire N__25506;
    wire N__25503;
    wire N__25500;
    wire N__25497;
    wire N__25494;
    wire N__25491;
    wire N__25490;
    wire N__25487;
    wire N__25486;
    wire N__25483;
    wire N__25480;
    wire N__25477;
    wire N__25470;
    wire N__25467;
    wire N__25464;
    wire N__25461;
    wire N__25458;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25440;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25428;
    wire N__25425;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25413;
    wire N__25410;
    wire N__25407;
    wire N__25404;
    wire N__25401;
    wire N__25400;
    wire N__25397;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25377;
    wire N__25376;
    wire N__25373;
    wire N__25370;
    wire N__25369;
    wire N__25366;
    wire N__25363;
    wire N__25360;
    wire N__25353;
    wire N__25350;
    wire N__25349;
    wire N__25346;
    wire N__25343;
    wire N__25342;
    wire N__25339;
    wire N__25336;
    wire N__25333;
    wire N__25326;
    wire N__25323;
    wire N__25320;
    wire N__25317;
    wire N__25314;
    wire N__25311;
    wire N__25308;
    wire N__25305;
    wire N__25302;
    wire N__25299;
    wire N__25296;
    wire N__25293;
    wire N__25290;
    wire N__25287;
    wire N__25284;
    wire N__25281;
    wire N__25278;
    wire N__25275;
    wire N__25272;
    wire N__25271;
    wire N__25268;
    wire N__25265;
    wire N__25262;
    wire N__25259;
    wire N__25254;
    wire N__25251;
    wire N__25248;
    wire N__25245;
    wire N__25242;
    wire N__25239;
    wire N__25236;
    wire N__25235;
    wire N__25232;
    wire N__25231;
    wire N__25228;
    wire N__25225;
    wire N__25222;
    wire N__25219;
    wire N__25212;
    wire N__25209;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25201;
    wire N__25198;
    wire N__25195;
    wire N__25192;
    wire N__25185;
    wire N__25182;
    wire N__25179;
    wire N__25178;
    wire N__25177;
    wire N__25174;
    wire N__25171;
    wire N__25168;
    wire N__25165;
    wire N__25162;
    wire N__25159;
    wire N__25152;
    wire N__25151;
    wire N__25150;
    wire N__25147;
    wire N__25142;
    wire N__25139;
    wire N__25136;
    wire N__25133;
    wire N__25128;
    wire N__25125;
    wire N__25122;
    wire N__25119;
    wire N__25116;
    wire N__25113;
    wire N__25110;
    wire N__25107;
    wire N__25104;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25092;
    wire N__25089;
    wire N__25086;
    wire N__25083;
    wire N__25080;
    wire N__25077;
    wire N__25074;
    wire N__25071;
    wire N__25068;
    wire N__25065;
    wire N__25062;
    wire N__25059;
    wire N__25056;
    wire N__25053;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25032;
    wire N__25029;
    wire N__25026;
    wire N__25023;
    wire N__25020;
    wire N__25017;
    wire N__25014;
    wire N__25011;
    wire N__25010;
    wire N__25007;
    wire N__25006;
    wire N__25003;
    wire N__25000;
    wire N__24997;
    wire N__24990;
    wire N__24987;
    wire N__24984;
    wire N__24981;
    wire N__24978;
    wire N__24977;
    wire N__24974;
    wire N__24971;
    wire N__24968;
    wire N__24965;
    wire N__24962;
    wire N__24959;
    wire N__24954;
    wire N__24951;
    wire N__24948;
    wire N__24945;
    wire N__24942;
    wire N__24939;
    wire N__24936;
    wire N__24935;
    wire N__24934;
    wire N__24931;
    wire N__24928;
    wire N__24925;
    wire N__24922;
    wire N__24919;
    wire N__24912;
    wire N__24909;
    wire N__24906;
    wire N__24903;
    wire N__24900;
    wire N__24897;
    wire N__24894;
    wire N__24891;
    wire N__24888;
    wire N__24885;
    wire N__24884;
    wire N__24881;
    wire N__24880;
    wire N__24877;
    wire N__24874;
    wire N__24871;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24831;
    wire N__24830;
    wire N__24827;
    wire N__24824;
    wire N__24821;
    wire N__24818;
    wire N__24813;
    wire N__24810;
    wire N__24807;
    wire N__24804;
    wire N__24801;
    wire N__24798;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24788;
    wire N__24785;
    wire N__24782;
    wire N__24779;
    wire N__24778;
    wire N__24775;
    wire N__24772;
    wire N__24769;
    wire N__24762;
    wire N__24759;
    wire N__24756;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24736;
    wire N__24731;
    wire N__24728;
    wire N__24723;
    wire N__24720;
    wire N__24717;
    wire N__24714;
    wire N__24711;
    wire N__24708;
    wire N__24707;
    wire N__24704;
    wire N__24701;
    wire N__24698;
    wire N__24695;
    wire N__24692;
    wire N__24687;
    wire N__24684;
    wire N__24681;
    wire N__24678;
    wire N__24675;
    wire N__24672;
    wire N__24669;
    wire N__24666;
    wire N__24663;
    wire N__24660;
    wire N__24657;
    wire N__24654;
    wire N__24651;
    wire N__24648;
    wire N__24645;
    wire N__24642;
    wire N__24639;
    wire N__24636;
    wire N__24633;
    wire N__24630;
    wire N__24627;
    wire N__24624;
    wire N__24621;
    wire N__24618;
    wire N__24617;
    wire N__24616;
    wire N__24613;
    wire N__24608;
    wire N__24603;
    wire N__24600;
    wire N__24597;
    wire N__24594;
    wire N__24591;
    wire N__24588;
    wire N__24585;
    wire N__24584;
    wire N__24581;
    wire N__24578;
    wire N__24577;
    wire N__24574;
    wire N__24571;
    wire N__24568;
    wire N__24561;
    wire N__24558;
    wire N__24555;
    wire N__24552;
    wire N__24549;
    wire N__24546;
    wire N__24543;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24535;
    wire N__24532;
    wire N__24529;
    wire N__24526;
    wire N__24519;
    wire N__24516;
    wire N__24513;
    wire N__24510;
    wire N__24507;
    wire N__24504;
    wire N__24501;
    wire N__24498;
    wire N__24495;
    wire N__24492;
    wire N__24489;
    wire N__24486;
    wire N__24483;
    wire N__24480;
    wire N__24477;
    wire N__24474;
    wire N__24471;
    wire N__24468;
    wire N__24467;
    wire N__24464;
    wire N__24463;
    wire N__24460;
    wire N__24457;
    wire N__24454;
    wire N__24451;
    wire N__24444;
    wire N__24441;
    wire N__24438;
    wire N__24435;
    wire N__24432;
    wire N__24429;
    wire N__24426;
    wire N__24423;
    wire N__24420;
    wire N__24417;
    wire N__24416;
    wire N__24415;
    wire N__24412;
    wire N__24409;
    wire N__24406;
    wire N__24403;
    wire N__24398;
    wire N__24393;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24381;
    wire N__24378;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24368;
    wire N__24365;
    wire N__24362;
    wire N__24359;
    wire N__24356;
    wire N__24353;
    wire N__24352;
    wire N__24349;
    wire N__24346;
    wire N__24343;
    wire N__24336;
    wire N__24333;
    wire N__24330;
    wire N__24327;
    wire N__24324;
    wire N__24321;
    wire N__24318;
    wire N__24315;
    wire N__24312;
    wire N__24309;
    wire N__24308;
    wire N__24307;
    wire N__24304;
    wire N__24299;
    wire N__24294;
    wire N__24291;
    wire N__24288;
    wire N__24285;
    wire N__24282;
    wire N__24279;
    wire N__24278;
    wire N__24277;
    wire N__24274;
    wire N__24271;
    wire N__24268;
    wire N__24265;
    wire N__24262;
    wire N__24259;
    wire N__24256;
    wire N__24253;
    wire N__24246;
    wire N__24243;
    wire N__24240;
    wire N__24237;
    wire N__24234;
    wire N__24231;
    wire N__24228;
    wire N__24227;
    wire N__24224;
    wire N__24221;
    wire N__24220;
    wire N__24217;
    wire N__24214;
    wire N__24211;
    wire N__24204;
    wire N__24201;
    wire N__24198;
    wire N__24195;
    wire N__24192;
    wire N__24189;
    wire N__24186;
    wire N__24183;
    wire N__24180;
    wire N__24177;
    wire N__24174;
    wire N__24171;
    wire N__24168;
    wire N__24165;
    wire N__24162;
    wire N__24159;
    wire N__24158;
    wire N__24157;
    wire N__24154;
    wire N__24149;
    wire N__24144;
    wire N__24141;
    wire N__24138;
    wire N__24135;
    wire N__24132;
    wire N__24129;
    wire N__24128;
    wire N__24125;
    wire N__24124;
    wire N__24121;
    wire N__24116;
    wire N__24113;
    wire N__24110;
    wire N__24107;
    wire N__24102;
    wire N__24099;
    wire N__24096;
    wire N__24093;
    wire N__24092;
    wire N__24091;
    wire N__24088;
    wire N__24083;
    wire N__24078;
    wire N__24075;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24065;
    wire N__24062;
    wire N__24059;
    wire N__24054;
    wire N__24051;
    wire N__24048;
    wire N__24045;
    wire N__24042;
    wire N__24039;
    wire N__24036;
    wire N__24035;
    wire N__24032;
    wire N__24029;
    wire N__24026;
    wire N__24021;
    wire N__24018;
    wire N__24015;
    wire N__24012;
    wire N__24009;
    wire N__24006;
    wire N__24003;
    wire N__24000;
    wire N__23997;
    wire N__23994;
    wire N__23991;
    wire N__23990;
    wire N__23987;
    wire N__23984;
    wire N__23983;
    wire N__23980;
    wire N__23977;
    wire N__23974;
    wire N__23967;
    wire N__23964;
    wire N__23961;
    wire N__23958;
    wire N__23955;
    wire N__23952;
    wire N__23949;
    wire N__23946;
    wire N__23945;
    wire N__23942;
    wire N__23939;
    wire N__23934;
    wire N__23931;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23919;
    wire N__23916;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23906;
    wire N__23905;
    wire N__23902;
    wire N__23899;
    wire N__23896;
    wire N__23889;
    wire N__23886;
    wire N__23883;
    wire N__23880;
    wire N__23877;
    wire N__23874;
    wire N__23871;
    wire N__23870;
    wire N__23867;
    wire N__23864;
    wire N__23859;
    wire N__23856;
    wire N__23853;
    wire N__23850;
    wire N__23847;
    wire N__23844;
    wire N__23841;
    wire N__23838;
    wire N__23835;
    wire N__23832;
    wire N__23831;
    wire N__23828;
    wire N__23827;
    wire N__23824;
    wire N__23821;
    wire N__23818;
    wire N__23811;
    wire N__23808;
    wire N__23805;
    wire N__23802;
    wire N__23799;
    wire N__23796;
    wire N__23793;
    wire N__23790;
    wire N__23787;
    wire N__23784;
    wire N__23781;
    wire N__23778;
    wire N__23775;
    wire N__23772;
    wire N__23769;
    wire N__23766;
    wire N__23763;
    wire N__23760;
    wire N__23757;
    wire N__23756;
    wire N__23753;
    wire N__23750;
    wire N__23747;
    wire N__23744;
    wire N__23741;
    wire N__23738;
    wire N__23733;
    wire N__23730;
    wire N__23727;
    wire N__23726;
    wire N__23723;
    wire N__23720;
    wire N__23715;
    wire N__23712;
    wire N__23709;
    wire N__23708;
    wire N__23705;
    wire N__23702;
    wire N__23697;
    wire N__23694;
    wire N__23691;
    wire N__23688;
    wire N__23685;
    wire N__23682;
    wire N__23679;
    wire N__23676;
    wire N__23673;
    wire N__23670;
    wire N__23667;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23655;
    wire N__23652;
    wire N__23649;
    wire N__23646;
    wire N__23643;
    wire N__23640;
    wire N__23637;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23620;
    wire N__23617;
    wire N__23614;
    wire N__23611;
    wire N__23604;
    wire N__23601;
    wire N__23598;
    wire N__23595;
    wire N__23592;
    wire N__23589;
    wire N__23586;
    wire N__23583;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23562;
    wire N__23559;
    wire N__23556;
    wire N__23553;
    wire N__23552;
    wire N__23551;
    wire N__23548;
    wire N__23543;
    wire N__23538;
    wire N__23535;
    wire N__23532;
    wire N__23529;
    wire N__23526;
    wire N__23523;
    wire N__23520;
    wire N__23517;
    wire N__23514;
    wire N__23511;
    wire N__23508;
    wire N__23505;
    wire N__23502;
    wire N__23499;
    wire N__23496;
    wire N__23493;
    wire N__23490;
    wire N__23487;
    wire N__23484;
    wire N__23481;
    wire N__23478;
    wire N__23475;
    wire N__23472;
    wire N__23469;
    wire N__23466;
    wire N__23463;
    wire N__23462;
    wire N__23459;
    wire N__23456;
    wire N__23453;
    wire N__23450;
    wire N__23447;
    wire N__23442;
    wire N__23439;
    wire N__23436;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23424;
    wire N__23421;
    wire N__23418;
    wire N__23415;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23400;
    wire N__23397;
    wire N__23394;
    wire N__23391;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23376;
    wire N__23373;
    wire N__23370;
    wire N__23367;
    wire N__23364;
    wire N__23361;
    wire N__23358;
    wire N__23355;
    wire N__23352;
    wire N__23349;
    wire N__23346;
    wire N__23343;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23331;
    wire N__23328;
    wire N__23325;
    wire N__23322;
    wire N__23319;
    wire N__23316;
    wire N__23313;
    wire N__23310;
    wire N__23307;
    wire N__23304;
    wire N__23303;
    wire N__23300;
    wire N__23297;
    wire N__23292;
    wire N__23289;
    wire N__23286;
    wire N__23283;
    wire N__23280;
    wire N__23277;
    wire N__23274;
    wire N__23271;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23259;
    wire N__23256;
    wire N__23253;
    wire N__23250;
    wire N__23247;
    wire N__23244;
    wire N__23241;
    wire N__23238;
    wire N__23235;
    wire N__23234;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23217;
    wire N__23214;
    wire N__23211;
    wire N__23208;
    wire N__23205;
    wire N__23202;
    wire N__23199;
    wire N__23196;
    wire N__23193;
    wire N__23190;
    wire N__23187;
    wire N__23184;
    wire N__23181;
    wire N__23178;
    wire N__23175;
    wire N__23172;
    wire N__23169;
    wire N__23166;
    wire N__23163;
    wire N__23160;
    wire N__23157;
    wire N__23154;
    wire N__23151;
    wire N__23148;
    wire N__23145;
    wire N__23142;
    wire N__23139;
    wire N__23136;
    wire N__23133;
    wire N__23130;
    wire N__23127;
    wire N__23124;
    wire N__23121;
    wire N__23118;
    wire N__23115;
    wire N__23112;
    wire N__23109;
    wire N__23106;
    wire N__23103;
    wire N__23100;
    wire N__23097;
    wire N__23096;
    wire N__23093;
    wire N__23090;
    wire N__23085;
    wire N__23082;
    wire N__23079;
    wire N__23076;
    wire N__23073;
    wire N__23070;
    wire N__23067;
    wire N__23064;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23052;
    wire N__23049;
    wire N__23046;
    wire N__23043;
    wire N__23040;
    wire N__23037;
    wire N__23034;
    wire N__23031;
    wire N__23028;
    wire N__23025;
    wire N__23022;
    wire N__23019;
    wire N__23016;
    wire N__23013;
    wire N__23010;
    wire N__23007;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22995;
    wire N__22992;
    wire N__22989;
    wire N__22986;
    wire N__22983;
    wire N__22980;
    wire N__22977;
    wire N__22974;
    wire N__22971;
    wire N__22968;
    wire N__22965;
    wire N__22962;
    wire N__22959;
    wire N__22956;
    wire N__22953;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22941;
    wire N__22938;
    wire N__22935;
    wire N__22932;
    wire N__22929;
    wire N__22926;
    wire N__22923;
    wire N__22920;
    wire N__22917;
    wire N__22914;
    wire N__22911;
    wire N__22908;
    wire N__22905;
    wire N__22902;
    wire N__22899;
    wire N__22896;
    wire N__22893;
    wire N__22890;
    wire N__22887;
    wire N__22884;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22860;
    wire N__22857;
    wire N__22854;
    wire N__22851;
    wire N__22848;
    wire N__22845;
    wire N__22844;
    wire N__22843;
    wire N__22840;
    wire N__22837;
    wire N__22834;
    wire N__22831;
    wire N__22828;
    wire N__22825;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22800;
    wire N__22799;
    wire N__22796;
    wire N__22793;
    wire N__22790;
    wire N__22785;
    wire N__22782;
    wire N__22779;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22767;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22757;
    wire N__22756;
    wire N__22753;
    wire N__22750;
    wire N__22747;
    wire N__22744;
    wire N__22741;
    wire N__22738;
    wire N__22731;
    wire N__22728;
    wire N__22725;
    wire N__22722;
    wire N__22719;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22694;
    wire N__22691;
    wire N__22690;
    wire N__22687;
    wire N__22684;
    wire N__22681;
    wire N__22678;
    wire N__22675;
    wire N__22672;
    wire N__22665;
    wire N__22662;
    wire N__22659;
    wire N__22656;
    wire N__22653;
    wire N__22650;
    wire N__22647;
    wire N__22644;
    wire N__22641;
    wire N__22638;
    wire N__22635;
    wire N__22632;
    wire N__22629;
    wire N__22626;
    wire N__22623;
    wire N__22620;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22608;
    wire N__22605;
    wire N__22602;
    wire N__22599;
    wire N__22596;
    wire N__22593;
    wire N__22590;
    wire N__22587;
    wire N__22584;
    wire N__22583;
    wire N__22582;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22566;
    wire N__22563;
    wire N__22560;
    wire N__22557;
    wire N__22554;
    wire N__22551;
    wire N__22548;
    wire N__22545;
    wire N__22542;
    wire N__22539;
    wire N__22536;
    wire N__22533;
    wire N__22530;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22518;
    wire N__22515;
    wire N__22512;
    wire N__22509;
    wire N__22506;
    wire N__22503;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22491;
    wire N__22488;
    wire N__22485;
    wire N__22482;
    wire N__22479;
    wire N__22476;
    wire N__22473;
    wire N__22470;
    wire N__22467;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22455;
    wire N__22452;
    wire N__22449;
    wire N__22446;
    wire N__22443;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22428;
    wire N__22425;
    wire N__22422;
    wire N__22419;
    wire N__22416;
    wire N__22413;
    wire N__22410;
    wire N__22407;
    wire N__22404;
    wire N__22401;
    wire N__22398;
    wire N__22395;
    wire N__22392;
    wire N__22389;
    wire N__22386;
    wire N__22383;
    wire N__22380;
    wire N__22377;
    wire N__22374;
    wire N__22371;
    wire N__22368;
    wire N__22365;
    wire N__22362;
    wire N__22359;
    wire N__22356;
    wire N__22353;
    wire N__22350;
    wire N__22347;
    wire N__22344;
    wire N__22341;
    wire N__22338;
    wire N__22335;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22320;
    wire N__22317;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22284;
    wire N__22281;
    wire N__22278;
    wire N__22275;
    wire N__22272;
    wire N__22269;
    wire N__22266;
    wire N__22263;
    wire N__22260;
    wire N__22257;
    wire N__22254;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22242;
    wire N__22239;
    wire N__22236;
    wire N__22233;
    wire N__22230;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22212;
    wire N__22209;
    wire N__22206;
    wire N__22203;
    wire N__22200;
    wire N__22197;
    wire N__22194;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22182;
    wire N__22179;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22167;
    wire N__22164;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22152;
    wire N__22149;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22125;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22110;
    wire N__22107;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22097;
    wire N__22094;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22071;
    wire N__22070;
    wire N__22065;
    wire N__22062;
    wire N__22059;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22047;
    wire N__22044;
    wire N__22043;
    wire N__22040;
    wire N__22037;
    wire N__22032;
    wire N__22029;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22019;
    wire N__22014;
    wire N__22011;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__21999;
    wire N__21996;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21972;
    wire N__21969;
    wire N__21968;
    wire N__21963;
    wire N__21960;
    wire N__21959;
    wire N__21956;
    wire N__21951;
    wire N__21948;
    wire N__21945;
    wire N__21942;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21924;
    wire N__21921;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21903;
    wire N__21900;
    wire N__21897;
    wire N__21894;
    wire N__21891;
    wire N__21888;
    wire N__21885;
    wire N__21882;
    wire N__21879;
    wire N__21876;
    wire N__21873;
    wire N__21870;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21858;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21819;
    wire N__21816;
    wire N__21813;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21801;
    wire N__21798;
    wire N__21795;
    wire N__21792;
    wire N__21789;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21759;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21732;
    wire N__21729;
    wire N__21726;
    wire N__21723;
    wire N__21720;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21708;
    wire N__21705;
    wire N__21702;
    wire N__21699;
    wire N__21696;
    wire N__21693;
    wire N__21690;
    wire N__21687;
    wire N__21684;
    wire N__21681;
    wire N__21678;
    wire N__21675;
    wire N__21672;
    wire N__21669;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire GNDG0;
    wire bfn_1_19_0_;
    wire n12696;
    wire n12697;
    wire n12698;
    wire n12699;
    wire n12700;
    wire n12701;
    wire n12702;
    wire n12703;
    wire bfn_1_20_0_;
    wire n12704;
    wire n12705;
    wire n12706;
    wire n12707;
    wire n12708;
    wire n12709;
    wire n12710;
    wire n12711;
    wire bfn_1_21_0_;
    wire n12712;
    wire n12713;
    wire n12714;
    wire n12715;
    wire n12716;
    wire bfn_1_22_0_;
    wire n12811;
    wire n12812;
    wire n12813;
    wire n12814;
    wire n12815;
    wire n12816;
    wire n12817;
    wire n12818;
    wire bfn_1_23_0_;
    wire n12819;
    wire n12820;
    wire n12821;
    wire n12822;
    wire n12823;
    wire n12824;
    wire n12825;
    wire n12826;
    wire bfn_1_24_0_;
    wire n12827;
    wire n12828;
    wire n12829;
    wire n12830;
    wire n12831;
    wire n12832;
    wire n12833;
    wire n12834;
    wire bfn_1_25_0_;
    wire n12835;
    wire n12836;
    wire n2882;
    wire n2900;
    wire n2876;
    wire n2908_cascade_;
    wire n2895;
    wire n2927_cascade_;
    wire n3024_cascade_;
    wire n14730_cascade_;
    wire n3021_cascade_;
    wire n14728;
    wire n14150_cascade_;
    wire n3128_cascade_;
    wire n14148;
    wire n3120_cascade_;
    wire n3122_cascade_;
    wire n14146;
    wire \debounce.reg_A_2 ;
    wire \debounce.reg_A_1 ;
    wire \debounce.reg_A_0 ;
    wire reg_B_0;
    wire \debounce.n6_cascade_ ;
    wire \debounce.n16_cascade_ ;
    wire \debounce.n17 ;
    wire reg_B_2;
    wire n14129_cascade_;
    wire \debounce.cnt_reg_0 ;
    wire bfn_1_31_0_;
    wire \debounce.cnt_reg_1 ;
    wire \debounce.n13013 ;
    wire \debounce.cnt_reg_2 ;
    wire \debounce.n13014 ;
    wire \debounce.cnt_reg_3 ;
    wire \debounce.n13015 ;
    wire \debounce.cnt_reg_4 ;
    wire \debounce.n13016 ;
    wire \debounce.cnt_reg_5 ;
    wire \debounce.n13017 ;
    wire \debounce.cnt_reg_6 ;
    wire \debounce.n13018 ;
    wire \debounce.cnt_reg_7 ;
    wire \debounce.n13019 ;
    wire \debounce.n13020 ;
    wire \debounce.cnt_reg_8 ;
    wire bfn_1_32_0_;
    wire \debounce.n13021 ;
    wire \debounce.cnt_reg_9 ;
    wire \debounce.cnt_next_9__N_424 ;
    wire bfn_2_13_0_;
    wire n12762;
    wire n12763;
    wire n12764;
    wire n12765;
    wire n12766;
    wire n12767;
    wire n12768;
    wire n12769;
    wire bfn_2_14_0_;
    wire n12770;
    wire n12771;
    wire n12772;
    wire n12773;
    wire n12774;
    wire n12775;
    wire n12776;
    wire n12777;
    wire bfn_2_15_0_;
    wire n12778;
    wire n12779;
    wire n2682;
    wire n12780;
    wire n12781;
    wire n12782;
    wire n12783;
    wire n12784;
    wire n12785;
    wire bfn_2_16_0_;
    wire n2801;
    wire bfn_2_17_0_;
    wire n12786;
    wire n12787;
    wire n12788;
    wire n12789;
    wire n12790;
    wire n12791;
    wire n12792;
    wire n12793;
    wire bfn_2_18_0_;
    wire n12794;
    wire n12795;
    wire n12796;
    wire n12797;
    wire n12798;
    wire n12799;
    wire n12800;
    wire n12801;
    wire bfn_2_19_0_;
    wire n12802;
    wire n2783;
    wire n12803;
    wire n12804;
    wire n12805;
    wire n12806;
    wire n12807;
    wire n12808;
    wire n12809;
    wire bfn_2_20_0_;
    wire n12810;
    wire n2683;
    wire n2677;
    wire n2678;
    wire n2797;
    wire n2694;
    wire n2793;
    wire n2726_cascade_;
    wire n2621_cascade_;
    wire n2688;
    wire n2696;
    wire n2795;
    wire n2728_cascade_;
    wire n2691;
    wire n2723;
    wire n2790;
    wire n2723_cascade_;
    wire n2693;
    wire n2697;
    wire n2681;
    wire n2794;
    wire n2826_cascade_;
    wire n14362_cascade_;
    wire n2789;
    wire n14346;
    wire n14350_cascade_;
    wire n14356;
    wire n2782;
    wire n2715;
    wire n2785;
    wire n2684;
    wire n2716;
    wire n2679;
    wire n2709;
    wire n2711_cascade_;
    wire n14368;
    wire n2796;
    wire n2742_cascade_;
    wire n2828;
    wire n2788;
    wire n2687;
    wire n2792;
    wire n2725;
    wire n2791;
    wire bfn_2_25_0_;
    wire n12837;
    wire n12838;
    wire n12839;
    wire n12840;
    wire n12841;
    wire n12842;
    wire n2994;
    wire n12843;
    wire n12844;
    wire n2993;
    wire bfn_2_26_0_;
    wire n2992;
    wire n12845;
    wire n12846;
    wire n2990;
    wire n12847;
    wire n2989;
    wire n12848;
    wire n12849;
    wire n12850;
    wire n12851;
    wire n12852;
    wire n2985;
    wire bfn_2_27_0_;
    wire n12853;
    wire n12854;
    wire n12855;
    wire n12856;
    wire n12857;
    wire n12858;
    wire n12859;
    wire n12860;
    wire n2977;
    wire bfn_2_28_0_;
    wire n12861;
    wire n2975;
    wire n12862;
    wire n12863;
    wire bfn_2_29_0_;
    wire n12892;
    wire n12893;
    wire n12894;
    wire n12895;
    wire n12896;
    wire n12897;
    wire n12898;
    wire n12899;
    wire bfn_2_30_0_;
    wire n12900;
    wire n12901;
    wire n12902;
    wire n12903;
    wire n12904;
    wire n3120;
    wire n3187;
    wire n12905;
    wire n12906;
    wire n12907;
    wire bfn_2_31_0_;
    wire n12908;
    wire n12909;
    wire n12910;
    wire n12911;
    wire n12912;
    wire n12913;
    wire n12914;
    wire n12915;
    wire bfn_2_32_0_;
    wire n12916;
    wire n12917;
    wire n12918;
    wire n12919;
    wire n12920;
    wire bfn_3_14_0_;
    wire n12676;
    wire n12677;
    wire n12678;
    wire n12679;
    wire n12680;
    wire n12681;
    wire n12682;
    wire n12683;
    wire bfn_3_15_0_;
    wire n12684;
    wire n12685;
    wire n12686;
    wire n12687;
    wire n12688;
    wire n12689;
    wire n12690;
    wire n12691;
    wire bfn_3_16_0_;
    wire n12692;
    wire n12693;
    wire n12694;
    wire n12695;
    wire n2233;
    wire n2300;
    wire n2233_cascade_;
    wire n2299;
    wire n2331_cascade_;
    wire n2301;
    wire n2222;
    wire n2222_cascade_;
    wire n2289;
    wire n2291;
    wire n2323_cascade_;
    wire n2219_cascade_;
    wire n2286;
    wire n2290;
    wire n2293;
    wire n2298;
    wire n2295;
    wire n2296;
    wire n11977;
    wire n14808_cascade_;
    wire n14594;
    wire n2219;
    wire n14598_cascade_;
    wire n14604_cascade_;
    wire n2247_cascade_;
    wire n2297;
    wire n2288;
    wire n2391;
    wire n2287;
    wire n2386;
    wire n2319_cascade_;
    wire n11971;
    wire n2292;
    wire n2324;
    wire n2324_cascade_;
    wire n2319;
    wire n14384_cascade_;
    wire n14382;
    wire n14390;
    wire n2689;
    wire n2622_cascade_;
    wire n2721;
    wire n2728;
    wire n2726;
    wire n2721_cascade_;
    wire n14348;
    wire n2383;
    wire n2622;
    wire n2628_cascade_;
    wire n2692;
    wire n2724;
    wire n2695;
    wire n2628;
    wire n2727;
    wire n2700;
    wire n2732_cascade_;
    wire n2729;
    wire n11957_cascade_;
    wire n13808;
    wire n2621;
    wire n14668;
    wire n2698;
    wire n2730;
    wire n2699;
    wire n2701;
    wire n14650_cascade_;
    wire n14654_cascade_;
    wire n14660_cascade_;
    wire n14674;
    wire n2643_cascade_;
    wire n2686;
    wire n2718;
    wire n2690;
    wire n2623;
    wire n2722;
    wire n2732;
    wire n2799;
    wire n2711;
    wire n2778;
    wire n2786;
    wire n2719;
    wire n2685;
    wire n2717;
    wire n2784;
    wire n2717_cascade_;
    wire n2713;
    wire n2780;
    wire n2798;
    wire n2731;
    wire n2680;
    wire n2887;
    wire n2820;
    wire n14690_cascade_;
    wire n14688;
    wire n14696_cascade_;
    wire n2714;
    wire n2781;
    wire n2720;
    wire n2787;
    wire n2823;
    wire n2890;
    wire n2827;
    wire n2894;
    wire n2822;
    wire n2889;
    wire n2982;
    wire n2986;
    wire n2879;
    wire n2710;
    wire n2777;
    wire n2996;
    wire n3028_cascade_;
    wire n2988;
    wire n2880;
    wire n2979;
    wire n2912_cascade_;
    wire n2983;
    wire bfn_3_28_0_;
    wire n12864;
    wire n12865;
    wire n12866;
    wire n12867;
    wire n3096;
    wire n12868;
    wire n3028;
    wire n3095;
    wire n12869;
    wire n3094;
    wire n12870;
    wire n12871;
    wire n3026;
    wire n3093;
    wire bfn_3_29_0_;
    wire n3025;
    wire n3092;
    wire n12872;
    wire n3024;
    wire n3091;
    wire n12873;
    wire n3090;
    wire n12874;
    wire n3022;
    wire n3089;
    wire n12875;
    wire n3021;
    wire n3088;
    wire n12876;
    wire n3020;
    wire n3087;
    wire n12877;
    wire n3086;
    wire n12878;
    wire n12879;
    wire bfn_3_30_0_;
    wire n3017;
    wire n3084;
    wire n12880;
    wire n12881;
    wire n12882;
    wire n12883;
    wire n12884;
    wire n12885;
    wire n12886;
    wire n12887;
    wire bfn_3_31_0_;
    wire n12888;
    wire n12889;
    wire n12890;
    wire n12891;
    wire n3075;
    wire n3082;
    wire n3074;
    wire n3173;
    wire n3174;
    wire n3079;
    wire n3078;
    wire n3076;
    wire n3175;
    wire n3108_cascade_;
    wire n2232;
    wire n2231;
    wire n2221;
    wire n2229;
    wire n2129_cascade_;
    wire n2228;
    wire n2226;
    wire n2225;
    wire n2228_cascade_;
    wire n14588;
    wire n2201;
    wire bfn_4_17_0_;
    wire n2200;
    wire n12657;
    wire n2199;
    wire n12658;
    wire n12659;
    wire n2197;
    wire n12660;
    wire n2129;
    wire n2196;
    wire n12661;
    wire n12662;
    wire n2194;
    wire n12663;
    wire n12664;
    wire n2193;
    wire bfn_4_18_0_;
    wire n12665;
    wire n12666;
    wire n2190;
    wire n12667;
    wire n2189;
    wire n12668;
    wire n12669;
    wire n2187;
    wire n12670;
    wire n12671;
    wire n12672;
    wire bfn_4_19_0_;
    wire n12673;
    wire n12674;
    wire n12675;
    wire n2214;
    wire n2294;
    wire n2186;
    wire n2218;
    wire n2285;
    wire n2218_cascade_;
    wire n2188;
    wire n2220;
    wire n14392;
    wire n2313;
    wire n14398_cascade_;
    wire n2327;
    wire n2346_cascade_;
    wire n2394;
    wire n2284;
    wire n2316;
    wire n2282;
    wire n2314;
    wire n2314_cascade_;
    wire n2381;
    wire n2392;
    wire n2325;
    wire n2320;
    wire n2387;
    wire n2382;
    wire n2396;
    wire n2329;
    wire n2328;
    wire n2395;
    wire n2427_cascade_;
    wire n14620_cascade_;
    wire n2526_cascade_;
    wire n14816;
    wire n2524_cascade_;
    wire n14574_cascade_;
    wire n2523_cascade_;
    wire n14576;
    wire n2527_cascade_;
    wire n2626;
    wire n2617;
    wire n2625;
    wire n2617_cascade_;
    wire n14812;
    wire n2633;
    wire n2633_cascade_;
    wire n12059;
    wire n2618;
    wire n2614;
    wire n2613;
    wire n2619;
    wire n2897;
    wire n2712;
    wire n2779;
    wire n2878;
    wire n2811_cascade_;
    wire n2733;
    wire n2800;
    wire n2832_cascade_;
    wire n2833;
    wire n2830;
    wire n11953_cascade_;
    wire n13857;
    wire n2815;
    wire n14702;
    wire n2812;
    wire n2813;
    wire n14708_cascade_;
    wire n2811;
    wire n2809;
    wire n14714_cascade_;
    wire n2808;
    wire n2816;
    wire n2841_cascade_;
    wire n2883;
    wire n2885;
    wire n2818;
    wire n3081;
    wire n2810;
    wire n2877;
    wire n2976;
    wire n2886;
    wire n2819;
    wire n2918;
    wire n2927;
    wire n2926;
    wire n2918_cascade_;
    wire n2825;
    wire n2892;
    wire n2921;
    wire n2922;
    wire n2924_cascade_;
    wire n2919;
    wire n14212_cascade_;
    wire n14216;
    wire n2817;
    wire n2884;
    wire n2916;
    wire n2981;
    wire n2929;
    wire n14222;
    wire n2915;
    wire n14224_cascade_;
    wire n2914;
    wire n2910;
    wire n14230_cascade_;
    wire n2912;
    wire n2908;
    wire n2907;
    wire n14236_cascade_;
    wire n2909;
    wire n2940_cascade_;
    wire n2997;
    wire n2911;
    wire n2978;
    wire n2995;
    wire n3000;
    wire n3015;
    wire n14736;
    wire n3014;
    wire n14742_cascade_;
    wire n3011;
    wire n3009;
    wire n14748_cascade_;
    wire n3006;
    wire n3008;
    wire n14754_cascade_;
    wire n3007;
    wire n3099;
    wire n3039_cascade_;
    wire n3018;
    wire n3085;
    wire n3098;
    wire n3130_cascade_;
    wire n3101;
    wire n3097;
    wire n3100;
    wire n3132_cascade_;
    wire n11945;
    wire n3080;
    wire n3013;
    wire n23_adj_715_cascade_;
    wire n3123;
    wire n3190;
    wire n3121;
    wire n3188;
    wire n3192;
    wire n3125;
    wire n3127;
    wire n3194;
    wire n3226_cascade_;
    wire n3119;
    wire n3186;
    wire n3218_cascade_;
    wire n3180;
    wire n3212_cascade_;
    wire n14798;
    wire n3107;
    wire n3106;
    wire n3105;
    wire n3195;
    wire n3138_cascade_;
    wire n3128;
    wire n3181;
    wire n3184;
    wire n3117;
    wire n3083;
    wire n13831;
    wire n3114;
    wire n3115_cascade_;
    wire n14156;
    wire n3113;
    wire n14162_cascade_;
    wire n14168_cascade_;
    wire n3108;
    wire n14174;
    wire n3010;
    wire n3077;
    wire n14264;
    wire n14260;
    wire n2130;
    wire n14324_cascade_;
    wire n13787;
    wire n2127;
    wire n2127_cascade_;
    wire n14318;
    wire n2131;
    wire n2198;
    wire n2131_cascade_;
    wire n2230;
    wire n14584;
    wire n2191;
    wire n2223;
    wire n2192;
    wire n2224;
    wire n14330;
    wire n2116_cascade_;
    wire n2148_cascade_;
    wire n2195;
    wire n2227;
    wire n2128;
    wire n2126;
    wire n2128_cascade_;
    wire n14316;
    wire n2125;
    wire n2185;
    wire n2217;
    wire n2183;
    wire n2116;
    wire n2215;
    wire n2184;
    wire n2122;
    wire n2124;
    wire n2401;
    wire n2390;
    wire n2323;
    wire n2118;
    wire n2393;
    wire n2326;
    wire n2330;
    wire n2397;
    wire n2322;
    wire n2389;
    wire n2399;
    wire n2332;
    wire n2388;
    wire n2321;
    wire n2420_cascade_;
    wire n14622;
    wire n2398;
    wire n2331;
    wire n2430_cascade_;
    wire n2400;
    wire n2333;
    wire n2432_cascade_;
    wire n11967;
    wire n2528_cascade_;
    wire n2627;
    wire n2384;
    wire n2317;
    wire n13828;
    wire n14628;
    wire n2318;
    wire n2385;
    wire n2417_cascade_;
    wire n14634;
    wire n14640_cascade_;
    wire n2445_cascade_;
    wire n2530_cascade_;
    wire n14646;
    wire n2533_cascade_;
    wire n12063;
    wire n2632;
    wire n14188;
    wire n2515_cascade_;
    wire n14117;
    wire n14194_cascade_;
    wire n2544_cascade_;
    wire n2631;
    wire n2513_cascade_;
    wire n2612;
    wire n2629;
    wire n2899;
    wire n2832;
    wire n2630;
    wire n2620;
    wire n2901;
    wire n2824;
    wire n2891;
    wire n2923;
    wire n2923_cascade_;
    wire n14214;
    wire n2896;
    wire n2829;
    wire n2928;
    wire n2821;
    wire n2888;
    wire n2881;
    wire n2814;
    wire n2893;
    wire n2826;
    wire n2925;
    wire n2615;
    wire n2831;
    wire n2898;
    wire n2930;
    wire n2991;
    wire n2924;
    wire n2913;
    wire n2980;
    wire n3012;
    wire n2933;
    wire n12053;
    wire n2987;
    wire n2920;
    wire n2999;
    wire n2932;
    wire n3001;
    wire n3033;
    wire n3033_cascade_;
    wire n3032;
    wire n3182;
    wire n3115;
    wire n2998;
    wire n2931;
    wire n3030;
    wire n3029;
    wire n3031;
    wire n3030_cascade_;
    wire n11947;
    wire n3019;
    wire n3027;
    wire n13871_cascade_;
    wire n3023;
    wire n14078;
    wire n3199;
    wire n3132;
    wire n3129;
    wire n3196;
    wire n3228_cascade_;
    wire n14768;
    wire n3200;
    wire n3133;
    wire n3198;
    wire n3131;
    wire n2917;
    wire n2984;
    wire n3016;
    wire n3124;
    wire n3191;
    wire n14804;
    wire n14025;
    wire n3237_cascade_;
    wire n13_adj_713;
    wire n3179;
    wire n3112;
    wire n14770;
    wire n14776_cascade_;
    wire n3122;
    wire n3189;
    wire n3116;
    wire n3183;
    wire n3185;
    wire n3118;
    wire n27_adj_716_cascade_;
    wire n14266;
    wire n35_adj_719;
    wire n17_adj_714_cascade_;
    wire n3109;
    wire n3176;
    wire n33_adj_718_cascade_;
    wire n14272;
    wire n14268;
    wire n14262_cascade_;
    wire n14282;
    wire n3111;
    wire n3178;
    wire n3110;
    wire n3177;
    wire n2283;
    wire n2216;
    wire n2315;
    wire bfn_6_17_0_;
    wire n12639;
    wire n2099;
    wire n12640;
    wire n2098;
    wire n12641;
    wire n2097;
    wire n12642;
    wire n2096;
    wire n12643;
    wire n2095;
    wire n12644;
    wire n2094;
    wire n12645;
    wire n12646;
    wire n2093;
    wire bfn_6_18_0_;
    wire n2092;
    wire n12647;
    wire n12648;
    wire n2090;
    wire n12649;
    wire n12650;
    wire n12651;
    wire n12652;
    wire n2086;
    wire n12653;
    wire n12654;
    wire bfn_6_19_0_;
    wire n2084;
    wire n12655;
    wire n12656;
    wire n2115;
    wire n2091;
    wire n2123;
    wire n14558_cascade_;
    wire n2101;
    wire n2049_cascade_;
    wire n2018;
    wire n2085;
    wire n2018_cascade_;
    wire n2117;
    wire n2089;
    wire n2121;
    wire n2501;
    wire bfn_6_21_0_;
    wire n12717;
    wire n2432;
    wire n2499;
    wire n12718;
    wire n2431;
    wire n2498;
    wire n12719;
    wire n2430;
    wire n2497;
    wire n12720;
    wire n2429;
    wire n2496;
    wire n12721;
    wire n2428;
    wire n2495;
    wire n12722;
    wire n2427;
    wire n2494;
    wire n12723;
    wire n12724;
    wire bfn_6_22_0_;
    wire n2425;
    wire n2492;
    wire n12725;
    wire n2424;
    wire n2491;
    wire n12726;
    wire n12727;
    wire n12728;
    wire n2421;
    wire n2488;
    wire n12729;
    wire n2420;
    wire n2487;
    wire n12730;
    wire n12731;
    wire n12732;
    wire bfn_6_23_0_;
    wire n2417;
    wire n2484;
    wire n12733;
    wire n2416;
    wire n2483;
    wire n12734;
    wire n2415;
    wire n2482;
    wire n12735;
    wire n2414;
    wire n2481;
    wire n12736;
    wire n2413;
    wire n2480;
    wire n12737;
    wire n2412;
    wire n12738;
    wire n2433;
    wire n2500;
    wire n2601;
    wire bfn_6_24_0_;
    wire n2533;
    wire n2600;
    wire n12739;
    wire n2532;
    wire n2599;
    wire n12740;
    wire n2531;
    wire n2598;
    wire n12741;
    wire n2530;
    wire n2597;
    wire n12742;
    wire n2529;
    wire n2596;
    wire n12743;
    wire n2528;
    wire n2595;
    wire n12744;
    wire n2527;
    wire n2594;
    wire n12745;
    wire n12746;
    wire n2526;
    wire n2593;
    wire bfn_6_25_0_;
    wire n12747;
    wire n2524;
    wire n2591;
    wire n12748;
    wire n2523;
    wire n2590;
    wire n12749;
    wire n2589;
    wire n12750;
    wire n2588;
    wire n12751;
    wire n2520;
    wire n2587;
    wire n12752;
    wire n2519;
    wire n2586;
    wire n12753;
    wire n12754;
    wire n2585;
    wire bfn_6_26_0_;
    wire n12755;
    wire n2516;
    wire n2583;
    wire n12756;
    wire n2515;
    wire n2582;
    wire n12757;
    wire n2514;
    wire n2581;
    wire n12758;
    wire n2513;
    wire n2580;
    wire n12759;
    wire n12760;
    wire n2511;
    wire n12761;
    wire n2610;
    wire n2418;
    wire n2485;
    wire n2517;
    wire n2584;
    wire n2517_cascade_;
    wire n2616;
    wire n2512;
    wire n2579;
    wire n2611;
    wire n3130;
    wire n3197;
    wire n3193;
    wire n3126;
    wire n3201;
    wire n3233_cascade_;
    wire n11943_cascade_;
    wire n13875;
    wire n29_adj_717_cascade_;
    wire n14270;
    wire n11941_cascade_;
    wire n11878;
    wire n14782;
    wire n14788;
    wire n14300_cascade_;
    wire n14302_cascade_;
    wire n14304_cascade_;
    wire n14306_cascade_;
    wire n14308;
    wire n5_adj_704;
    wire n12039;
    wire n14292_cascade_;
    wire n14284;
    wire n14286_cascade_;
    wire n14288;
    wire n14294;
    wire n14296_cascade_;
    wire n14298;
    wire n45_adj_720;
    wire ENCODER0_A_N;
    wire n1922_cascade_;
    wire n2021;
    wire n2088;
    wire n2021_cascade_;
    wire n2120;
    wire n2020;
    wire n2087;
    wire n2020_cascade_;
    wire n2119;
    wire n14446_cascade_;
    wire n11985;
    wire n14450_cascade_;
    wire n1950_cascade_;
    wire n2017;
    wire n2025;
    wire n2028;
    wire n2026;
    wire n2025_cascade_;
    wire n2027;
    wire n2032;
    wire n2031;
    wire n2032_cascade_;
    wire n2022;
    wire n2024;
    wire n2023;
    wire n14544;
    wire n11981;
    wire n2029;
    wire n14550_cascade_;
    wire n2030;
    wire n14552;
    wire n2100;
    wire n2033;
    wire n2132;
    wire n2132_cascade_;
    wire n2133;
    wire n11909;
    wire n307;
    wire n310;
    wire n312;
    wire n313;
    wire n314;
    wire n317;
    wire n14184;
    wire n2490;
    wire n2423;
    wire n2522;
    wire n2489;
    wire n2422;
    wire n2521;
    wire n2426;
    wire n2493;
    wire n2525;
    wire n2592;
    wire n2525_cascade_;
    wire n2624;
    wire n2486;
    wire n2419;
    wire n2518;
    wire n315;
    wire n311;
    wire bfn_7_25_0_;
    wire n15485;
    wire n3237;
    wire n12952;
    wire n15451;
    wire n3138;
    wire n12953;
    wire n15418;
    wire n3039;
    wire n12954;
    wire n15384;
    wire n2940;
    wire n12955;
    wire n15352;
    wire n2841;
    wire n12956;
    wire n15322;
    wire n2742;
    wire n12957;
    wire n15292;
    wire n2643;
    wire encoder0_position_scaled_7;
    wire n12958;
    wire n12959;
    wire n15830;
    wire n2544;
    wire bfn_7_26_0_;
    wire n15802;
    wire n2445;
    wire n12960;
    wire n15775;
    wire n2346;
    wire n12961;
    wire n15748;
    wire n2247;
    wire n12962;
    wire n15722;
    wire n2148;
    wire n12963;
    wire n15697;
    wire n2049;
    wire n12964;
    wire n12965;
    wire n15652;
    wire n12966;
    wire n12967;
    wire bfn_7_27_0_;
    wire n12968;
    wire n12969;
    wire n12970;
    wire n12971;
    wire n12972;
    wire n12973;
    wire n12974;
    wire n12051;
    wire n15490;
    wire n319;
    wire bfn_7_29_0_;
    wire n318;
    wire n3301;
    wire n12921;
    wire n3233;
    wire n3300;
    wire n12922;
    wire n3232;
    wire n3299;
    wire n12923;
    wire n3231;
    wire n12924;
    wire n3298;
    wire n3230;
    wire n15079;
    wire n12925;
    wire n3229;
    wire n3296;
    wire n12926;
    wire n3228;
    wire n3295;
    wire n12927;
    wire n12928;
    wire n3227;
    wire n3294;
    wire bfn_7_30_0_;
    wire n3226;
    wire n3293;
    wire n12929;
    wire n3225;
    wire n3292;
    wire n12930;
    wire n3224;
    wire n3291;
    wire n12931;
    wire n3223;
    wire n3290;
    wire n12932;
    wire n3222;
    wire n3289;
    wire n12933;
    wire n3221;
    wire n3288;
    wire n12934;
    wire n3220;
    wire n3287;
    wire n12935;
    wire n12936;
    wire n3219;
    wire n3286;
    wire bfn_7_31_0_;
    wire n3218;
    wire n3285;
    wire n12937;
    wire n3217;
    wire n3284;
    wire n12938;
    wire n3216;
    wire n3283;
    wire n12939;
    wire n3215;
    wire n3282;
    wire n12940;
    wire n3214;
    wire n3281;
    wire n12941;
    wire n3213;
    wire n3280;
    wire n12942;
    wire n3212;
    wire n3279;
    wire n12943;
    wire n12944;
    wire n3211;
    wire n3278;
    wire bfn_7_32_0_;
    wire n3210;
    wire n3277;
    wire n12945;
    wire n3209;
    wire n3276;
    wire n12946;
    wire n3208;
    wire n3275;
    wire n12947;
    wire n3207;
    wire n3274;
    wire n12948;
    wire n3206;
    wire n3273;
    wire n12949;
    wire n3205;
    wire n3272;
    wire n12950;
    wire n3204;
    wire n12951;
    wire n3271;
    wire n2001;
    wire bfn_9_16_0_;
    wire n2000;
    wire n12622;
    wire n1999;
    wire n12623;
    wire n1998;
    wire n12624;
    wire n1997;
    wire n12625;
    wire n1996;
    wire n12626;
    wire n1995;
    wire n12627;
    wire n1994;
    wire n12628;
    wire n12629;
    wire n1993;
    wire bfn_9_17_0_;
    wire n1992;
    wire n12630;
    wire n1991;
    wire n12631;
    wire n1990;
    wire n12632;
    wire n1922;
    wire n1989;
    wire n12633;
    wire n1988;
    wire n12634;
    wire n12635;
    wire n1986;
    wire n12636;
    wire n12637;
    wire n1985;
    wire bfn_9_18_0_;
    wire n15674;
    wire n12638;
    wire n2016;
    wire n1921;
    wire n14530;
    wire n1918;
    wire n1919;
    wire n305;
    wire n306;
    wire n308;
    wire n309;
    wire n33_adj_651;
    wire n33;
    wire bfn_9_22_0_;
    wire n32;
    wire n12975;
    wire n31_adj_649;
    wire n31;
    wire n12976;
    wire n30_adj_648;
    wire n12977;
    wire n29_adj_647;
    wire n29;
    wire n12978;
    wire n28_adj_646;
    wire n28;
    wire n12979;
    wire n27_adj_645;
    wire n27;
    wire n12980;
    wire n26_adj_644;
    wire n26;
    wire n12981;
    wire n12982;
    wire n25_adj_643;
    wire n25;
    wire bfn_9_23_0_;
    wire n24_adj_642;
    wire n24;
    wire n12983;
    wire n23_adj_641;
    wire n23;
    wire n12984;
    wire n22;
    wire n12985;
    wire n21;
    wire n12986;
    wire n20;
    wire n12987;
    wire n19_adj_637;
    wire n19;
    wire n12988;
    wire n18_adj_636;
    wire n18;
    wire n12989;
    wire n12990;
    wire bfn_9_24_0_;
    wire n12991;
    wire n12992;
    wire n14_adj_632;
    wire n14;
    wire n12993;
    wire n12994;
    wire n12995;
    wire n12996;
    wire n12997;
    wire n12998;
    wire bfn_9_25_0_;
    wire n12999;
    wire n13000;
    wire n13001;
    wire n13002;
    wire n4_adj_622;
    wire n13003;
    wire n13004;
    wire n13005;
    wire encoder0_position_scaled_8;
    wire encoder0_position_scaled_14;
    wire encoder0_position_scaled_10;
    wire encoder0_position_scaled_12;
    wire encoder0_position_scaled_13;
    wire encoder0_position_scaled_15;
    wire n15508;
    wire encoder0_position_scaled_18;
    wire encoder0_position_scaled_23;
    wire encoder0_position_scaled_17;
    wire dti_N_333_cascade_;
    wire reg_B_1;
    wire n14129;
    wire n1377;
    wire bfn_9_29_0_;
    wire n13006;
    wire n13007;
    wire n13008;
    wire n13009;
    wire n15072;
    wire n13010;
    wire n13011;
    wire n11526;
    wire n13012;
    wire n15075;
    wire n15071;
    wire dti_counter_5;
    wire dti_counter_6;
    wire n14_adj_705_cascade_;
    wire dti_counter_2;
    wire n10_adj_706;
    wire dti_counter_0;
    wire n15081;
    wire dti_counter_3;
    wire n15074;
    wire dti_counter_4;
    wire n15073;
    wire dti_counter_7;
    wire n15070;
    wire dti_counter_1;
    wire n15076;
    wire commutation_state_prev_0;
    wire n14929;
    wire n14928;
    wire LED_c;
    wire n1831_cascade_;
    wire n1930;
    wire n1931;
    wire n1933;
    wire n1929;
    wire n14524_cascade_;
    wire n14526_cascade_;
    wire n1851_cascade_;
    wire n1928;
    wire n1925;
    wire n1928_cascade_;
    wire n1923;
    wire n14440;
    wire n1932;
    wire encoder0_position_0;
    wire bfn_10_18_0_;
    wire \quad_counter0.n13095 ;
    wire encoder0_position_2;
    wire \quad_counter0.n13096 ;
    wire \quad_counter0.n13097 ;
    wire encoder0_position_4;
    wire \quad_counter0.n13098 ;
    wire encoder0_position_5;
    wire \quad_counter0.n13099 ;
    wire encoder0_position_6;
    wire \quad_counter0.n13100 ;
    wire encoder0_position_7;
    wire \quad_counter0.n13101 ;
    wire \quad_counter0.n13102 ;
    wire encoder0_position_8;
    wire bfn_10_19_0_;
    wire encoder0_position_9;
    wire \quad_counter0.n13103 ;
    wire encoder0_position_10;
    wire \quad_counter0.n13104 ;
    wire \quad_counter0.n13105 ;
    wire \quad_counter0.n13106 ;
    wire \quad_counter0.n13107 ;
    wire encoder0_position_14;
    wire \quad_counter0.n13108 ;
    wire encoder0_position_15;
    wire \quad_counter0.n13109 ;
    wire \quad_counter0.n13110 ;
    wire bfn_10_20_0_;
    wire \quad_counter0.n13111 ;
    wire \quad_counter0.n13112 ;
    wire encoder0_position_19;
    wire \quad_counter0.n13113 ;
    wire \quad_counter0.n13114 ;
    wire \quad_counter0.n13115 ;
    wire \quad_counter0.n13116 ;
    wire \quad_counter0.n13117 ;
    wire \quad_counter0.n13118 ;
    wire bfn_10_21_0_;
    wire \quad_counter0.n13119 ;
    wire \quad_counter0.n13120 ;
    wire \quad_counter0.n13121 ;
    wire \quad_counter0.n13122 ;
    wire \quad_counter0.n13123 ;
    wire \quad_counter0.n13124 ;
    wire \quad_counter0.n13125 ;
    wire bfn_10_22_0_;
    wire n12496;
    wire n12497;
    wire n12498;
    wire n12499;
    wire n12500;
    wire n2563;
    wire n13656;
    wire n403;
    wire n13_adj_631;
    wire n38;
    wire n402;
    wire n39;
    wire n2562;
    wire n5187;
    wire encoder0_position_11;
    wire n22_adj_640;
    wire encoder0_position_12;
    wire n21_adj_639;
    wire encoder0_position_13;
    wire n20_adj_638;
    wire n15_adj_633;
    wire n6_adj_624;
    wire direction_N_537;
    wire direction_N_537_cascade_;
    wire n1302;
    wire n8_adj_626;
    wire n5_adj_623;
    wire n2_adj_620;
    wire n9_adj_627;
    wire encoder0_position_scaled_5;
    wire encoder0_position_scaled_1;
    wire \quad_counter0.direction_N_540 ;
    wire encoder0_position_scaled_9;
    wire encoder0_position_scaled_20;
    wire encoder0_position_scaled_11;
    wire encoder0_position_scaled_21;
    wire encoder0_position_scaled_19;
    wire pwm_setpoint_4;
    wire encoder0_position_scaled_22;
    wire \quad_counter0.a_prev ;
    wire \quad_counter0.direction_N_536 ;
    wire n26_adj_703;
    wire bfn_10_29_0_;
    wire n25_adj_702;
    wire n13070;
    wire n24_adj_701;
    wire n13071;
    wire n23_adj_700;
    wire n13072;
    wire n22_adj_699;
    wire n13073;
    wire n21_adj_698;
    wire n13074;
    wire n20_adj_697;
    wire n13075;
    wire n19_adj_696;
    wire n13076;
    wire n13077;
    wire n18_adj_695;
    wire bfn_10_30_0_;
    wire n17_adj_694;
    wire n13078;
    wire n16_adj_693;
    wire n13079;
    wire n15_adj_692;
    wire n13080;
    wire n14_adj_691;
    wire n13081;
    wire n13_adj_690;
    wire n13082;
    wire n12_adj_689;
    wire n13083;
    wire n11_adj_688;
    wire n13084;
    wire n13085;
    wire n10_adj_687;
    wire bfn_10_31_0_;
    wire n9_adj_686;
    wire n13086;
    wire n8_adj_685;
    wire n13087;
    wire n7_adj_684;
    wire n13088;
    wire n6_adj_683;
    wire n13089;
    wire blink_counter_21;
    wire n13090;
    wire blink_counter_22;
    wire n13091;
    wire blink_counter_23;
    wire n13092;
    wire n13093;
    wire blink_counter_24;
    wire bfn_10_32_0_;
    wire n13094;
    wire blink_counter_25;
    wire n1833_cascade_;
    wire n11989;
    wire n304;
    wire n1901;
    wire bfn_11_17_0_;
    wire n1833;
    wire n1900;
    wire n12606;
    wire n1832;
    wire n1899;
    wire n12607;
    wire n1831;
    wire n1898;
    wire n12608;
    wire n1897;
    wire n12609;
    wire n1896;
    wire n12610;
    wire n12611;
    wire n12612;
    wire n12613;
    wire n1893;
    wire bfn_11_18_0_;
    wire n12614;
    wire n1891;
    wire n12615;
    wire n1890;
    wire n12616;
    wire n1889;
    wire n12617;
    wire n12618;
    wire n1887;
    wire n12619;
    wire n1886;
    wire n12620;
    wire n12621;
    wire bfn_11_19_0_;
    wire n1892;
    wire n1924;
    wire n1924_cascade_;
    wire n14438;
    wire n1822;
    wire n1822_cascade_;
    wire n14534;
    wire n1895;
    wire n1927;
    wire n1894;
    wire n1926;
    wire n1829;
    wire n1885;
    wire n1917;
    wire n30;
    wire encoder0_position_3;
    wire n316;
    wire n1888;
    wire n1851;
    wire n1920;
    wire n1987;
    wire n1920_cascade_;
    wire n1950;
    wire n2019;
    wire n1819;
    wire n16;
    wire encoder0_position_29;
    wire n404;
    wire encoder0_position_17;
    wire n16_adj_634;
    wire n7_adj_625;
    wire n3_adj_621;
    wire n2566;
    wire n7;
    wire n13662_cascade_;
    wire encoder0_position_26;
    wire n2565;
    wire encoder0_position_27;
    wire n13660_cascade_;
    wire n832_cascade_;
    wire n2564;
    wire n13658_cascade_;
    wire encoder0_position_28;
    wire encoder0_position_scaled_4;
    wire n929_cascade_;
    wire encoder0_position_30;
    wire n13654;
    wire n829_cascade_;
    wire n12027;
    wire n861_cascade_;
    wire n6;
    wire n4;
    wire n40;
    wire n5;
    wire n5_adj_682;
    wire n3;
    wire n5_adj_682_cascade_;
    wire n13653;
    wire bfn_11_24_0_;
    wire n12501;
    wire n12502;
    wire n831;
    wire n898;
    wire n12503;
    wire n830;
    wire n897;
    wire n12504;
    wire n12505;
    wire n12506;
    wire n2;
    wire n14568;
    wire n2561;
    wire n828;
    wire encoder0_position_scaled_3;
    wire encoder0_position_scaled_6;
    wire encoder0_position_scaled_2;
    wire n25_adj_597;
    wire bfn_11_26_0_;
    wire n12426;
    wire n12427;
    wire n22_adj_594;
    wire n12428;
    wire n21_adj_593;
    wire pwm_setpoint_23_N_171_4;
    wire n12429;
    wire n20_adj_592;
    wire pwm_setpoint_23_N_171_5;
    wire n12430;
    wire n12431;
    wire n18_adj_590;
    wire pwm_setpoint_23_N_171_7;
    wire n12432;
    wire n12433;
    wire n17_adj_589;
    wire pwm_setpoint_23_N_171_8;
    wire bfn_11_27_0_;
    wire n16_adj_588;
    wire n12434;
    wire n15_adj_587;
    wire n12435;
    wire n14_adj_586;
    wire pwm_setpoint_23_N_171_11;
    wire n12436;
    wire n12437;
    wire n12_adj_584;
    wire pwm_setpoint_23_N_171_13;
    wire n12438;
    wire n11_adj_583;
    wire n12439;
    wire n10_adj_582;
    wire n12440;
    wire n12441;
    wire n9_adj_581;
    wire bfn_11_28_0_;
    wire n12442;
    wire pwm_setpoint_23_N_171_18;
    wire n12443;
    wire n12444;
    wire n12445;
    wire n12446;
    wire n12447;
    wire n12448;
    wire n16_adj_664_cascade_;
    wire n24_adj_669_cascade_;
    wire n8_adj_657;
    wire n15144;
    wire pwm_setpoint_23_N_171_21;
    wire pwm_setpoint_23_N_171_9;
    wire pwm_setpoint_9;
    wire pwm_setpoint_23_N_171_14;
    wire pwm_setpoint_23_N_171_22;
    wire n9_adj_658;
    wire pwm_setpoint_8;
    wire n17_adj_665;
    wire n19_adj_666;
    wire n15178;
    wire n17_adj_665_cascade_;
    wire pwm_setpoint_23_N_171_16;
    wire n15174;
    wire pwm_setpoint_23_N_171_17;
    wire pwm_setpoint_16;
    wire pwm_setpoint_7;
    wire pwm_setpoint_23_N_171_10;
    wire pwm_setpoint_11;
    wire n15204;
    wire pwm_setpoint_17;
    wire n35_cascade_;
    wire n12_adj_661;
    wire n1825;
    wire n1825_cascade_;
    wire n14520;
    wire n1828;
    wire n1830;
    wire n1752_cascade_;
    wire n1826;
    wire n1824;
    wire n1823;
    wire n1726_cascade_;
    wire n14244_cascade_;
    wire n14250_cascade_;
    wire n14254;
    wire n1721_cascade_;
    wire n1820;
    wire n1827;
    wire n1722_cascade_;
    wire n1821;
    wire n1731_cascade_;
    wire n11991;
    wire n1801;
    wire bfn_12_20_0_;
    wire n1800;
    wire n12591;
    wire n1732;
    wire n1799;
    wire n12592;
    wire n1731;
    wire n1798;
    wire n12593;
    wire n1797;
    wire n12594;
    wire n1796;
    wire n12595;
    wire n1795;
    wire n12596;
    wire n1794;
    wire n12597;
    wire n12598;
    wire n1726;
    wire n1793;
    wire bfn_12_21_0_;
    wire n1792;
    wire n12599;
    wire n1791;
    wire n12600;
    wire n1723;
    wire n1790;
    wire n12601;
    wire n1722;
    wire n1789;
    wire n12602;
    wire n1721;
    wire n1788;
    wire n12603;
    wire n1720;
    wire n1787;
    wire n12604;
    wire n12605;
    wire n1818;
    wire n10_adj_628;
    wire n17;
    wire n303;
    wire n15;
    wire encoder0_position_18;
    wire n899;
    wire n832;
    wire n900;
    wire n833;
    wire n932_cascade_;
    wire encoder0_position_25;
    wire n8;
    wire n41;
    wire n901;
    wire n41_cascade_;
    wire n933_cascade_;
    wire n10;
    wire encoder0_position_23;
    wire encoder0_position_24;
    wire n9;
    wire n295_cascade_;
    wire n11955_cascade_;
    wire n14460;
    wire n960_cascade_;
    wire n861;
    wire n829;
    wire n896;
    wire bfn_12_25_0_;
    wire n24_adj_552;
    wire n12473;
    wire n23_adj_553;
    wire n12474;
    wire n22_adj_554;
    wire n12475;
    wire n21_adj_555;
    wire duty_4;
    wire n12476;
    wire n20_adj_556;
    wire duty_5;
    wire n12477;
    wire n19_adj_557;
    wire n12478;
    wire n18_adj_558;
    wire duty_7;
    wire n12479;
    wire n12480;
    wire n17_adj_559;
    wire duty_8;
    wire bfn_12_26_0_;
    wire n16_adj_560;
    wire duty_9;
    wire n12481;
    wire n15_adj_561;
    wire duty_10;
    wire n12482;
    wire n14_adj_562;
    wire duty_11;
    wire n12483;
    wire n13_adj_563;
    wire n12484;
    wire n12_adj_564;
    wire duty_13;
    wire n12485;
    wire n11_adj_565;
    wire duty_14;
    wire n12486;
    wire n10_adj_566;
    wire n12487;
    wire n12488;
    wire duty_16;
    wire bfn_12_27_0_;
    wire n8_adj_568;
    wire n12489;
    wire n7_adj_569;
    wire n12490;
    wire n6_adj_570;
    wire n12491;
    wire n5_adj_571;
    wire n12492;
    wire n4_adj_572;
    wire n12493;
    wire n3_adj_573;
    wire n12494;
    wire n2_adj_574;
    wire n12495;
    wire duty_17;
    wire n8_adj_580;
    wire duty_21;
    wire n4_adj_576;
    wire duty_18;
    wire n7_adj_579;
    wire pwm_setpoint_23_N_171_19;
    wire pwm_setpoint_23_N_171_20;
    wire pwm_setpoint_23_N_171_0;
    wire duty_0;
    wire pwm_setpoint_0;
    wire duty_20;
    wire n5_adj_577;
    wire pwm_setpoint_22;
    wire n45_cascade_;
    wire pwm_setpoint_20;
    wire n41_adj_678_cascade_;
    wire n40_adj_677;
    wire n45;
    wire n15223;
    wire n15165;
    wire n15243;
    wire duty_22;
    wire n3_adj_575;
    wire pwm_setpoint_19;
    wire n39_adj_676_cascade_;
    wire n15254;
    wire pwm_setpoint_21;
    wire pwm_setpoint_23_N_171_12;
    wire n39_adj_676;
    wire n41_adj_678;
    wire n15091;
    wire n4_adj_655;
    wire pwm_setpoint_12;
    wire n25_adj_670;
    wire n15110;
    wire n23_adj_668;
    wire n25_adj_670_cascade_;
    wire n43;
    wire n15146;
    wire n13_adj_662;
    wire n15_adj_663;
    wire n15229;
    wire duty_12;
    wire n13_adj_585;
    wire n31_adj_674_cascade_;
    wire n15230;
    wire n15237;
    wire n15195_cascade_;
    wire n15241;
    wire n15097;
    wire n10_adj_659;
    wire n30_adj_673;
    wire n33_adj_675;
    wire n15104;
    wire n31_adj_674;
    wire n35;
    wire n15247;
    wire n15099_cascade_;
    wire n15220;
    wire pwm_setpoint_18;
    wire n15257_cascade_;
    wire n37;
    wire n15258;
    wire bfn_13_17_0_;
    wire n1700;
    wire n12577;
    wire n1699;
    wire n12578;
    wire n12579;
    wire n12580;
    wire n12581;
    wire n12582;
    wire n1694;
    wire n12583;
    wire n12584;
    wire bfn_13_18_0_;
    wire n12585;
    wire n1691;
    wire n12586;
    wire n1690;
    wire n12587;
    wire n1689;
    wire n12588;
    wire n1688;
    wire n12589;
    wire n12590;
    wire n1719;
    wire n1695;
    wire n1727;
    wire n1696;
    wire n1653_cascade_;
    wire n1728;
    wire n1697;
    wire n1692;
    wire n1724;
    wire n1693_adj_614;
    wire n1725;
    wire n15611;
    wire n1625_adj_605;
    wire n1625_adj_605_cascade_;
    wire n1698;
    wire n1730;
    wire n1730_cascade_;
    wire n1729;
    wire n14514;
    wire n11_adj_629;
    wire n1701;
    wire n1653;
    wire n1733;
    wire n1752;
    wire n15630;
    wire n1621_adj_601;
    wire ENCODER0_B_N;
    wire encoder0_position_1;
    wire n32_adj_650;
    wire encoder0_position_16;
    wire n17_adj_635;
    wire n1129_cascade_;
    wire n11933_cascade_;
    wire n13728_cascade_;
    wire n1059_cascade_;
    wire n1132_cascade_;
    wire n295;
    wire n1001;
    wire bfn_13_24_0_;
    wire n933;
    wire n1000;
    wire n12507;
    wire n932;
    wire n999;
    wire n12508;
    wire n931;
    wire n998;
    wire n12509;
    wire n930;
    wire n997;
    wire n12510;
    wire n929;
    wire n996;
    wire n12511;
    wire n928;
    wire n995;
    wire n12512;
    wire n960;
    wire n927;
    wire n12513;
    wire encoder0_position_scaled_0;
    wire n25_adj_551;
    wire n11872_cascade_;
    wire n14034_cascade_;
    wire n14116_cascade_;
    wire n10_adj_598;
    wire pwm_setpoint_23_N_171_2;
    wire pwm_setpoint_23_N_171_3;
    wire duty_3;
    wire n10_adj_681;
    wire n16_adj_710_cascade_;
    wire n15_adj_711;
    wire duty_2;
    wire n23_adj_595;
    wire duty_15;
    wire pwm_setpoint_23_N_171_15;
    wire pwm_setpoint_15;
    wire \quad_counter0.a_new_0 ;
    wire \quad_counter0.b_new_0 ;
    wire a_new_1;
    wire \quad_counter0.a_prev_N_543 ;
    wire \quad_counter0.b_new_1 ;
    wire \quad_counter0.debounce_cnt ;
    wire \quad_counter0.a_prev_N_543_cascade_ ;
    wire b_prev;
    wire n15121;
    wire pwm_setpoint_23_N_171_6;
    wire pwm_setpoint_6;
    wire pwm_setpoint_2;
    wire pwm_setpoint_3;
    wire duty_19;
    wire n6_adj_578;
    wire \PWM.n13991 ;
    wire n4_adj_599;
    wire commutation_state_prev_1;
    wire n5137;
    wire dti;
    wire n5201_cascade_;
    wire pwm_setpoint_13;
    wire n27_adj_671;
    wire \PWM.n17 ;
    wire \PWM.n26_cascade_ ;
    wire \PWM.n27 ;
    wire \PWM.n29_cascade_ ;
    wire \PWM.n28 ;
    wire commutation_state_prev_2;
    wire h2;
    wire h3;
    wire h1;
    wire n6_adj_721;
    wire commutation_state_7__N_261;
    wire pwm_setpoint_5;
    wire n11_adj_660;
    wire pwm_setpoint_14;
    wire n29_adj_672;
    wire n21_adj_667;
    wire pwm_setpoint_10;
    wire n21_adj_667_cascade_;
    wire n6_adj_656;
    wire n15203;
    wire n14420_cascade_;
    wire n1630_adj_610;
    wire n1629_adj_609;
    wire n1630_adj_610_cascade_;
    wire n1624_adj_604;
    wire n14502;
    wire n1623_adj_603;
    wire n1624_adj_604_cascade_;
    wire n13748;
    wire n14508;
    wire n1627_adj_607;
    wire n1523_cascade_;
    wire n1622_adj_602;
    wire n14426;
    wire n14428_cascade_;
    wire n1554_cascade_;
    wire n1427_cascade_;
    wire n1628_adj_608;
    wire n11;
    wire encoder0_position_22;
    wire n1626_adj_606;
    wire duty_6;
    wire n19_adj_591;
    wire bfn_14_20_0_;
    wire n12541;
    wire n12542;
    wire n12543;
    wire n12544;
    wire n1396;
    wire n12545;
    wire n1395;
    wire n12546;
    wire n12547;
    wire n12548;
    wire bfn_14_21_0_;
    wire n1392;
    wire n12549;
    wire n12550;
    wire n12551;
    wire n15553;
    wire n1401;
    wire n12019;
    wire n14406_cascade_;
    wire n14464;
    wire n1233_cascade_;
    wire n297;
    wire n1201;
    wire bfn_14_23_0_;
    wire n1133;
    wire n1200;
    wire n12522;
    wire n12523;
    wire n1131;
    wire n1198;
    wire n12524;
    wire n1130;
    wire n1197;
    wire n12525;
    wire n12526;
    wire n12527;
    wire n12528;
    wire n12529;
    wire bfn_14_24_0_;
    wire n12530;
    wire n15522;
    wire n13;
    wire encoder0_position_20;
    wire n1125;
    wire n20_adj_618_cascade_;
    wire n13197;
    wire n13197_cascade_;
    wire n24_adj_653;
    wire direction_N_342_cascade_;
    wire direction_N_342;
    wire n13675;
    wire n23_adj_709_cascade_;
    wire n25_adj_707;
    wire direction_N_340;
    wire n24_adj_708;
    wire n23_adj_654;
    wire pwm_setpoint_23_N_171_1;
    wire pwm_setpoint_1;
    wire n16_adj_679_cascade_;
    wire n15_adj_680;
    wire n25_adj_652;
    wire n16_adj_619_cascade_;
    wire n22_adj_617;
    wire n24_adj_616;
    wire encoder0_position_scaled_16;
    wire n9_adj_567;
    wire duty_1;
    wire n24_adj_596;
    wire pwm_setpoint_23__N_195;
    wire pwm_counter_0;
    wire bfn_14_28_0_;
    wire pwm_counter_1;
    wire \PWM.n13022 ;
    wire pwm_counter_2;
    wire \PWM.n13023 ;
    wire pwm_counter_3;
    wire \PWM.n13024 ;
    wire pwm_counter_4;
    wire \PWM.n13025 ;
    wire pwm_counter_5;
    wire \PWM.n13026 ;
    wire pwm_counter_6;
    wire \PWM.n13027 ;
    wire pwm_counter_7;
    wire \PWM.n13028 ;
    wire \PWM.n13029 ;
    wire pwm_counter_8;
    wire bfn_14_29_0_;
    wire pwm_counter_9;
    wire \PWM.n13030 ;
    wire pwm_counter_10;
    wire \PWM.n13031 ;
    wire pwm_counter_11;
    wire \PWM.n13032 ;
    wire pwm_counter_12;
    wire \PWM.n13033 ;
    wire pwm_counter_13;
    wire \PWM.n13034 ;
    wire pwm_counter_14;
    wire \PWM.n13035 ;
    wire pwm_counter_15;
    wire \PWM.n13036 ;
    wire \PWM.n13037 ;
    wire pwm_counter_16;
    wire bfn_14_30_0_;
    wire pwm_counter_17;
    wire \PWM.n13038 ;
    wire pwm_counter_18;
    wire \PWM.n13039 ;
    wire pwm_counter_19;
    wire \PWM.n13040 ;
    wire pwm_counter_20;
    wire \PWM.n13041 ;
    wire pwm_counter_21;
    wire \PWM.n13042 ;
    wire pwm_counter_22;
    wire \PWM.n13043 ;
    wire \PWM.n13044 ;
    wire \PWM.n13045 ;
    wire bfn_14_31_0_;
    wire \PWM.n13046 ;
    wire \PWM.n13047 ;
    wire \PWM.n13048 ;
    wire \PWM.n13049 ;
    wire \PWM.n13050 ;
    wire \PWM.n13051 ;
    wire \PWM.n13052 ;
    wire \PWM.pwm_counter_31__N_407 ;
    wire pwm_counter_24;
    wire pwm_counter_29;
    wire pwm_counter_27;
    wire pwm_counter_26;
    wire pwm_counter_30;
    wire pwm_counter_25;
    wire n12_adj_615_cascade_;
    wire pwm_counter_28;
    wire n1631_adj_611;
    wire n1554;
    wire n1632_adj_612;
    wire n302;
    wire n1632_adj_612_cascade_;
    wire n1633_adj_613;
    wire n11919;
    wire n1393;
    wire n1425_cascade_;
    wire n14484;
    wire n14490_cascade_;
    wire n1455_cascade_;
    wire n1531_cascade_;
    wire n11997;
    wire n1455;
    wire n1394;
    wire n1391;
    wire n299;
    wire n11925_cascade_;
    wire n1398;
    wire n1430_cascade_;
    wire n13739;
    wire n13720;
    wire n1400;
    wire n1356_cascade_;
    wire n1333;
    wire n1432_cascade_;
    wire n11923;
    wire n1328;
    wire n1328_cascade_;
    wire n14414;
    wire n1327;
    wire n1331;
    wire n1332;
    wire n1399;
    wire n1332_cascade_;
    wire n1329;
    wire n11927;
    wire n13723_cascade_;
    wire n1257_cascade_;
    wire n1325;
    wire n12;
    wire encoder0_position_31;
    wire n1326;
    wire n1195;
    wire n1227_cascade_;
    wire n14476;
    wire n1199;
    wire n1132;
    wire n1127;
    wire n1194;
    wire n1127_cascade_;
    wire n1126;
    wire n1193;
    wire n1225_cascade_;
    wire n1324;
    wire n1129;
    wire n1196;
    wire n1158;
    wire n1059;
    wire n1128;
    wire bfn_15_25_0_;
    wire n1693;
    wire encoder0_position_target_0;
    wire n12449;
    wire encoder0_position_target_1;
    wire n12450;
    wire encoder0_position_target_2;
    wire n12451;
    wire encoder0_position_target_3;
    wire n12452;
    wire encoder0_position_target_4;
    wire n12453;
    wire encoder0_position_target_5;
    wire n12454;
    wire encoder0_position_target_6;
    wire n12455;
    wire n12456;
    wire encoder0_position_target_7;
    wire bfn_15_26_0_;
    wire encoder0_position_target_8;
    wire n12457;
    wire encoder0_position_target_9;
    wire n12458;
    wire encoder0_position_target_10;
    wire n12459;
    wire encoder0_position_target_11;
    wire n12460;
    wire encoder0_position_target_12;
    wire n12461;
    wire encoder0_position_target_13;
    wire n12462;
    wire encoder0_position_target_14;
    wire n12463;
    wire n12464;
    wire encoder0_position_target_15;
    wire bfn_15_27_0_;
    wire encoder0_position_target_16;
    wire n12465;
    wire encoder0_position_target_17;
    wire n12466;
    wire encoder0_position_target_18;
    wire n12467;
    wire encoder0_position_target_19;
    wire n12468;
    wire encoder0_position_target_20;
    wire n12469;
    wire encoder0_position_target_21;
    wire n12470;
    wire encoder0_position_target_22;
    wire n12471;
    wire n12472;
    wire direction_c;
    wire bfn_15_28_0_;
    wire encoder0_position_target_23;
    wire pwm_setpoint_23;
    wire pwm_counter_23;
    wire n15245;
    wire pwm_counter_31;
    wire n5180;
    wire n5182;
    wire duty_23;
    wire n300;
    wire n1501;
    wire bfn_16_17_0_;
    wire n1433;
    wire n1500;
    wire n12552;
    wire n1432;
    wire n1499;
    wire n12553;
    wire n1431;
    wire n1498;
    wire n12554;
    wire n1430;
    wire n1497;
    wire n12555;
    wire n1496;
    wire n12556;
    wire n1428;
    wire n1495;
    wire n12557;
    wire n1427;
    wire n1494;
    wire n12558;
    wire n12559;
    wire n1426;
    wire n1493;
    wire bfn_16_18_0_;
    wire n1425;
    wire n1492;
    wire n12560;
    wire n1424;
    wire n1491;
    wire n12561;
    wire n1423;
    wire n1490;
    wire n12562;
    wire n15572;
    wire n1422;
    wire n12563;
    wire n301;
    wire n1601;
    wire bfn_16_19_0_;
    wire n1533;
    wire n1600;
    wire n12564;
    wire n1532;
    wire n1599;
    wire n12565;
    wire n1531;
    wire n1598;
    wire n12566;
    wire n1530;
    wire n1597;
    wire n12567;
    wire n1529;
    wire n1596;
    wire n12568;
    wire n1528;
    wire n1595;
    wire n12569;
    wire n1527;
    wire n1594;
    wire n12570;
    wire n12571;
    wire n1526;
    wire n1593;
    wire bfn_16_20_0_;
    wire n1525;
    wire n1592;
    wire n12572;
    wire n1524;
    wire n1591;
    wire n12573;
    wire n1523;
    wire n1590;
    wire n12574;
    wire n1522;
    wire n1589;
    wire n12575;
    wire n1521;
    wire n15591;
    wire n12576;
    wire n1620_adj_600;
    wire encoder0_position_21;
    wire n12_adj_630;
    wire n1397;
    wire n1356;
    wire n1429;
    wire n298;
    wire n1301;
    wire bfn_16_21_0_;
    wire n1233;
    wire n1300;
    wire n12531;
    wire n1232;
    wire n1299;
    wire n12532;
    wire n12533;
    wire n1230;
    wire n1297;
    wire n12534;
    wire n1229;
    wire n1296;
    wire n12535;
    wire n1228;
    wire n1295;
    wire n12536;
    wire n1227;
    wire n1294;
    wire n12537;
    wire n12538;
    wire n1226;
    wire n1293;
    wire bfn_16_22_0_;
    wire n1225;
    wire n1292;
    wire n12539;
    wire n15537;
    wire n1224;
    wire n12540;
    wire n1323;
    wire n1298;
    wire n1231;
    wire n1257;
    wire n1330;
    wire n296;
    wire n1101;
    wire bfn_16_23_0_;
    wire n1033;
    wire n1100;
    wire n12514;
    wire n1032;
    wire n1099;
    wire n12515;
    wire n1031;
    wire n1098;
    wire n12516;
    wire n1030;
    wire n1097;
    wire n12517;
    wire n1029;
    wire n1096;
    wire n12518;
    wire n1028;
    wire n1095;
    wire n12519;
    wire n1027;
    wire n1094;
    wire n12520;
    wire n12521;
    wire CONSTANT_ONE_NET;
    wire n1026;
    wire bfn_16_24_0_;
    wire n1093;
    wire sweep_counter_0;
    wire bfn_16_25_0_;
    wire sweep_counter_1;
    wire n13053;
    wire sweep_counter_2;
    wire n13054;
    wire sweep_counter_3;
    wire n13055;
    wire sweep_counter_4;
    wire n13056;
    wire sweep_counter_5;
    wire n13057;
    wire sweep_counter_6;
    wire n13058;
    wire sweep_counter_7;
    wire n13059;
    wire n13060;
    wire bfn_16_26_0_;
    wire sweep_counter_9;
    wire n13061;
    wire sweep_counter_10;
    wire n13062;
    wire sweep_counter_11;
    wire n13063;
    wire n13064;
    wire n13065;
    wire n13066;
    wire sweep_counter_15;
    wire n13067;
    wire n13068;
    wire sweep_counter_16;
    wire bfn_16_27_0_;
    wire n13069;
    wire n5215;
    wire sweep_counter_8;
    wire sweep_counter_14;
    wire sweep_counter_13;
    wire sweep_counter_17;
    wire n6_adj_712_cascade_;
    wire sweep_counter_12;
    wire n13968;
    wire GHC;
    wire INHC_c_0;
    wire GHB;
    wire INHB_c_0;
    wire INLA_c_0;
    wire INLB_c_0;
    wire commutation_state_0;
    wire commutation_state_2;
    wire dir;
    wire commutation_state_1;
    wire INLC_c_0;
    wire CLK_N;
    wire n5201;
    wire n5253;
    wire GHA;
    wire pwm_out;
    wire INHA_c_0;
    wire _gnd_net_;

    defparam CS_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CS_CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CS_CLK_pad_iopad (
            .OE(N__56752),
            .DIN(N__56751),
            .DOUT(N__56750),
            .PACKAGEPIN(CS_CLK));
    defparam CS_CLK_pad_preio.PIN_TYPE=6'b011001;
    defparam CS_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CS_CLK_pad_preio (
            .PADOEN(N__56752),
            .PADOUT(N__56751),
            .PADIN(N__56750),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam CS_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CS_pad_iopad.PULLUP=1'b0;
    IO_PAD CS_pad_iopad (
            .OE(N__56743),
            .DIN(N__56742),
            .DOUT(N__56741),
            .PACKAGEPIN(CS));
    defparam CS_pad_preio.PIN_TYPE=6'b011001;
    defparam CS_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CS_pad_preio (
            .PADOEN(N__56743),
            .PADOUT(N__56742),
            .PADIN(N__56741),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam DE_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DE_pad_iopad.PULLUP=1'b0;
    IO_PAD DE_pad_iopad (
            .OE(N__56734),
            .DIN(N__56733),
            .DOUT(N__56732),
            .PACKAGEPIN(DE));
    defparam DE_pad_preio.PIN_TYPE=6'b011001;
    defparam DE_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DE_pad_preio (
            .PADOEN(N__56734),
            .PADOUT(N__56733),
            .PADIN(N__56732),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam ENCODER0_A_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ENCODER0_A_pad_iopad.PULLUP=1'b0;
    IO_PAD ENCODER0_A_pad_iopad (
            .OE(N__56725),
            .DIN(N__56724),
            .DOUT(N__56723),
            .PACKAGEPIN(ENCODER0_A));
    defparam ENCODER0_A_pad_preio.PIN_TYPE=6'b000001;
    defparam ENCODER0_A_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ENCODER0_A_pad_preio (
            .PADOEN(N__56725),
            .PADOUT(N__56724),
            .PADIN(N__56723),
            .CLOCKENABLE(),
            .DIN0(ENCODER0_A_N),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam ENCODER0_B_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ENCODER0_B_pad_iopad.PULLUP=1'b0;
    IO_PAD ENCODER0_B_pad_iopad (
            .OE(N__56716),
            .DIN(N__56715),
            .DOUT(N__56714),
            .PACKAGEPIN(ENCODER0_B));
    defparam ENCODER0_B_pad_preio.PIN_TYPE=6'b000001;
    defparam ENCODER0_B_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ENCODER0_B_pad_preio (
            .PADOEN(N__56716),
            .PADOUT(N__56715),
            .PADIN(N__56714),
            .CLOCKENABLE(),
            .DIN0(ENCODER0_B_N),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHA_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHA_pad_iopad.PULLUP=1'b0;
    IO_PAD INHA_pad_iopad (
            .OE(N__56707),
            .DIN(N__56706),
            .DOUT(N__56705),
            .PACKAGEPIN(INHA));
    defparam INHA_pad_preio.PIN_TYPE=6'b011001;
    defparam INHA_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHA_pad_preio (
            .PADOEN(N__56707),
            .PADOUT(N__56706),
            .PADIN(N__56705),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__55974),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHB_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHB_pad_iopad.PULLUP=1'b0;
    IO_PAD INHB_pad_iopad (
            .OE(N__56698),
            .DIN(N__56697),
            .DOUT(N__56696),
            .PACKAGEPIN(INHB));
    defparam INHB_pad_preio.PIN_TYPE=6'b011001;
    defparam INHB_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHB_pad_preio (
            .PADOEN(N__56698),
            .PADOUT(N__56697),
            .PADIN(N__56696),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__56565),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INHC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INHC_pad_iopad.PULLUP=1'b0;
    IO_PAD INHC_pad_iopad (
            .OE(N__56689),
            .DIN(N__56688),
            .DOUT(N__56687),
            .PACKAGEPIN(INHC));
    defparam INHC_pad_preio.PIN_TYPE=6'b011001;
    defparam INHC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INHC_pad_preio (
            .PADOEN(N__56689),
            .PADOUT(N__56688),
            .PADIN(N__56687),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__55728),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLA_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLA_pad_iopad.PULLUP=1'b0;
    IO_PAD INLA_pad_iopad (
            .OE(N__56680),
            .DIN(N__56679),
            .DOUT(N__56678),
            .PACKAGEPIN(INLA));
    defparam INLA_pad_preio.PIN_TYPE=6'b011001;
    defparam INLA_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLA_pad_preio (
            .PADOEN(N__56680),
            .PADOUT(N__56679),
            .PADIN(N__56678),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__56553),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLB_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLB_pad_iopad.PULLUP=1'b0;
    IO_PAD INLB_pad_iopad (
            .OE(N__56671),
            .DIN(N__56670),
            .DOUT(N__56669),
            .PACKAGEPIN(INLB));
    defparam INLB_pad_preio.PIN_TYPE=6'b011001;
    defparam INLB_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLB_pad_preio (
            .PADOEN(N__56671),
            .PADOUT(N__56670),
            .PADIN(N__56669),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__56538),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam INLC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam INLC_pad_iopad.PULLUP=1'b0;
    IO_PAD INLC_pad_iopad (
            .OE(N__56662),
            .DIN(N__56661),
            .DOUT(N__56660),
            .PACKAGEPIN(INLC));
    defparam INLC_pad_preio.PIN_TYPE=6'b011001;
    defparam INLC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO INLC_pad_preio (
            .PADOEN(N__56662),
            .PADOUT(N__56661),
            .PADIN(N__56660),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__56277),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__56653),
            .DIN(N__56652),
            .DOUT(N__56651),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__56653),
            .PADOUT(N__56652),
            .PADIN(N__56651),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__39138),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam NEOPXL_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam NEOPXL_pad_iopad.PULLUP=1'b0;
    IO_PAD NEOPXL_pad_iopad (
            .OE(N__56644),
            .DIN(N__56643),
            .DOUT(N__56642),
            .PACKAGEPIN(NEOPXL));
    defparam NEOPXL_pad_preio.PIN_TYPE=6'b011001;
    defparam NEOPXL_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO NEOPXL_pad_preio (
            .PADOEN(N__56644),
            .PADOUT(N__56643),
            .PADIN(N__56642),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam TX_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TX_pad_iopad.PULLUP=1'b0;
    IO_PAD TX_pad_iopad (
            .OE(N__56635),
            .DIN(N__56634),
            .DOUT(N__56633),
            .PACKAGEPIN(TX));
    defparam TX_pad_preio.PIN_TYPE=6'b011001;
    defparam TX_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO TX_pad_preio (
            .PADOEN(N__56635),
            .PADOUT(N__56634),
            .PADIN(N__56633),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__56626),
            .DIN(N__56625),
            .DOUT(N__56624),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__56626),
            .PADOUT(N__56625),
            .PADIN(N__56624),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall1_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall1_input_iopad.PULLUP=1'b1;
    IO_PAD hall1_input_iopad (
            .OE(N__56617),
            .DIN(N__56616),
            .DOUT(N__56615),
            .PACKAGEPIN(HALL1));
    defparam hall1_input_preio.PIN_TYPE=6'b000000;
    defparam hall1_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall1_input_preio (
            .PADOEN(N__56617),
            .PADOUT(N__56616),
            .PADIN(N__56615),
            .CLOCKENABLE(VCCG0),
            .DIN0(\debounce.reg_A_2 ),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(N__56204),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall2_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall2_input_iopad.PULLUP=1'b1;
    IO_PAD hall2_input_iopad (
            .OE(N__56608),
            .DIN(N__56607),
            .DOUT(N__56606),
            .PACKAGEPIN(HALL2));
    defparam hall2_input_preio.PIN_TYPE=6'b000000;
    defparam hall2_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall2_input_preio (
            .PADOEN(N__56608),
            .PADOUT(N__56607),
            .PADIN(N__56606),
            .CLOCKENABLE(VCCG0),
            .DIN0(\debounce.reg_A_1 ),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(N__56200),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam hall3_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam hall3_input_iopad.PULLUP=1'b1;
    IO_PAD hall3_input_iopad (
            .OE(N__56599),
            .DIN(N__56598),
            .DOUT(N__56597),
            .PACKAGEPIN(HALL3));
    defparam hall3_input_preio.PIN_TYPE=6'b000000;
    defparam hall3_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO hall3_input_preio (
            .PADOEN(N__56599),
            .PADOUT(N__56598),
            .PADIN(N__56597),
            .CLOCKENABLE(VCCG0),
            .DIN0(\debounce.reg_A_0 ),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(N__56200),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__56590),
            .DIN(N__56589),
            .DOUT(N__56588),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__56590),
            .PADOUT(N__56589),
            .PADIN(N__56588),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__13452 (
            .O(N__56571),
            .I(N__56568));
    LocalMux I__13451 (
            .O(N__56568),
            .I(GHB));
    IoInMux I__13450 (
            .O(N__56565),
            .I(N__56562));
    LocalMux I__13449 (
            .O(N__56562),
            .I(N__56559));
    Span12Mux_s0_v I__13448 (
            .O(N__56559),
            .I(N__56556));
    Odrv12 I__13447 (
            .O(N__56556),
            .I(INHB_c_0));
    IoInMux I__13446 (
            .O(N__56553),
            .I(N__56550));
    LocalMux I__13445 (
            .O(N__56550),
            .I(N__56547));
    Span4Mux_s1_v I__13444 (
            .O(N__56547),
            .I(N__56544));
    Span4Mux_h I__13443 (
            .O(N__56544),
            .I(N__56541));
    Odrv4 I__13442 (
            .O(N__56541),
            .I(INLA_c_0));
    IoInMux I__13441 (
            .O(N__56538),
            .I(N__56535));
    LocalMux I__13440 (
            .O(N__56535),
            .I(N__56532));
    Span4Mux_s1_v I__13439 (
            .O(N__56532),
            .I(N__56529));
    Span4Mux_h I__13438 (
            .O(N__56529),
            .I(N__56526));
    Odrv4 I__13437 (
            .O(N__56526),
            .I(INLB_c_0));
    InMux I__13436 (
            .O(N__56523),
            .I(N__56497));
    InMux I__13435 (
            .O(N__56522),
            .I(N__56497));
    InMux I__13434 (
            .O(N__56521),
            .I(N__56497));
    InMux I__13433 (
            .O(N__56520),
            .I(N__56497));
    InMux I__13432 (
            .O(N__56519),
            .I(N__56497));
    InMux I__13431 (
            .O(N__56518),
            .I(N__56494));
    InMux I__13430 (
            .O(N__56517),
            .I(N__56491));
    InMux I__13429 (
            .O(N__56516),
            .I(N__56488));
    InMux I__13428 (
            .O(N__56515),
            .I(N__56485));
    InMux I__13427 (
            .O(N__56514),
            .I(N__56476));
    InMux I__13426 (
            .O(N__56513),
            .I(N__56476));
    InMux I__13425 (
            .O(N__56512),
            .I(N__56476));
    InMux I__13424 (
            .O(N__56511),
            .I(N__56476));
    InMux I__13423 (
            .O(N__56510),
            .I(N__56469));
    InMux I__13422 (
            .O(N__56509),
            .I(N__56469));
    InMux I__13421 (
            .O(N__56508),
            .I(N__56469));
    LocalMux I__13420 (
            .O(N__56497),
            .I(N__56466));
    LocalMux I__13419 (
            .O(N__56494),
            .I(N__56461));
    LocalMux I__13418 (
            .O(N__56491),
            .I(N__56461));
    LocalMux I__13417 (
            .O(N__56488),
            .I(N__56450));
    LocalMux I__13416 (
            .O(N__56485),
            .I(N__56450));
    LocalMux I__13415 (
            .O(N__56476),
            .I(N__56450));
    LocalMux I__13414 (
            .O(N__56469),
            .I(N__56450));
    Span12Mux_v I__13413 (
            .O(N__56466),
            .I(N__56450));
    Span4Mux_h I__13412 (
            .O(N__56461),
            .I(N__56447));
    Odrv12 I__13411 (
            .O(N__56450),
            .I(commutation_state_0));
    Odrv4 I__13410 (
            .O(N__56447),
            .I(commutation_state_0));
    CascadeMux I__13409 (
            .O(N__56442),
            .I(N__56436));
    CascadeMux I__13408 (
            .O(N__56441),
            .I(N__56433));
    CascadeMux I__13407 (
            .O(N__56440),
            .I(N__56428));
    CascadeMux I__13406 (
            .O(N__56439),
            .I(N__56425));
    InMux I__13405 (
            .O(N__56436),
            .I(N__56416));
    InMux I__13404 (
            .O(N__56433),
            .I(N__56416));
    InMux I__13403 (
            .O(N__56432),
            .I(N__56416));
    InMux I__13402 (
            .O(N__56431),
            .I(N__56416));
    InMux I__13401 (
            .O(N__56428),
            .I(N__56413));
    InMux I__13400 (
            .O(N__56425),
            .I(N__56410));
    LocalMux I__13399 (
            .O(N__56416),
            .I(N__56407));
    LocalMux I__13398 (
            .O(N__56413),
            .I(N__56398));
    LocalMux I__13397 (
            .O(N__56410),
            .I(N__56398));
    Span4Mux_s2_v I__13396 (
            .O(N__56407),
            .I(N__56395));
    CascadeMux I__13395 (
            .O(N__56406),
            .I(N__56392));
    CascadeMux I__13394 (
            .O(N__56405),
            .I(N__56389));
    InMux I__13393 (
            .O(N__56404),
            .I(N__56384));
    InMux I__13392 (
            .O(N__56403),
            .I(N__56384));
    Span4Mux_s2_v I__13391 (
            .O(N__56398),
            .I(N__56381));
    Span4Mux_h I__13390 (
            .O(N__56395),
            .I(N__56378));
    InMux I__13389 (
            .O(N__56392),
            .I(N__56373));
    InMux I__13388 (
            .O(N__56389),
            .I(N__56373));
    LocalMux I__13387 (
            .O(N__56384),
            .I(commutation_state_2));
    Odrv4 I__13386 (
            .O(N__56381),
            .I(commutation_state_2));
    Odrv4 I__13385 (
            .O(N__56378),
            .I(commutation_state_2));
    LocalMux I__13384 (
            .O(N__56373),
            .I(commutation_state_2));
    CascadeMux I__13383 (
            .O(N__56364),
            .I(N__56360));
    CascadeMux I__13382 (
            .O(N__56363),
            .I(N__56356));
    InMux I__13381 (
            .O(N__56360),
            .I(N__56344));
    InMux I__13380 (
            .O(N__56359),
            .I(N__56344));
    InMux I__13379 (
            .O(N__56356),
            .I(N__56344));
    InMux I__13378 (
            .O(N__56355),
            .I(N__56344));
    InMux I__13377 (
            .O(N__56354),
            .I(N__56341));
    InMux I__13376 (
            .O(N__56353),
            .I(N__56338));
    LocalMux I__13375 (
            .O(N__56344),
            .I(N__56333));
    LocalMux I__13374 (
            .O(N__56341),
            .I(N__56333));
    LocalMux I__13373 (
            .O(N__56338),
            .I(dir));
    Odrv12 I__13372 (
            .O(N__56333),
            .I(dir));
    InMux I__13371 (
            .O(N__56328),
            .I(N__56316));
    InMux I__13370 (
            .O(N__56327),
            .I(N__56307));
    InMux I__13369 (
            .O(N__56326),
            .I(N__56307));
    InMux I__13368 (
            .O(N__56325),
            .I(N__56307));
    InMux I__13367 (
            .O(N__56324),
            .I(N__56307));
    InMux I__13366 (
            .O(N__56323),
            .I(N__56304));
    InMux I__13365 (
            .O(N__56322),
            .I(N__56297));
    InMux I__13364 (
            .O(N__56321),
            .I(N__56297));
    InMux I__13363 (
            .O(N__56320),
            .I(N__56297));
    InMux I__13362 (
            .O(N__56319),
            .I(N__56294));
    LocalMux I__13361 (
            .O(N__56316),
            .I(N__56287));
    LocalMux I__13360 (
            .O(N__56307),
            .I(N__56287));
    LocalMux I__13359 (
            .O(N__56304),
            .I(N__56287));
    LocalMux I__13358 (
            .O(N__56297),
            .I(N__56284));
    LocalMux I__13357 (
            .O(N__56294),
            .I(commutation_state_1));
    Odrv12 I__13356 (
            .O(N__56287),
            .I(commutation_state_1));
    Odrv4 I__13355 (
            .O(N__56284),
            .I(commutation_state_1));
    IoInMux I__13354 (
            .O(N__56277),
            .I(N__56274));
    LocalMux I__13353 (
            .O(N__56274),
            .I(N__56271));
    Span12Mux_s6_v I__13352 (
            .O(N__56271),
            .I(N__56268));
    Span12Mux_h I__13351 (
            .O(N__56268),
            .I(N__56265));
    Odrv12 I__13350 (
            .O(N__56265),
            .I(INLC_c_0));
    ClkMux I__13349 (
            .O(N__56262),
            .I(N__56070));
    ClkMux I__13348 (
            .O(N__56261),
            .I(N__56070));
    ClkMux I__13347 (
            .O(N__56260),
            .I(N__56070));
    ClkMux I__13346 (
            .O(N__56259),
            .I(N__56070));
    ClkMux I__13345 (
            .O(N__56258),
            .I(N__56070));
    ClkMux I__13344 (
            .O(N__56257),
            .I(N__56070));
    ClkMux I__13343 (
            .O(N__56256),
            .I(N__56070));
    ClkMux I__13342 (
            .O(N__56255),
            .I(N__56070));
    ClkMux I__13341 (
            .O(N__56254),
            .I(N__56070));
    ClkMux I__13340 (
            .O(N__56253),
            .I(N__56070));
    ClkMux I__13339 (
            .O(N__56252),
            .I(N__56070));
    ClkMux I__13338 (
            .O(N__56251),
            .I(N__56070));
    ClkMux I__13337 (
            .O(N__56250),
            .I(N__56070));
    ClkMux I__13336 (
            .O(N__56249),
            .I(N__56070));
    ClkMux I__13335 (
            .O(N__56248),
            .I(N__56070));
    ClkMux I__13334 (
            .O(N__56247),
            .I(N__56070));
    ClkMux I__13333 (
            .O(N__56246),
            .I(N__56070));
    ClkMux I__13332 (
            .O(N__56245),
            .I(N__56070));
    ClkMux I__13331 (
            .O(N__56244),
            .I(N__56070));
    ClkMux I__13330 (
            .O(N__56243),
            .I(N__56070));
    ClkMux I__13329 (
            .O(N__56242),
            .I(N__56070));
    ClkMux I__13328 (
            .O(N__56241),
            .I(N__56070));
    ClkMux I__13327 (
            .O(N__56240),
            .I(N__56070));
    ClkMux I__13326 (
            .O(N__56239),
            .I(N__56070));
    ClkMux I__13325 (
            .O(N__56238),
            .I(N__56070));
    ClkMux I__13324 (
            .O(N__56237),
            .I(N__56070));
    ClkMux I__13323 (
            .O(N__56236),
            .I(N__56070));
    ClkMux I__13322 (
            .O(N__56235),
            .I(N__56070));
    ClkMux I__13321 (
            .O(N__56234),
            .I(N__56070));
    ClkMux I__13320 (
            .O(N__56233),
            .I(N__56070));
    ClkMux I__13319 (
            .O(N__56232),
            .I(N__56070));
    ClkMux I__13318 (
            .O(N__56231),
            .I(N__56070));
    ClkMux I__13317 (
            .O(N__56230),
            .I(N__56070));
    ClkMux I__13316 (
            .O(N__56229),
            .I(N__56070));
    ClkMux I__13315 (
            .O(N__56228),
            .I(N__56070));
    ClkMux I__13314 (
            .O(N__56227),
            .I(N__56070));
    ClkMux I__13313 (
            .O(N__56226),
            .I(N__56070));
    ClkMux I__13312 (
            .O(N__56225),
            .I(N__56070));
    ClkMux I__13311 (
            .O(N__56224),
            .I(N__56070));
    ClkMux I__13310 (
            .O(N__56223),
            .I(N__56070));
    ClkMux I__13309 (
            .O(N__56222),
            .I(N__56070));
    ClkMux I__13308 (
            .O(N__56221),
            .I(N__56070));
    ClkMux I__13307 (
            .O(N__56220),
            .I(N__56070));
    ClkMux I__13306 (
            .O(N__56219),
            .I(N__56070));
    ClkMux I__13305 (
            .O(N__56218),
            .I(N__56070));
    ClkMux I__13304 (
            .O(N__56217),
            .I(N__56070));
    ClkMux I__13303 (
            .O(N__56216),
            .I(N__56070));
    ClkMux I__13302 (
            .O(N__56215),
            .I(N__56070));
    ClkMux I__13301 (
            .O(N__56214),
            .I(N__56070));
    ClkMux I__13300 (
            .O(N__56213),
            .I(N__56070));
    ClkMux I__13299 (
            .O(N__56212),
            .I(N__56070));
    ClkMux I__13298 (
            .O(N__56211),
            .I(N__56070));
    ClkMux I__13297 (
            .O(N__56210),
            .I(N__56070));
    ClkMux I__13296 (
            .O(N__56209),
            .I(N__56070));
    ClkMux I__13295 (
            .O(N__56208),
            .I(N__56070));
    ClkMux I__13294 (
            .O(N__56207),
            .I(N__56070));
    ClkMux I__13293 (
            .O(N__56206),
            .I(N__56070));
    ClkMux I__13292 (
            .O(N__56205),
            .I(N__56070));
    ClkMux I__13291 (
            .O(N__56204),
            .I(N__56070));
    ClkMux I__13290 (
            .O(N__56203),
            .I(N__56070));
    ClkMux I__13289 (
            .O(N__56202),
            .I(N__56070));
    ClkMux I__13288 (
            .O(N__56201),
            .I(N__56070));
    ClkMux I__13287 (
            .O(N__56200),
            .I(N__56070));
    ClkMux I__13286 (
            .O(N__56199),
            .I(N__56070));
    GlobalMux I__13285 (
            .O(N__56070),
            .I(N__56067));
    gio2CtrlBuf I__13284 (
            .O(N__56067),
            .I(CLK_N));
    CEMux I__13283 (
            .O(N__56064),
            .I(N__56060));
    CEMux I__13282 (
            .O(N__56063),
            .I(N__56057));
    LocalMux I__13281 (
            .O(N__56060),
            .I(N__56053));
    LocalMux I__13280 (
            .O(N__56057),
            .I(N__56050));
    CEMux I__13279 (
            .O(N__56056),
            .I(N__56047));
    Span4Mux_h I__13278 (
            .O(N__56053),
            .I(N__56040));
    Span4Mux_h I__13277 (
            .O(N__56050),
            .I(N__56040));
    LocalMux I__13276 (
            .O(N__56047),
            .I(N__56040));
    Span4Mux_h I__13275 (
            .O(N__56040),
            .I(N__56037));
    Odrv4 I__13274 (
            .O(N__56037),
            .I(n5201));
    SRMux I__13273 (
            .O(N__56034),
            .I(N__56031));
    LocalMux I__13272 (
            .O(N__56031),
            .I(N__56026));
    SRMux I__13271 (
            .O(N__56030),
            .I(N__56023));
    SRMux I__13270 (
            .O(N__56029),
            .I(N__56020));
    Span4Mux_h I__13269 (
            .O(N__56026),
            .I(N__56015));
    LocalMux I__13268 (
            .O(N__56023),
            .I(N__56015));
    LocalMux I__13267 (
            .O(N__56020),
            .I(N__56012));
    Span4Mux_h I__13266 (
            .O(N__56015),
            .I(N__56009));
    Span12Mux_s3_v I__13265 (
            .O(N__56012),
            .I(N__56006));
    Odrv4 I__13264 (
            .O(N__56009),
            .I(n5253));
    Odrv12 I__13263 (
            .O(N__56006),
            .I(n5253));
    InMux I__13262 (
            .O(N__56001),
            .I(N__55998));
    LocalMux I__13261 (
            .O(N__55998),
            .I(GHA));
    InMux I__13260 (
            .O(N__55995),
            .I(N__55990));
    InMux I__13259 (
            .O(N__55994),
            .I(N__55985));
    InMux I__13258 (
            .O(N__55993),
            .I(N__55985));
    LocalMux I__13257 (
            .O(N__55990),
            .I(N__55980));
    LocalMux I__13256 (
            .O(N__55985),
            .I(N__55980));
    Span4Mux_s2_v I__13255 (
            .O(N__55980),
            .I(N__55977));
    Odrv4 I__13254 (
            .O(N__55977),
            .I(pwm_out));
    IoInMux I__13253 (
            .O(N__55974),
            .I(N__55971));
    LocalMux I__13252 (
            .O(N__55971),
            .I(N__55968));
    IoSpan4Mux I__13251 (
            .O(N__55968),
            .I(N__55965));
    Span4Mux_s0_v I__13250 (
            .O(N__55965),
            .I(N__55962));
    Odrv4 I__13249 (
            .O(N__55962),
            .I(INHA_c_0));
    InMux I__13248 (
            .O(N__55959),
            .I(N__55956));
    LocalMux I__13247 (
            .O(N__55956),
            .I(N__55952));
    InMux I__13246 (
            .O(N__55955),
            .I(N__55949));
    Span4Mux_h I__13245 (
            .O(N__55952),
            .I(N__55946));
    LocalMux I__13244 (
            .O(N__55949),
            .I(sweep_counter_15));
    Odrv4 I__13243 (
            .O(N__55946),
            .I(sweep_counter_15));
    InMux I__13242 (
            .O(N__55941),
            .I(n13067));
    InMux I__13241 (
            .O(N__55938),
            .I(N__55934));
    InMux I__13240 (
            .O(N__55937),
            .I(N__55931));
    LocalMux I__13239 (
            .O(N__55934),
            .I(N__55928));
    LocalMux I__13238 (
            .O(N__55931),
            .I(sweep_counter_16));
    Odrv4 I__13237 (
            .O(N__55928),
            .I(sweep_counter_16));
    InMux I__13236 (
            .O(N__55923),
            .I(bfn_16_27_0_));
    InMux I__13235 (
            .O(N__55920),
            .I(n13069));
    SRMux I__13234 (
            .O(N__55917),
            .I(N__55913));
    CEMux I__13233 (
            .O(N__55916),
            .I(N__55908));
    LocalMux I__13232 (
            .O(N__55913),
            .I(N__55905));
    SRMux I__13231 (
            .O(N__55912),
            .I(N__55902));
    CEMux I__13230 (
            .O(N__55911),
            .I(N__55899));
    LocalMux I__13229 (
            .O(N__55908),
            .I(N__55894));
    Span4Mux_v I__13228 (
            .O(N__55905),
            .I(N__55891));
    LocalMux I__13227 (
            .O(N__55902),
            .I(N__55888));
    LocalMux I__13226 (
            .O(N__55899),
            .I(N__55885));
    CEMux I__13225 (
            .O(N__55898),
            .I(N__55882));
    SRMux I__13224 (
            .O(N__55897),
            .I(N__55878));
    Span4Mux_h I__13223 (
            .O(N__55894),
            .I(N__55875));
    Span4Mux_v I__13222 (
            .O(N__55891),
            .I(N__55872));
    Span4Mux_h I__13221 (
            .O(N__55888),
            .I(N__55869));
    Span4Mux_v I__13220 (
            .O(N__55885),
            .I(N__55866));
    LocalMux I__13219 (
            .O(N__55882),
            .I(N__55863));
    CEMux I__13218 (
            .O(N__55881),
            .I(N__55860));
    LocalMux I__13217 (
            .O(N__55878),
            .I(N__55857));
    Span4Mux_v I__13216 (
            .O(N__55875),
            .I(N__55850));
    Span4Mux_h I__13215 (
            .O(N__55872),
            .I(N__55850));
    Span4Mux_v I__13214 (
            .O(N__55869),
            .I(N__55850));
    Span4Mux_h I__13213 (
            .O(N__55866),
            .I(N__55841));
    Span4Mux_v I__13212 (
            .O(N__55863),
            .I(N__55841));
    LocalMux I__13211 (
            .O(N__55860),
            .I(N__55841));
    Span4Mux_h I__13210 (
            .O(N__55857),
            .I(N__55841));
    Odrv4 I__13209 (
            .O(N__55850),
            .I(n5215));
    Odrv4 I__13208 (
            .O(N__55841),
            .I(n5215));
    InMux I__13207 (
            .O(N__55836),
            .I(N__55832));
    InMux I__13206 (
            .O(N__55835),
            .I(N__55829));
    LocalMux I__13205 (
            .O(N__55832),
            .I(N__55826));
    LocalMux I__13204 (
            .O(N__55829),
            .I(sweep_counter_8));
    Odrv4 I__13203 (
            .O(N__55826),
            .I(sweep_counter_8));
    InMux I__13202 (
            .O(N__55821),
            .I(N__55817));
    InMux I__13201 (
            .O(N__55820),
            .I(N__55814));
    LocalMux I__13200 (
            .O(N__55817),
            .I(N__55811));
    LocalMux I__13199 (
            .O(N__55814),
            .I(sweep_counter_14));
    Odrv4 I__13198 (
            .O(N__55811),
            .I(sweep_counter_14));
    InMux I__13197 (
            .O(N__55806),
            .I(N__55802));
    InMux I__13196 (
            .O(N__55805),
            .I(N__55799));
    LocalMux I__13195 (
            .O(N__55802),
            .I(N__55796));
    LocalMux I__13194 (
            .O(N__55799),
            .I(sweep_counter_13));
    Odrv4 I__13193 (
            .O(N__55796),
            .I(sweep_counter_13));
    InMux I__13192 (
            .O(N__55791),
            .I(N__55787));
    InMux I__13191 (
            .O(N__55790),
            .I(N__55784));
    LocalMux I__13190 (
            .O(N__55787),
            .I(sweep_counter_17));
    LocalMux I__13189 (
            .O(N__55784),
            .I(sweep_counter_17));
    CascadeMux I__13188 (
            .O(N__55779),
            .I(n6_adj_712_cascade_));
    InMux I__13187 (
            .O(N__55776),
            .I(N__55772));
    InMux I__13186 (
            .O(N__55775),
            .I(N__55769));
    LocalMux I__13185 (
            .O(N__55772),
            .I(N__55766));
    LocalMux I__13184 (
            .O(N__55769),
            .I(sweep_counter_12));
    Odrv4 I__13183 (
            .O(N__55766),
            .I(sweep_counter_12));
    InMux I__13182 (
            .O(N__55761),
            .I(N__55757));
    InMux I__13181 (
            .O(N__55760),
            .I(N__55754));
    LocalMux I__13180 (
            .O(N__55757),
            .I(N__55751));
    LocalMux I__13179 (
            .O(N__55754),
            .I(N__55748));
    Span4Mux_h I__13178 (
            .O(N__55751),
            .I(N__55745));
    Span4Mux_h I__13177 (
            .O(N__55748),
            .I(N__55742));
    Span4Mux_v I__13176 (
            .O(N__55745),
            .I(N__55739));
    Odrv4 I__13175 (
            .O(N__55742),
            .I(n13968));
    Odrv4 I__13174 (
            .O(N__55739),
            .I(n13968));
    InMux I__13173 (
            .O(N__55734),
            .I(N__55731));
    LocalMux I__13172 (
            .O(N__55731),
            .I(GHC));
    IoInMux I__13171 (
            .O(N__55728),
            .I(N__55725));
    LocalMux I__13170 (
            .O(N__55725),
            .I(N__55722));
    Span12Mux_s0_v I__13169 (
            .O(N__55722),
            .I(N__55719));
    Odrv12 I__13168 (
            .O(N__55719),
            .I(INHC_c_0));
    InMux I__13167 (
            .O(N__55716),
            .I(N__55712));
    InMux I__13166 (
            .O(N__55715),
            .I(N__55709));
    LocalMux I__13165 (
            .O(N__55712),
            .I(N__55706));
    LocalMux I__13164 (
            .O(N__55709),
            .I(sweep_counter_6));
    Odrv4 I__13163 (
            .O(N__55706),
            .I(sweep_counter_6));
    InMux I__13162 (
            .O(N__55701),
            .I(n13058));
    InMux I__13161 (
            .O(N__55698),
            .I(N__55695));
    LocalMux I__13160 (
            .O(N__55695),
            .I(N__55691));
    InMux I__13159 (
            .O(N__55694),
            .I(N__55688));
    Span4Mux_h I__13158 (
            .O(N__55691),
            .I(N__55685));
    LocalMux I__13157 (
            .O(N__55688),
            .I(sweep_counter_7));
    Odrv4 I__13156 (
            .O(N__55685),
            .I(sweep_counter_7));
    InMux I__13155 (
            .O(N__55680),
            .I(n13059));
    InMux I__13154 (
            .O(N__55677),
            .I(bfn_16_26_0_));
    CascadeMux I__13153 (
            .O(N__55674),
            .I(N__55671));
    InMux I__13152 (
            .O(N__55671),
            .I(N__55668));
    LocalMux I__13151 (
            .O(N__55668),
            .I(N__55664));
    InMux I__13150 (
            .O(N__55667),
            .I(N__55661));
    Span4Mux_h I__13149 (
            .O(N__55664),
            .I(N__55658));
    LocalMux I__13148 (
            .O(N__55661),
            .I(sweep_counter_9));
    Odrv4 I__13147 (
            .O(N__55658),
            .I(sweep_counter_9));
    InMux I__13146 (
            .O(N__55653),
            .I(n13061));
    InMux I__13145 (
            .O(N__55650),
            .I(N__55647));
    LocalMux I__13144 (
            .O(N__55647),
            .I(N__55643));
    InMux I__13143 (
            .O(N__55646),
            .I(N__55640));
    Span4Mux_h I__13142 (
            .O(N__55643),
            .I(N__55637));
    LocalMux I__13141 (
            .O(N__55640),
            .I(sweep_counter_10));
    Odrv4 I__13140 (
            .O(N__55637),
            .I(sweep_counter_10));
    InMux I__13139 (
            .O(N__55632),
            .I(n13062));
    InMux I__13138 (
            .O(N__55629),
            .I(N__55626));
    LocalMux I__13137 (
            .O(N__55626),
            .I(N__55622));
    InMux I__13136 (
            .O(N__55625),
            .I(N__55619));
    Span4Mux_h I__13135 (
            .O(N__55622),
            .I(N__55616));
    LocalMux I__13134 (
            .O(N__55619),
            .I(sweep_counter_11));
    Odrv4 I__13133 (
            .O(N__55616),
            .I(sweep_counter_11));
    InMux I__13132 (
            .O(N__55611),
            .I(n13063));
    InMux I__13131 (
            .O(N__55608),
            .I(n13064));
    InMux I__13130 (
            .O(N__55605),
            .I(n13065));
    InMux I__13129 (
            .O(N__55602),
            .I(n13066));
    CascadeMux I__13128 (
            .O(N__55599),
            .I(N__55596));
    InMux I__13127 (
            .O(N__55596),
            .I(N__55593));
    LocalMux I__13126 (
            .O(N__55593),
            .I(N__55588));
    InMux I__13125 (
            .O(N__55592),
            .I(N__55583));
    InMux I__13124 (
            .O(N__55591),
            .I(N__55583));
    Span4Mux_v I__13123 (
            .O(N__55588),
            .I(N__55580));
    LocalMux I__13122 (
            .O(N__55583),
            .I(n1027));
    Odrv4 I__13121 (
            .O(N__55580),
            .I(n1027));
    InMux I__13120 (
            .O(N__55575),
            .I(N__55572));
    LocalMux I__13119 (
            .O(N__55572),
            .I(N__55569));
    Odrv4 I__13118 (
            .O(N__55569),
            .I(n1094));
    InMux I__13117 (
            .O(N__55566),
            .I(n12520));
    CascadeMux I__13116 (
            .O(N__55563),
            .I(N__55559));
    InMux I__13115 (
            .O(N__55562),
            .I(N__55521));
    InMux I__13114 (
            .O(N__55559),
            .I(N__55521));
    CascadeMux I__13113 (
            .O(N__55558),
            .I(N__55518));
    CascadeMux I__13112 (
            .O(N__55557),
            .I(N__55515));
    CascadeMux I__13111 (
            .O(N__55556),
            .I(N__55512));
    CascadeMux I__13110 (
            .O(N__55555),
            .I(N__55509));
    CascadeMux I__13109 (
            .O(N__55554),
            .I(N__55506));
    CascadeMux I__13108 (
            .O(N__55553),
            .I(N__55503));
    CascadeMux I__13107 (
            .O(N__55552),
            .I(N__55500));
    CascadeMux I__13106 (
            .O(N__55551),
            .I(N__55497));
    CascadeMux I__13105 (
            .O(N__55550),
            .I(N__55487));
    CascadeMux I__13104 (
            .O(N__55549),
            .I(N__55482));
    CascadeMux I__13103 (
            .O(N__55548),
            .I(N__55479));
    CascadeMux I__13102 (
            .O(N__55547),
            .I(N__55473));
    InMux I__13101 (
            .O(N__55546),
            .I(N__55470));
    InMux I__13100 (
            .O(N__55545),
            .I(N__55463));
    InMux I__13099 (
            .O(N__55544),
            .I(N__55463));
    InMux I__13098 (
            .O(N__55543),
            .I(N__55463));
    InMux I__13097 (
            .O(N__55542),
            .I(N__55456));
    InMux I__13096 (
            .O(N__55541),
            .I(N__55456));
    InMux I__13095 (
            .O(N__55540),
            .I(N__55456));
    CascadeMux I__13094 (
            .O(N__55539),
            .I(N__55450));
    CascadeMux I__13093 (
            .O(N__55538),
            .I(N__55447));
    CascadeMux I__13092 (
            .O(N__55537),
            .I(N__55441));
    CascadeMux I__13091 (
            .O(N__55536),
            .I(N__55438));
    CascadeMux I__13090 (
            .O(N__55535),
            .I(N__55428));
    CascadeMux I__13089 (
            .O(N__55534),
            .I(N__55422));
    CascadeMux I__13088 (
            .O(N__55533),
            .I(N__55415));
    CascadeMux I__13087 (
            .O(N__55532),
            .I(N__55412));
    CascadeMux I__13086 (
            .O(N__55531),
            .I(N__55409));
    CascadeMux I__13085 (
            .O(N__55530),
            .I(N__55406));
    CascadeMux I__13084 (
            .O(N__55529),
            .I(N__55403));
    CascadeMux I__13083 (
            .O(N__55528),
            .I(N__55400));
    CascadeMux I__13082 (
            .O(N__55527),
            .I(N__55397));
    CascadeMux I__13081 (
            .O(N__55526),
            .I(N__55394));
    LocalMux I__13080 (
            .O(N__55521),
            .I(N__55389));
    InMux I__13079 (
            .O(N__55518),
            .I(N__55380));
    InMux I__13078 (
            .O(N__55515),
            .I(N__55380));
    InMux I__13077 (
            .O(N__55512),
            .I(N__55380));
    InMux I__13076 (
            .O(N__55509),
            .I(N__55380));
    InMux I__13075 (
            .O(N__55506),
            .I(N__55371));
    InMux I__13074 (
            .O(N__55503),
            .I(N__55371));
    InMux I__13073 (
            .O(N__55500),
            .I(N__55371));
    InMux I__13072 (
            .O(N__55497),
            .I(N__55371));
    InMux I__13071 (
            .O(N__55496),
            .I(N__55368));
    InMux I__13070 (
            .O(N__55495),
            .I(N__55361));
    InMux I__13069 (
            .O(N__55494),
            .I(N__55361));
    InMux I__13068 (
            .O(N__55493),
            .I(N__55361));
    CascadeMux I__13067 (
            .O(N__55492),
            .I(N__55358));
    CascadeMux I__13066 (
            .O(N__55491),
            .I(N__55352));
    CascadeMux I__13065 (
            .O(N__55490),
            .I(N__55341));
    InMux I__13064 (
            .O(N__55487),
            .I(N__55333));
    InMux I__13063 (
            .O(N__55486),
            .I(N__55333));
    InMux I__13062 (
            .O(N__55485),
            .I(N__55333));
    InMux I__13061 (
            .O(N__55482),
            .I(N__55322));
    InMux I__13060 (
            .O(N__55479),
            .I(N__55322));
    InMux I__13059 (
            .O(N__55478),
            .I(N__55322));
    InMux I__13058 (
            .O(N__55477),
            .I(N__55322));
    InMux I__13057 (
            .O(N__55476),
            .I(N__55322));
    InMux I__13056 (
            .O(N__55473),
            .I(N__55319));
    LocalMux I__13055 (
            .O(N__55470),
            .I(N__55312));
    LocalMux I__13054 (
            .O(N__55463),
            .I(N__55312));
    LocalMux I__13053 (
            .O(N__55456),
            .I(N__55312));
    InMux I__13052 (
            .O(N__55455),
            .I(N__55305));
    InMux I__13051 (
            .O(N__55454),
            .I(N__55305));
    InMux I__13050 (
            .O(N__55453),
            .I(N__55305));
    InMux I__13049 (
            .O(N__55450),
            .I(N__55294));
    InMux I__13048 (
            .O(N__55447),
            .I(N__55294));
    InMux I__13047 (
            .O(N__55446),
            .I(N__55294));
    InMux I__13046 (
            .O(N__55445),
            .I(N__55294));
    InMux I__13045 (
            .O(N__55444),
            .I(N__55294));
    InMux I__13044 (
            .O(N__55441),
            .I(N__55289));
    InMux I__13043 (
            .O(N__55438),
            .I(N__55289));
    InMux I__13042 (
            .O(N__55437),
            .I(N__55270));
    InMux I__13041 (
            .O(N__55436),
            .I(N__55270));
    InMux I__13040 (
            .O(N__55435),
            .I(N__55263));
    InMux I__13039 (
            .O(N__55434),
            .I(N__55263));
    InMux I__13038 (
            .O(N__55433),
            .I(N__55263));
    InMux I__13037 (
            .O(N__55432),
            .I(N__55252));
    InMux I__13036 (
            .O(N__55431),
            .I(N__55252));
    InMux I__13035 (
            .O(N__55428),
            .I(N__55252));
    InMux I__13034 (
            .O(N__55427),
            .I(N__55252));
    InMux I__13033 (
            .O(N__55426),
            .I(N__55252));
    InMux I__13032 (
            .O(N__55425),
            .I(N__55241));
    InMux I__13031 (
            .O(N__55422),
            .I(N__55241));
    InMux I__13030 (
            .O(N__55421),
            .I(N__55241));
    InMux I__13029 (
            .O(N__55420),
            .I(N__55241));
    InMux I__13028 (
            .O(N__55419),
            .I(N__55241));
    InMux I__13027 (
            .O(N__55418),
            .I(N__55237));
    InMux I__13026 (
            .O(N__55415),
            .I(N__55228));
    InMux I__13025 (
            .O(N__55412),
            .I(N__55228));
    InMux I__13024 (
            .O(N__55409),
            .I(N__55228));
    InMux I__13023 (
            .O(N__55406),
            .I(N__55228));
    InMux I__13022 (
            .O(N__55403),
            .I(N__55219));
    InMux I__13021 (
            .O(N__55400),
            .I(N__55219));
    InMux I__13020 (
            .O(N__55397),
            .I(N__55219));
    InMux I__13019 (
            .O(N__55394),
            .I(N__55219));
    CascadeMux I__13018 (
            .O(N__55393),
            .I(N__55215));
    CascadeMux I__13017 (
            .O(N__55392),
            .I(N__55206));
    Span4Mux_v I__13016 (
            .O(N__55389),
            .I(N__55192));
    LocalMux I__13015 (
            .O(N__55380),
            .I(N__55192));
    LocalMux I__13014 (
            .O(N__55371),
            .I(N__55192));
    LocalMux I__13013 (
            .O(N__55368),
            .I(N__55192));
    LocalMux I__13012 (
            .O(N__55361),
            .I(N__55192));
    InMux I__13011 (
            .O(N__55358),
            .I(N__55183));
    InMux I__13010 (
            .O(N__55357),
            .I(N__55183));
    InMux I__13009 (
            .O(N__55356),
            .I(N__55183));
    InMux I__13008 (
            .O(N__55355),
            .I(N__55183));
    InMux I__13007 (
            .O(N__55352),
            .I(N__55174));
    InMux I__13006 (
            .O(N__55351),
            .I(N__55174));
    InMux I__13005 (
            .O(N__55350),
            .I(N__55174));
    InMux I__13004 (
            .O(N__55349),
            .I(N__55174));
    InMux I__13003 (
            .O(N__55348),
            .I(N__55167));
    InMux I__13002 (
            .O(N__55347),
            .I(N__55167));
    InMux I__13001 (
            .O(N__55346),
            .I(N__55167));
    CascadeMux I__13000 (
            .O(N__55345),
            .I(N__55161));
    InMux I__12999 (
            .O(N__55344),
            .I(N__55152));
    InMux I__12998 (
            .O(N__55341),
            .I(N__55152));
    CascadeMux I__12997 (
            .O(N__55340),
            .I(N__55148));
    LocalMux I__12996 (
            .O(N__55333),
            .I(N__55141));
    LocalMux I__12995 (
            .O(N__55322),
            .I(N__55141));
    LocalMux I__12994 (
            .O(N__55319),
            .I(N__55141));
    Span4Mux_v I__12993 (
            .O(N__55312),
            .I(N__55132));
    LocalMux I__12992 (
            .O(N__55305),
            .I(N__55132));
    LocalMux I__12991 (
            .O(N__55294),
            .I(N__55132));
    LocalMux I__12990 (
            .O(N__55289),
            .I(N__55132));
    CascadeMux I__12989 (
            .O(N__55288),
            .I(N__55122));
    InMux I__12988 (
            .O(N__55287),
            .I(N__55110));
    InMux I__12987 (
            .O(N__55286),
            .I(N__55110));
    InMux I__12986 (
            .O(N__55285),
            .I(N__55110));
    InMux I__12985 (
            .O(N__55284),
            .I(N__55101));
    InMux I__12984 (
            .O(N__55283),
            .I(N__55101));
    InMux I__12983 (
            .O(N__55282),
            .I(N__55101));
    InMux I__12982 (
            .O(N__55281),
            .I(N__55101));
    InMux I__12981 (
            .O(N__55280),
            .I(N__55098));
    CascadeMux I__12980 (
            .O(N__55279),
            .I(N__55093));
    CascadeMux I__12979 (
            .O(N__55278),
            .I(N__55088));
    CascadeMux I__12978 (
            .O(N__55277),
            .I(N__55073));
    CascadeMux I__12977 (
            .O(N__55276),
            .I(N__55070));
    CascadeMux I__12976 (
            .O(N__55275),
            .I(N__55067));
    LocalMux I__12975 (
            .O(N__55270),
            .I(N__55046));
    LocalMux I__12974 (
            .O(N__55263),
            .I(N__55046));
    LocalMux I__12973 (
            .O(N__55252),
            .I(N__55046));
    LocalMux I__12972 (
            .O(N__55241),
            .I(N__55046));
    CascadeMux I__12971 (
            .O(N__55240),
            .I(N__55042));
    LocalMux I__12970 (
            .O(N__55237),
            .I(N__55023));
    LocalMux I__12969 (
            .O(N__55228),
            .I(N__55023));
    LocalMux I__12968 (
            .O(N__55219),
            .I(N__55023));
    InMux I__12967 (
            .O(N__55218),
            .I(N__55020));
    InMux I__12966 (
            .O(N__55215),
            .I(N__55011));
    InMux I__12965 (
            .O(N__55214),
            .I(N__55011));
    InMux I__12964 (
            .O(N__55213),
            .I(N__55011));
    InMux I__12963 (
            .O(N__55212),
            .I(N__55011));
    InMux I__12962 (
            .O(N__55211),
            .I(N__55004));
    InMux I__12961 (
            .O(N__55210),
            .I(N__55004));
    InMux I__12960 (
            .O(N__55209),
            .I(N__55004));
    InMux I__12959 (
            .O(N__55206),
            .I(N__54995));
    InMux I__12958 (
            .O(N__55205),
            .I(N__54995));
    InMux I__12957 (
            .O(N__55204),
            .I(N__54995));
    InMux I__12956 (
            .O(N__55203),
            .I(N__54995));
    Span4Mux_v I__12955 (
            .O(N__55192),
            .I(N__54988));
    LocalMux I__12954 (
            .O(N__55183),
            .I(N__54988));
    LocalMux I__12953 (
            .O(N__55174),
            .I(N__54988));
    LocalMux I__12952 (
            .O(N__55167),
            .I(N__54985));
    InMux I__12951 (
            .O(N__55166),
            .I(N__54974));
    InMux I__12950 (
            .O(N__55165),
            .I(N__54974));
    InMux I__12949 (
            .O(N__55164),
            .I(N__54974));
    InMux I__12948 (
            .O(N__55161),
            .I(N__54974));
    InMux I__12947 (
            .O(N__55160),
            .I(N__54974));
    InMux I__12946 (
            .O(N__55159),
            .I(N__54967));
    InMux I__12945 (
            .O(N__55158),
            .I(N__54967));
    InMux I__12944 (
            .O(N__55157),
            .I(N__54967));
    LocalMux I__12943 (
            .O(N__55152),
            .I(N__54964));
    InMux I__12942 (
            .O(N__55151),
            .I(N__54959));
    InMux I__12941 (
            .O(N__55148),
            .I(N__54959));
    Span4Mux_s3_h I__12940 (
            .O(N__55141),
            .I(N__54947));
    Span4Mux_v I__12939 (
            .O(N__55132),
            .I(N__54947));
    InMux I__12938 (
            .O(N__55131),
            .I(N__54944));
    InMux I__12937 (
            .O(N__55130),
            .I(N__54937));
    InMux I__12936 (
            .O(N__55129),
            .I(N__54937));
    InMux I__12935 (
            .O(N__55128),
            .I(N__54937));
    InMux I__12934 (
            .O(N__55127),
            .I(N__54932));
    InMux I__12933 (
            .O(N__55126),
            .I(N__54932));
    InMux I__12932 (
            .O(N__55125),
            .I(N__54925));
    InMux I__12931 (
            .O(N__55122),
            .I(N__54925));
    InMux I__12930 (
            .O(N__55121),
            .I(N__54925));
    InMux I__12929 (
            .O(N__55120),
            .I(N__54922));
    InMux I__12928 (
            .O(N__55119),
            .I(N__54915));
    InMux I__12927 (
            .O(N__55118),
            .I(N__54915));
    InMux I__12926 (
            .O(N__55117),
            .I(N__54915));
    LocalMux I__12925 (
            .O(N__55110),
            .I(N__54908));
    LocalMux I__12924 (
            .O(N__55101),
            .I(N__54908));
    LocalMux I__12923 (
            .O(N__55098),
            .I(N__54908));
    InMux I__12922 (
            .O(N__55097),
            .I(N__54903));
    InMux I__12921 (
            .O(N__55096),
            .I(N__54903));
    InMux I__12920 (
            .O(N__55093),
            .I(N__54894));
    InMux I__12919 (
            .O(N__55092),
            .I(N__54894));
    InMux I__12918 (
            .O(N__55091),
            .I(N__54894));
    InMux I__12917 (
            .O(N__55088),
            .I(N__54894));
    InMux I__12916 (
            .O(N__55087),
            .I(N__54887));
    InMux I__12915 (
            .O(N__55086),
            .I(N__54884));
    CascadeMux I__12914 (
            .O(N__55085),
            .I(N__54857));
    CascadeMux I__12913 (
            .O(N__55084),
            .I(N__54854));
    CascadeMux I__12912 (
            .O(N__55083),
            .I(N__54851));
    CascadeMux I__12911 (
            .O(N__55082),
            .I(N__54848));
    CascadeMux I__12910 (
            .O(N__55081),
            .I(N__54845));
    CascadeMux I__12909 (
            .O(N__55080),
            .I(N__54842));
    CascadeMux I__12908 (
            .O(N__55079),
            .I(N__54839));
    CascadeMux I__12907 (
            .O(N__55078),
            .I(N__54836));
    CascadeMux I__12906 (
            .O(N__55077),
            .I(N__54833));
    CascadeMux I__12905 (
            .O(N__55076),
            .I(N__54830));
    InMux I__12904 (
            .O(N__55073),
            .I(N__54823));
    InMux I__12903 (
            .O(N__55070),
            .I(N__54823));
    InMux I__12902 (
            .O(N__55067),
            .I(N__54823));
    CascadeMux I__12901 (
            .O(N__55066),
            .I(N__54820));
    CascadeMux I__12900 (
            .O(N__55065),
            .I(N__54817));
    CascadeMux I__12899 (
            .O(N__55064),
            .I(N__54814));
    CascadeMux I__12898 (
            .O(N__55063),
            .I(N__54810));
    CascadeMux I__12897 (
            .O(N__55062),
            .I(N__54807));
    CascadeMux I__12896 (
            .O(N__55061),
            .I(N__54804));
    CascadeMux I__12895 (
            .O(N__55060),
            .I(N__54801));
    CascadeMux I__12894 (
            .O(N__55059),
            .I(N__54798));
    CascadeMux I__12893 (
            .O(N__55058),
            .I(N__54795));
    CascadeMux I__12892 (
            .O(N__55057),
            .I(N__54789));
    CascadeMux I__12891 (
            .O(N__55056),
            .I(N__54780));
    CascadeMux I__12890 (
            .O(N__55055),
            .I(N__54777));
    Span4Mux_v I__12889 (
            .O(N__55046),
            .I(N__54773));
    InMux I__12888 (
            .O(N__55045),
            .I(N__54770));
    InMux I__12887 (
            .O(N__55042),
            .I(N__54767));
    CascadeMux I__12886 (
            .O(N__55041),
            .I(N__54764));
    CascadeMux I__12885 (
            .O(N__55040),
            .I(N__54759));
    CascadeMux I__12884 (
            .O(N__55039),
            .I(N__54753));
    CascadeMux I__12883 (
            .O(N__55038),
            .I(N__54750));
    CascadeMux I__12882 (
            .O(N__55037),
            .I(N__54747));
    CascadeMux I__12881 (
            .O(N__55036),
            .I(N__54740));
    CascadeMux I__12880 (
            .O(N__55035),
            .I(N__54737));
    CascadeMux I__12879 (
            .O(N__55034),
            .I(N__54733));
    InMux I__12878 (
            .O(N__55033),
            .I(N__54714));
    InMux I__12877 (
            .O(N__55032),
            .I(N__54714));
    InMux I__12876 (
            .O(N__55031),
            .I(N__54714));
    CascadeMux I__12875 (
            .O(N__55030),
            .I(N__54710));
    Span4Mux_v I__12874 (
            .O(N__55023),
            .I(N__54702));
    LocalMux I__12873 (
            .O(N__55020),
            .I(N__54695));
    LocalMux I__12872 (
            .O(N__55011),
            .I(N__54695));
    LocalMux I__12871 (
            .O(N__55004),
            .I(N__54690));
    LocalMux I__12870 (
            .O(N__54995),
            .I(N__54690));
    Span4Mux_h I__12869 (
            .O(N__54988),
            .I(N__54677));
    Span4Mux_v I__12868 (
            .O(N__54985),
            .I(N__54677));
    LocalMux I__12867 (
            .O(N__54974),
            .I(N__54677));
    LocalMux I__12866 (
            .O(N__54967),
            .I(N__54677));
    Span4Mux_v I__12865 (
            .O(N__54964),
            .I(N__54677));
    LocalMux I__12864 (
            .O(N__54959),
            .I(N__54677));
    InMux I__12863 (
            .O(N__54958),
            .I(N__54668));
    InMux I__12862 (
            .O(N__54957),
            .I(N__54668));
    InMux I__12861 (
            .O(N__54956),
            .I(N__54668));
    InMux I__12860 (
            .O(N__54955),
            .I(N__54668));
    InMux I__12859 (
            .O(N__54954),
            .I(N__54663));
    InMux I__12858 (
            .O(N__54953),
            .I(N__54663));
    CascadeMux I__12857 (
            .O(N__54952),
            .I(N__54658));
    Span4Mux_h I__12856 (
            .O(N__54947),
            .I(N__54640));
    LocalMux I__12855 (
            .O(N__54944),
            .I(N__54627));
    LocalMux I__12854 (
            .O(N__54937),
            .I(N__54627));
    LocalMux I__12853 (
            .O(N__54932),
            .I(N__54627));
    LocalMux I__12852 (
            .O(N__54925),
            .I(N__54627));
    LocalMux I__12851 (
            .O(N__54922),
            .I(N__54627));
    LocalMux I__12850 (
            .O(N__54915),
            .I(N__54627));
    Span4Mux_v I__12849 (
            .O(N__54908),
            .I(N__54624));
    LocalMux I__12848 (
            .O(N__54903),
            .I(N__54621));
    LocalMux I__12847 (
            .O(N__54894),
            .I(N__54618));
    InMux I__12846 (
            .O(N__54893),
            .I(N__54615));
    InMux I__12845 (
            .O(N__54892),
            .I(N__54608));
    InMux I__12844 (
            .O(N__54891),
            .I(N__54608));
    InMux I__12843 (
            .O(N__54890),
            .I(N__54608));
    LocalMux I__12842 (
            .O(N__54887),
            .I(N__54603));
    LocalMux I__12841 (
            .O(N__54884),
            .I(N__54603));
    InMux I__12840 (
            .O(N__54883),
            .I(N__54596));
    InMux I__12839 (
            .O(N__54882),
            .I(N__54596));
    InMux I__12838 (
            .O(N__54881),
            .I(N__54596));
    CascadeMux I__12837 (
            .O(N__54880),
            .I(N__54593));
    CascadeMux I__12836 (
            .O(N__54879),
            .I(N__54583));
    CascadeMux I__12835 (
            .O(N__54878),
            .I(N__54569));
    CascadeMux I__12834 (
            .O(N__54877),
            .I(N__54566));
    CascadeMux I__12833 (
            .O(N__54876),
            .I(N__54561));
    CascadeMux I__12832 (
            .O(N__54875),
            .I(N__54558));
    CascadeMux I__12831 (
            .O(N__54874),
            .I(N__54553));
    CascadeMux I__12830 (
            .O(N__54873),
            .I(N__54550));
    CascadeMux I__12829 (
            .O(N__54872),
            .I(N__54547));
    CascadeMux I__12828 (
            .O(N__54871),
            .I(N__54544));
    CascadeMux I__12827 (
            .O(N__54870),
            .I(N__54541));
    CascadeMux I__12826 (
            .O(N__54869),
            .I(N__54538));
    CascadeMux I__12825 (
            .O(N__54868),
            .I(N__54535));
    CascadeMux I__12824 (
            .O(N__54867),
            .I(N__54531));
    CascadeMux I__12823 (
            .O(N__54866),
            .I(N__54528));
    CascadeMux I__12822 (
            .O(N__54865),
            .I(N__54525));
    CascadeMux I__12821 (
            .O(N__54864),
            .I(N__54522));
    CascadeMux I__12820 (
            .O(N__54863),
            .I(N__54519));
    CascadeMux I__12819 (
            .O(N__54862),
            .I(N__54516));
    CascadeMux I__12818 (
            .O(N__54861),
            .I(N__54512));
    CascadeMux I__12817 (
            .O(N__54860),
            .I(N__54509));
    InMux I__12816 (
            .O(N__54857),
            .I(N__54499));
    InMux I__12815 (
            .O(N__54854),
            .I(N__54499));
    InMux I__12814 (
            .O(N__54851),
            .I(N__54499));
    InMux I__12813 (
            .O(N__54848),
            .I(N__54492));
    InMux I__12812 (
            .O(N__54845),
            .I(N__54492));
    InMux I__12811 (
            .O(N__54842),
            .I(N__54492));
    InMux I__12810 (
            .O(N__54839),
            .I(N__54483));
    InMux I__12809 (
            .O(N__54836),
            .I(N__54483));
    InMux I__12808 (
            .O(N__54833),
            .I(N__54483));
    InMux I__12807 (
            .O(N__54830),
            .I(N__54483));
    LocalMux I__12806 (
            .O(N__54823),
            .I(N__54480));
    InMux I__12805 (
            .O(N__54820),
            .I(N__54477));
    InMux I__12804 (
            .O(N__54817),
            .I(N__54466));
    InMux I__12803 (
            .O(N__54814),
            .I(N__54466));
    InMux I__12802 (
            .O(N__54813),
            .I(N__54466));
    InMux I__12801 (
            .O(N__54810),
            .I(N__54466));
    InMux I__12800 (
            .O(N__54807),
            .I(N__54466));
    InMux I__12799 (
            .O(N__54804),
            .I(N__54457));
    InMux I__12798 (
            .O(N__54801),
            .I(N__54457));
    InMux I__12797 (
            .O(N__54798),
            .I(N__54457));
    InMux I__12796 (
            .O(N__54795),
            .I(N__54457));
    InMux I__12795 (
            .O(N__54794),
            .I(N__54452));
    InMux I__12794 (
            .O(N__54793),
            .I(N__54452));
    InMux I__12793 (
            .O(N__54792),
            .I(N__54447));
    InMux I__12792 (
            .O(N__54789),
            .I(N__54447));
    InMux I__12791 (
            .O(N__54788),
            .I(N__54438));
    InMux I__12790 (
            .O(N__54787),
            .I(N__54438));
    InMux I__12789 (
            .O(N__54786),
            .I(N__54431));
    InMux I__12788 (
            .O(N__54785),
            .I(N__54431));
    InMux I__12787 (
            .O(N__54784),
            .I(N__54431));
    InMux I__12786 (
            .O(N__54783),
            .I(N__54424));
    InMux I__12785 (
            .O(N__54780),
            .I(N__54424));
    InMux I__12784 (
            .O(N__54777),
            .I(N__54424));
    CascadeMux I__12783 (
            .O(N__54776),
            .I(N__54418));
    Span4Mux_h I__12782 (
            .O(N__54773),
            .I(N__54407));
    LocalMux I__12781 (
            .O(N__54770),
            .I(N__54407));
    LocalMux I__12780 (
            .O(N__54767),
            .I(N__54407));
    InMux I__12779 (
            .O(N__54764),
            .I(N__54402));
    InMux I__12778 (
            .O(N__54763),
            .I(N__54402));
    InMux I__12777 (
            .O(N__54762),
            .I(N__54391));
    InMux I__12776 (
            .O(N__54759),
            .I(N__54391));
    InMux I__12775 (
            .O(N__54758),
            .I(N__54391));
    InMux I__12774 (
            .O(N__54757),
            .I(N__54391));
    InMux I__12773 (
            .O(N__54756),
            .I(N__54391));
    InMux I__12772 (
            .O(N__54753),
            .I(N__54382));
    InMux I__12771 (
            .O(N__54750),
            .I(N__54382));
    InMux I__12770 (
            .O(N__54747),
            .I(N__54382));
    InMux I__12769 (
            .O(N__54746),
            .I(N__54382));
    CascadeMux I__12768 (
            .O(N__54745),
            .I(N__54376));
    CascadeMux I__12767 (
            .O(N__54744),
            .I(N__54370));
    InMux I__12766 (
            .O(N__54743),
            .I(N__54364));
    InMux I__12765 (
            .O(N__54740),
            .I(N__54357));
    InMux I__12764 (
            .O(N__54737),
            .I(N__54357));
    InMux I__12763 (
            .O(N__54736),
            .I(N__54357));
    InMux I__12762 (
            .O(N__54733),
            .I(N__54352));
    InMux I__12761 (
            .O(N__54732),
            .I(N__54352));
    CascadeMux I__12760 (
            .O(N__54731),
            .I(N__54348));
    CascadeMux I__12759 (
            .O(N__54730),
            .I(N__54342));
    CascadeMux I__12758 (
            .O(N__54729),
            .I(N__54339));
    CascadeMux I__12757 (
            .O(N__54728),
            .I(N__54336));
    CascadeMux I__12756 (
            .O(N__54727),
            .I(N__54333));
    CascadeMux I__12755 (
            .O(N__54726),
            .I(N__54330));
    CascadeMux I__12754 (
            .O(N__54725),
            .I(N__54321));
    CascadeMux I__12753 (
            .O(N__54724),
            .I(N__54318));
    CascadeMux I__12752 (
            .O(N__54723),
            .I(N__54315));
    CascadeMux I__12751 (
            .O(N__54722),
            .I(N__54312));
    CascadeMux I__12750 (
            .O(N__54721),
            .I(N__54309));
    LocalMux I__12749 (
            .O(N__54714),
            .I(N__54306));
    InMux I__12748 (
            .O(N__54713),
            .I(N__54297));
    InMux I__12747 (
            .O(N__54710),
            .I(N__54297));
    InMux I__12746 (
            .O(N__54709),
            .I(N__54297));
    InMux I__12745 (
            .O(N__54708),
            .I(N__54297));
    CascadeMux I__12744 (
            .O(N__54707),
            .I(N__54294));
    CascadeMux I__12743 (
            .O(N__54706),
            .I(N__54289));
    CascadeMux I__12742 (
            .O(N__54705),
            .I(N__54284));
    Span4Mux_h I__12741 (
            .O(N__54702),
            .I(N__54280));
    InMux I__12740 (
            .O(N__54701),
            .I(N__54275));
    InMux I__12739 (
            .O(N__54700),
            .I(N__54275));
    Span4Mux_v I__12738 (
            .O(N__54695),
            .I(N__54270));
    Span4Mux_v I__12737 (
            .O(N__54690),
            .I(N__54270));
    Span4Mux_h I__12736 (
            .O(N__54677),
            .I(N__54263));
    LocalMux I__12735 (
            .O(N__54668),
            .I(N__54263));
    LocalMux I__12734 (
            .O(N__54663),
            .I(N__54263));
    InMux I__12733 (
            .O(N__54662),
            .I(N__54258));
    InMux I__12732 (
            .O(N__54661),
            .I(N__54258));
    InMux I__12731 (
            .O(N__54658),
            .I(N__54253));
    InMux I__12730 (
            .O(N__54657),
            .I(N__54253));
    CascadeMux I__12729 (
            .O(N__54656),
            .I(N__54249));
    CascadeMux I__12728 (
            .O(N__54655),
            .I(N__54237));
    CascadeMux I__12727 (
            .O(N__54654),
            .I(N__54233));
    InMux I__12726 (
            .O(N__54653),
            .I(N__54230));
    InMux I__12725 (
            .O(N__54652),
            .I(N__54223));
    InMux I__12724 (
            .O(N__54651),
            .I(N__54223));
    InMux I__12723 (
            .O(N__54650),
            .I(N__54223));
    InMux I__12722 (
            .O(N__54649),
            .I(N__54218));
    InMux I__12721 (
            .O(N__54648),
            .I(N__54218));
    InMux I__12720 (
            .O(N__54647),
            .I(N__54215));
    InMux I__12719 (
            .O(N__54646),
            .I(N__54212));
    InMux I__12718 (
            .O(N__54645),
            .I(N__54205));
    InMux I__12717 (
            .O(N__54644),
            .I(N__54205));
    InMux I__12716 (
            .O(N__54643),
            .I(N__54205));
    Span4Mux_h I__12715 (
            .O(N__54640),
            .I(N__54186));
    Span4Mux_v I__12714 (
            .O(N__54627),
            .I(N__54186));
    Span4Mux_v I__12713 (
            .O(N__54624),
            .I(N__54186));
    Span4Mux_h I__12712 (
            .O(N__54621),
            .I(N__54186));
    Span4Mux_h I__12711 (
            .O(N__54618),
            .I(N__54186));
    LocalMux I__12710 (
            .O(N__54615),
            .I(N__54186));
    LocalMux I__12709 (
            .O(N__54608),
            .I(N__54186));
    Span4Mux_v I__12708 (
            .O(N__54603),
            .I(N__54186));
    LocalMux I__12707 (
            .O(N__54596),
            .I(N__54186));
    InMux I__12706 (
            .O(N__54593),
            .I(N__54177));
    InMux I__12705 (
            .O(N__54592),
            .I(N__54177));
    InMux I__12704 (
            .O(N__54591),
            .I(N__54177));
    InMux I__12703 (
            .O(N__54590),
            .I(N__54177));
    InMux I__12702 (
            .O(N__54589),
            .I(N__54168));
    InMux I__12701 (
            .O(N__54588),
            .I(N__54168));
    InMux I__12700 (
            .O(N__54587),
            .I(N__54168));
    InMux I__12699 (
            .O(N__54586),
            .I(N__54168));
    InMux I__12698 (
            .O(N__54583),
            .I(N__54163));
    InMux I__12697 (
            .O(N__54582),
            .I(N__54163));
    InMux I__12696 (
            .O(N__54581),
            .I(N__54154));
    InMux I__12695 (
            .O(N__54580),
            .I(N__54154));
    InMux I__12694 (
            .O(N__54579),
            .I(N__54154));
    InMux I__12693 (
            .O(N__54578),
            .I(N__54154));
    InMux I__12692 (
            .O(N__54577),
            .I(N__54145));
    InMux I__12691 (
            .O(N__54576),
            .I(N__54145));
    InMux I__12690 (
            .O(N__54575),
            .I(N__54145));
    InMux I__12689 (
            .O(N__54574),
            .I(N__54145));
    InMux I__12688 (
            .O(N__54573),
            .I(N__54140));
    InMux I__12687 (
            .O(N__54572),
            .I(N__54140));
    InMux I__12686 (
            .O(N__54569),
            .I(N__54131));
    InMux I__12685 (
            .O(N__54566),
            .I(N__54131));
    InMux I__12684 (
            .O(N__54565),
            .I(N__54131));
    InMux I__12683 (
            .O(N__54564),
            .I(N__54131));
    InMux I__12682 (
            .O(N__54561),
            .I(N__54122));
    InMux I__12681 (
            .O(N__54558),
            .I(N__54122));
    InMux I__12680 (
            .O(N__54557),
            .I(N__54122));
    InMux I__12679 (
            .O(N__54556),
            .I(N__54122));
    InMux I__12678 (
            .O(N__54553),
            .I(N__54113));
    InMux I__12677 (
            .O(N__54550),
            .I(N__54113));
    InMux I__12676 (
            .O(N__54547),
            .I(N__54113));
    InMux I__12675 (
            .O(N__54544),
            .I(N__54113));
    InMux I__12674 (
            .O(N__54541),
            .I(N__54106));
    InMux I__12673 (
            .O(N__54538),
            .I(N__54106));
    InMux I__12672 (
            .O(N__54535),
            .I(N__54106));
    InMux I__12671 (
            .O(N__54534),
            .I(N__54095));
    InMux I__12670 (
            .O(N__54531),
            .I(N__54095));
    InMux I__12669 (
            .O(N__54528),
            .I(N__54095));
    InMux I__12668 (
            .O(N__54525),
            .I(N__54095));
    InMux I__12667 (
            .O(N__54522),
            .I(N__54095));
    InMux I__12666 (
            .O(N__54519),
            .I(N__54090));
    InMux I__12665 (
            .O(N__54516),
            .I(N__54090));
    InMux I__12664 (
            .O(N__54515),
            .I(N__54083));
    InMux I__12663 (
            .O(N__54512),
            .I(N__54083));
    InMux I__12662 (
            .O(N__54509),
            .I(N__54083));
    InMux I__12661 (
            .O(N__54508),
            .I(N__54076));
    InMux I__12660 (
            .O(N__54507),
            .I(N__54076));
    InMux I__12659 (
            .O(N__54506),
            .I(N__54076));
    LocalMux I__12658 (
            .O(N__54499),
            .I(N__54067));
    LocalMux I__12657 (
            .O(N__54492),
            .I(N__54067));
    LocalMux I__12656 (
            .O(N__54483),
            .I(N__54067));
    Span4Mux_s2_h I__12655 (
            .O(N__54480),
            .I(N__54058));
    LocalMux I__12654 (
            .O(N__54477),
            .I(N__54058));
    LocalMux I__12653 (
            .O(N__54466),
            .I(N__54058));
    LocalMux I__12652 (
            .O(N__54457),
            .I(N__54058));
    LocalMux I__12651 (
            .O(N__54452),
            .I(N__54053));
    LocalMux I__12650 (
            .O(N__54447),
            .I(N__54053));
    InMux I__12649 (
            .O(N__54446),
            .I(N__54050));
    InMux I__12648 (
            .O(N__54445),
            .I(N__54043));
    InMux I__12647 (
            .O(N__54444),
            .I(N__54043));
    InMux I__12646 (
            .O(N__54443),
            .I(N__54043));
    LocalMux I__12645 (
            .O(N__54438),
            .I(N__54036));
    LocalMux I__12644 (
            .O(N__54431),
            .I(N__54036));
    LocalMux I__12643 (
            .O(N__54424),
            .I(N__54036));
    InMux I__12642 (
            .O(N__54423),
            .I(N__54025));
    InMux I__12641 (
            .O(N__54422),
            .I(N__54025));
    InMux I__12640 (
            .O(N__54421),
            .I(N__54025));
    InMux I__12639 (
            .O(N__54418),
            .I(N__54025));
    InMux I__12638 (
            .O(N__54417),
            .I(N__54025));
    CascadeMux I__12637 (
            .O(N__54416),
            .I(N__54017));
    CascadeMux I__12636 (
            .O(N__54415),
            .I(N__54014));
    CascadeMux I__12635 (
            .O(N__54414),
            .I(N__54011));
    Span4Mux_v I__12634 (
            .O(N__54407),
            .I(N__54001));
    LocalMux I__12633 (
            .O(N__54402),
            .I(N__54001));
    LocalMux I__12632 (
            .O(N__54391),
            .I(N__54001));
    LocalMux I__12631 (
            .O(N__54382),
            .I(N__54001));
    InMux I__12630 (
            .O(N__54381),
            .I(N__53994));
    InMux I__12629 (
            .O(N__54380),
            .I(N__53994));
    InMux I__12628 (
            .O(N__54379),
            .I(N__53994));
    InMux I__12627 (
            .O(N__54376),
            .I(N__53983));
    InMux I__12626 (
            .O(N__54375),
            .I(N__53983));
    InMux I__12625 (
            .O(N__54374),
            .I(N__53983));
    InMux I__12624 (
            .O(N__54373),
            .I(N__53983));
    InMux I__12623 (
            .O(N__54370),
            .I(N__53983));
    CascadeMux I__12622 (
            .O(N__54369),
            .I(N__53979));
    CascadeMux I__12621 (
            .O(N__54368),
            .I(N__53972));
    CascadeMux I__12620 (
            .O(N__54367),
            .I(N__53969));
    LocalMux I__12619 (
            .O(N__54364),
            .I(N__53960));
    LocalMux I__12618 (
            .O(N__54357),
            .I(N__53960));
    LocalMux I__12617 (
            .O(N__54352),
            .I(N__53960));
    InMux I__12616 (
            .O(N__54351),
            .I(N__53957));
    InMux I__12615 (
            .O(N__54348),
            .I(N__53950));
    InMux I__12614 (
            .O(N__54347),
            .I(N__53950));
    InMux I__12613 (
            .O(N__54346),
            .I(N__53950));
    InMux I__12612 (
            .O(N__54345),
            .I(N__53945));
    InMux I__12611 (
            .O(N__54342),
            .I(N__53945));
    InMux I__12610 (
            .O(N__54339),
            .I(N__53936));
    InMux I__12609 (
            .O(N__54336),
            .I(N__53936));
    InMux I__12608 (
            .O(N__54333),
            .I(N__53936));
    InMux I__12607 (
            .O(N__54330),
            .I(N__53936));
    CascadeMux I__12606 (
            .O(N__54329),
            .I(N__53932));
    CascadeMux I__12605 (
            .O(N__54328),
            .I(N__53929));
    CascadeMux I__12604 (
            .O(N__54327),
            .I(N__53926));
    CascadeMux I__12603 (
            .O(N__54326),
            .I(N__53923));
    CascadeMux I__12602 (
            .O(N__54325),
            .I(N__53920));
    InMux I__12601 (
            .O(N__54324),
            .I(N__53910));
    InMux I__12600 (
            .O(N__54321),
            .I(N__53910));
    InMux I__12599 (
            .O(N__54318),
            .I(N__53910));
    InMux I__12598 (
            .O(N__54315),
            .I(N__53903));
    InMux I__12597 (
            .O(N__54312),
            .I(N__53903));
    InMux I__12596 (
            .O(N__54309),
            .I(N__53903));
    Span4Mux_v I__12595 (
            .O(N__54306),
            .I(N__53898));
    LocalMux I__12594 (
            .O(N__54297),
            .I(N__53898));
    InMux I__12593 (
            .O(N__54294),
            .I(N__53891));
    InMux I__12592 (
            .O(N__54293),
            .I(N__53891));
    InMux I__12591 (
            .O(N__54292),
            .I(N__53891));
    InMux I__12590 (
            .O(N__54289),
            .I(N__53880));
    InMux I__12589 (
            .O(N__54288),
            .I(N__53880));
    InMux I__12588 (
            .O(N__54287),
            .I(N__53880));
    InMux I__12587 (
            .O(N__54284),
            .I(N__53880));
    InMux I__12586 (
            .O(N__54283),
            .I(N__53880));
    Span4Mux_h I__12585 (
            .O(N__54280),
            .I(N__53875));
    LocalMux I__12584 (
            .O(N__54275),
            .I(N__53875));
    Span4Mux_h I__12583 (
            .O(N__54270),
            .I(N__53868));
    Span4Mux_h I__12582 (
            .O(N__54263),
            .I(N__53868));
    LocalMux I__12581 (
            .O(N__54258),
            .I(N__53868));
    LocalMux I__12580 (
            .O(N__54253),
            .I(N__53865));
    InMux I__12579 (
            .O(N__54252),
            .I(N__53856));
    InMux I__12578 (
            .O(N__54249),
            .I(N__53856));
    InMux I__12577 (
            .O(N__54248),
            .I(N__53856));
    InMux I__12576 (
            .O(N__54247),
            .I(N__53856));
    CascadeMux I__12575 (
            .O(N__54246),
            .I(N__53852));
    CascadeMux I__12574 (
            .O(N__54245),
            .I(N__53847));
    CascadeMux I__12573 (
            .O(N__54244),
            .I(N__53843));
    CascadeMux I__12572 (
            .O(N__54243),
            .I(N__53838));
    CascadeMux I__12571 (
            .O(N__54242),
            .I(N__53835));
    CascadeMux I__12570 (
            .O(N__54241),
            .I(N__53831));
    CascadeMux I__12569 (
            .O(N__54240),
            .I(N__53828));
    InMux I__12568 (
            .O(N__54237),
            .I(N__53825));
    InMux I__12567 (
            .O(N__54236),
            .I(N__53820));
    InMux I__12566 (
            .O(N__54233),
            .I(N__53820));
    LocalMux I__12565 (
            .O(N__54230),
            .I(N__53810));
    LocalMux I__12564 (
            .O(N__54223),
            .I(N__53799));
    LocalMux I__12563 (
            .O(N__54218),
            .I(N__53799));
    LocalMux I__12562 (
            .O(N__54215),
            .I(N__53799));
    LocalMux I__12561 (
            .O(N__54212),
            .I(N__53799));
    LocalMux I__12560 (
            .O(N__54205),
            .I(N__53799));
    Span4Mux_h I__12559 (
            .O(N__54186),
            .I(N__53792));
    LocalMux I__12558 (
            .O(N__54177),
            .I(N__53792));
    LocalMux I__12557 (
            .O(N__54168),
            .I(N__53792));
    LocalMux I__12556 (
            .O(N__54163),
            .I(N__53778));
    LocalMux I__12555 (
            .O(N__54154),
            .I(N__53778));
    LocalMux I__12554 (
            .O(N__54145),
            .I(N__53778));
    LocalMux I__12553 (
            .O(N__54140),
            .I(N__53761));
    LocalMux I__12552 (
            .O(N__54131),
            .I(N__53761));
    LocalMux I__12551 (
            .O(N__54122),
            .I(N__53761));
    LocalMux I__12550 (
            .O(N__54113),
            .I(N__53761));
    LocalMux I__12549 (
            .O(N__54106),
            .I(N__53761));
    LocalMux I__12548 (
            .O(N__54095),
            .I(N__53761));
    LocalMux I__12547 (
            .O(N__54090),
            .I(N__53761));
    LocalMux I__12546 (
            .O(N__54083),
            .I(N__53761));
    LocalMux I__12545 (
            .O(N__54076),
            .I(N__53758));
    InMux I__12544 (
            .O(N__54075),
            .I(N__53753));
    InMux I__12543 (
            .O(N__54074),
            .I(N__53753));
    Span4Mux_v I__12542 (
            .O(N__54067),
            .I(N__53742));
    Span4Mux_v I__12541 (
            .O(N__54058),
            .I(N__53742));
    Span4Mux_s2_h I__12540 (
            .O(N__54053),
            .I(N__53742));
    LocalMux I__12539 (
            .O(N__54050),
            .I(N__53742));
    LocalMux I__12538 (
            .O(N__54043),
            .I(N__53742));
    Span4Mux_v I__12537 (
            .O(N__54036),
            .I(N__53737));
    LocalMux I__12536 (
            .O(N__54025),
            .I(N__53737));
    InMux I__12535 (
            .O(N__54024),
            .I(N__53728));
    InMux I__12534 (
            .O(N__54023),
            .I(N__53728));
    InMux I__12533 (
            .O(N__54022),
            .I(N__53728));
    InMux I__12532 (
            .O(N__54021),
            .I(N__53728));
    InMux I__12531 (
            .O(N__54020),
            .I(N__53717));
    InMux I__12530 (
            .O(N__54017),
            .I(N__53717));
    InMux I__12529 (
            .O(N__54014),
            .I(N__53717));
    InMux I__12528 (
            .O(N__54011),
            .I(N__53717));
    InMux I__12527 (
            .O(N__54010),
            .I(N__53717));
    Span4Mux_v I__12526 (
            .O(N__54001),
            .I(N__53710));
    LocalMux I__12525 (
            .O(N__53994),
            .I(N__53710));
    LocalMux I__12524 (
            .O(N__53983),
            .I(N__53710));
    InMux I__12523 (
            .O(N__53982),
            .I(N__53705));
    InMux I__12522 (
            .O(N__53979),
            .I(N__53705));
    InMux I__12521 (
            .O(N__53978),
            .I(N__53696));
    InMux I__12520 (
            .O(N__53977),
            .I(N__53696));
    InMux I__12519 (
            .O(N__53976),
            .I(N__53696));
    InMux I__12518 (
            .O(N__53975),
            .I(N__53696));
    InMux I__12517 (
            .O(N__53972),
            .I(N__53689));
    InMux I__12516 (
            .O(N__53969),
            .I(N__53689));
    InMux I__12515 (
            .O(N__53968),
            .I(N__53689));
    InMux I__12514 (
            .O(N__53967),
            .I(N__53686));
    Span4Mux_h I__12513 (
            .O(N__53960),
            .I(N__53677));
    LocalMux I__12512 (
            .O(N__53957),
            .I(N__53677));
    LocalMux I__12511 (
            .O(N__53950),
            .I(N__53677));
    LocalMux I__12510 (
            .O(N__53945),
            .I(N__53677));
    LocalMux I__12509 (
            .O(N__53936),
            .I(N__53674));
    InMux I__12508 (
            .O(N__53935),
            .I(N__53667));
    InMux I__12507 (
            .O(N__53932),
            .I(N__53667));
    InMux I__12506 (
            .O(N__53929),
            .I(N__53667));
    InMux I__12505 (
            .O(N__53926),
            .I(N__53660));
    InMux I__12504 (
            .O(N__53923),
            .I(N__53660));
    InMux I__12503 (
            .O(N__53920),
            .I(N__53660));
    CascadeMux I__12502 (
            .O(N__53919),
            .I(N__53656));
    CascadeMux I__12501 (
            .O(N__53918),
            .I(N__53653));
    CascadeMux I__12500 (
            .O(N__53917),
            .I(N__53650));
    LocalMux I__12499 (
            .O(N__53910),
            .I(N__53635));
    LocalMux I__12498 (
            .O(N__53903),
            .I(N__53635));
    Sp12to4 I__12497 (
            .O(N__53898),
            .I(N__53635));
    LocalMux I__12496 (
            .O(N__53891),
            .I(N__53635));
    LocalMux I__12495 (
            .O(N__53880),
            .I(N__53635));
    Span4Mux_h I__12494 (
            .O(N__53875),
            .I(N__53630));
    Span4Mux_v I__12493 (
            .O(N__53868),
            .I(N__53630));
    Span4Mux_v I__12492 (
            .O(N__53865),
            .I(N__53625));
    LocalMux I__12491 (
            .O(N__53856),
            .I(N__53625));
    InMux I__12490 (
            .O(N__53855),
            .I(N__53616));
    InMux I__12489 (
            .O(N__53852),
            .I(N__53616));
    InMux I__12488 (
            .O(N__53851),
            .I(N__53616));
    InMux I__12487 (
            .O(N__53850),
            .I(N__53616));
    InMux I__12486 (
            .O(N__53847),
            .I(N__53605));
    InMux I__12485 (
            .O(N__53846),
            .I(N__53605));
    InMux I__12484 (
            .O(N__53843),
            .I(N__53605));
    InMux I__12483 (
            .O(N__53842),
            .I(N__53605));
    InMux I__12482 (
            .O(N__53841),
            .I(N__53605));
    InMux I__12481 (
            .O(N__53838),
            .I(N__53594));
    InMux I__12480 (
            .O(N__53835),
            .I(N__53594));
    InMux I__12479 (
            .O(N__53834),
            .I(N__53594));
    InMux I__12478 (
            .O(N__53831),
            .I(N__53594));
    InMux I__12477 (
            .O(N__53828),
            .I(N__53594));
    LocalMux I__12476 (
            .O(N__53825),
            .I(N__53589));
    LocalMux I__12475 (
            .O(N__53820),
            .I(N__53589));
    InMux I__12474 (
            .O(N__53819),
            .I(N__53586));
    InMux I__12473 (
            .O(N__53818),
            .I(N__53579));
    InMux I__12472 (
            .O(N__53817),
            .I(N__53579));
    InMux I__12471 (
            .O(N__53816),
            .I(N__53579));
    InMux I__12470 (
            .O(N__53815),
            .I(N__53572));
    InMux I__12469 (
            .O(N__53814),
            .I(N__53572));
    InMux I__12468 (
            .O(N__53813),
            .I(N__53572));
    Span4Mux_v I__12467 (
            .O(N__53810),
            .I(N__53565));
    Span4Mux_v I__12466 (
            .O(N__53799),
            .I(N__53565));
    Span4Mux_v I__12465 (
            .O(N__53792),
            .I(N__53565));
    InMux I__12464 (
            .O(N__53791),
            .I(N__53562));
    InMux I__12463 (
            .O(N__53790),
            .I(N__53557));
    InMux I__12462 (
            .O(N__53789),
            .I(N__53557));
    InMux I__12461 (
            .O(N__53788),
            .I(N__53552));
    InMux I__12460 (
            .O(N__53787),
            .I(N__53552));
    InMux I__12459 (
            .O(N__53786),
            .I(N__53547));
    InMux I__12458 (
            .O(N__53785),
            .I(N__53547));
    Span4Mux_v I__12457 (
            .O(N__53778),
            .I(N__53542));
    Span4Mux_v I__12456 (
            .O(N__53761),
            .I(N__53542));
    Span4Mux_v I__12455 (
            .O(N__53758),
            .I(N__53537));
    LocalMux I__12454 (
            .O(N__53753),
            .I(N__53537));
    Span4Mux_h I__12453 (
            .O(N__53742),
            .I(N__53528));
    Span4Mux_v I__12452 (
            .O(N__53737),
            .I(N__53528));
    LocalMux I__12451 (
            .O(N__53728),
            .I(N__53528));
    LocalMux I__12450 (
            .O(N__53717),
            .I(N__53528));
    Span4Mux_v I__12449 (
            .O(N__53710),
            .I(N__53519));
    LocalMux I__12448 (
            .O(N__53705),
            .I(N__53519));
    LocalMux I__12447 (
            .O(N__53696),
            .I(N__53519));
    LocalMux I__12446 (
            .O(N__53689),
            .I(N__53519));
    LocalMux I__12445 (
            .O(N__53686),
            .I(N__53516));
    Span4Mux_v I__12444 (
            .O(N__53677),
            .I(N__53513));
    Span4Mux_v I__12443 (
            .O(N__53674),
            .I(N__53506));
    LocalMux I__12442 (
            .O(N__53667),
            .I(N__53506));
    LocalMux I__12441 (
            .O(N__53660),
            .I(N__53506));
    InMux I__12440 (
            .O(N__53659),
            .I(N__53497));
    InMux I__12439 (
            .O(N__53656),
            .I(N__53497));
    InMux I__12438 (
            .O(N__53653),
            .I(N__53497));
    InMux I__12437 (
            .O(N__53650),
            .I(N__53497));
    CascadeMux I__12436 (
            .O(N__53649),
            .I(N__53494));
    CascadeMux I__12435 (
            .O(N__53648),
            .I(N__53491));
    CascadeMux I__12434 (
            .O(N__53647),
            .I(N__53488));
    CascadeMux I__12433 (
            .O(N__53646),
            .I(N__53485));
    Span12Mux_v I__12432 (
            .O(N__53635),
            .I(N__53482));
    Span4Mux_v I__12431 (
            .O(N__53630),
            .I(N__53477));
    Span4Mux_v I__12430 (
            .O(N__53625),
            .I(N__53477));
    LocalMux I__12429 (
            .O(N__53616),
            .I(N__53472));
    LocalMux I__12428 (
            .O(N__53605),
            .I(N__53472));
    LocalMux I__12427 (
            .O(N__53594),
            .I(N__53461));
    Span12Mux_s8_v I__12426 (
            .O(N__53589),
            .I(N__53461));
    LocalMux I__12425 (
            .O(N__53586),
            .I(N__53461));
    LocalMux I__12424 (
            .O(N__53579),
            .I(N__53461));
    LocalMux I__12423 (
            .O(N__53572),
            .I(N__53461));
    Sp12to4 I__12422 (
            .O(N__53565),
            .I(N__53450));
    LocalMux I__12421 (
            .O(N__53562),
            .I(N__53450));
    LocalMux I__12420 (
            .O(N__53557),
            .I(N__53450));
    LocalMux I__12419 (
            .O(N__53552),
            .I(N__53450));
    LocalMux I__12418 (
            .O(N__53547),
            .I(N__53450));
    Span4Mux_h I__12417 (
            .O(N__53542),
            .I(N__53445));
    Span4Mux_v I__12416 (
            .O(N__53537),
            .I(N__53445));
    Span4Mux_v I__12415 (
            .O(N__53528),
            .I(N__53440));
    Span4Mux_v I__12414 (
            .O(N__53519),
            .I(N__53440));
    Span12Mux_s4_h I__12413 (
            .O(N__53516),
            .I(N__53435));
    Sp12to4 I__12412 (
            .O(N__53513),
            .I(N__53435));
    Span4Mux_h I__12411 (
            .O(N__53506),
            .I(N__53430));
    LocalMux I__12410 (
            .O(N__53497),
            .I(N__53430));
    InMux I__12409 (
            .O(N__53494),
            .I(N__53421));
    InMux I__12408 (
            .O(N__53491),
            .I(N__53421));
    InMux I__12407 (
            .O(N__53488),
            .I(N__53421));
    InMux I__12406 (
            .O(N__53485),
            .I(N__53421));
    Span12Mux_h I__12405 (
            .O(N__53482),
            .I(N__53418));
    Span4Mux_v I__12404 (
            .O(N__53477),
            .I(N__53415));
    Span12Mux_v I__12403 (
            .O(N__53472),
            .I(N__53408));
    Span12Mux_h I__12402 (
            .O(N__53461),
            .I(N__53408));
    Span12Mux_h I__12401 (
            .O(N__53450),
            .I(N__53408));
    Span4Mux_h I__12400 (
            .O(N__53445),
            .I(N__53403));
    Span4Mux_h I__12399 (
            .O(N__53440),
            .I(N__53403));
    Span12Mux_v I__12398 (
            .O(N__53435),
            .I(N__53396));
    Sp12to4 I__12397 (
            .O(N__53430),
            .I(N__53396));
    LocalMux I__12396 (
            .O(N__53421),
            .I(N__53396));
    Odrv12 I__12395 (
            .O(N__53418),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__12394 (
            .O(N__53415),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__12393 (
            .O(N__53408),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__12392 (
            .O(N__53403),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__12391 (
            .O(N__53396),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__12390 (
            .O(N__53385),
            .I(N__53381));
    CascadeMux I__12389 (
            .O(N__53384),
            .I(N__53378));
    InMux I__12388 (
            .O(N__53381),
            .I(N__53374));
    InMux I__12387 (
            .O(N__53378),
            .I(N__53371));
    InMux I__12386 (
            .O(N__53377),
            .I(N__53368));
    LocalMux I__12385 (
            .O(N__53374),
            .I(N__53365));
    LocalMux I__12384 (
            .O(N__53371),
            .I(n1026));
    LocalMux I__12383 (
            .O(N__53368),
            .I(n1026));
    Odrv12 I__12382 (
            .O(N__53365),
            .I(n1026));
    InMux I__12381 (
            .O(N__53358),
            .I(bfn_16_24_0_));
    InMux I__12380 (
            .O(N__53355),
            .I(N__53352));
    LocalMux I__12379 (
            .O(N__53352),
            .I(N__53349));
    Odrv4 I__12378 (
            .O(N__53349),
            .I(n1093));
    InMux I__12377 (
            .O(N__53346),
            .I(N__53342));
    InMux I__12376 (
            .O(N__53345),
            .I(N__53339));
    LocalMux I__12375 (
            .O(N__53342),
            .I(N__53336));
    LocalMux I__12374 (
            .O(N__53339),
            .I(sweep_counter_0));
    Odrv4 I__12373 (
            .O(N__53336),
            .I(sweep_counter_0));
    InMux I__12372 (
            .O(N__53331),
            .I(bfn_16_25_0_));
    InMux I__12371 (
            .O(N__53328),
            .I(N__53324));
    InMux I__12370 (
            .O(N__53327),
            .I(N__53321));
    LocalMux I__12369 (
            .O(N__53324),
            .I(N__53318));
    LocalMux I__12368 (
            .O(N__53321),
            .I(sweep_counter_1));
    Odrv4 I__12367 (
            .O(N__53318),
            .I(sweep_counter_1));
    InMux I__12366 (
            .O(N__53313),
            .I(n13053));
    InMux I__12365 (
            .O(N__53310),
            .I(N__53306));
    InMux I__12364 (
            .O(N__53309),
            .I(N__53303));
    LocalMux I__12363 (
            .O(N__53306),
            .I(N__53300));
    LocalMux I__12362 (
            .O(N__53303),
            .I(N__53295));
    Span4Mux_v I__12361 (
            .O(N__53300),
            .I(N__53295));
    Odrv4 I__12360 (
            .O(N__53295),
            .I(sweep_counter_2));
    InMux I__12359 (
            .O(N__53292),
            .I(n13054));
    InMux I__12358 (
            .O(N__53289),
            .I(N__53286));
    LocalMux I__12357 (
            .O(N__53286),
            .I(N__53282));
    InMux I__12356 (
            .O(N__53285),
            .I(N__53279));
    Span4Mux_v I__12355 (
            .O(N__53282),
            .I(N__53276));
    LocalMux I__12354 (
            .O(N__53279),
            .I(sweep_counter_3));
    Odrv4 I__12353 (
            .O(N__53276),
            .I(sweep_counter_3));
    InMux I__12352 (
            .O(N__53271),
            .I(n13055));
    InMux I__12351 (
            .O(N__53268),
            .I(N__53265));
    LocalMux I__12350 (
            .O(N__53265),
            .I(N__53261));
    InMux I__12349 (
            .O(N__53264),
            .I(N__53258));
    Span4Mux_h I__12348 (
            .O(N__53261),
            .I(N__53255));
    LocalMux I__12347 (
            .O(N__53258),
            .I(sweep_counter_4));
    Odrv4 I__12346 (
            .O(N__53255),
            .I(sweep_counter_4));
    InMux I__12345 (
            .O(N__53250),
            .I(n13056));
    InMux I__12344 (
            .O(N__53247),
            .I(N__53243));
    InMux I__12343 (
            .O(N__53246),
            .I(N__53240));
    LocalMux I__12342 (
            .O(N__53243),
            .I(N__53237));
    LocalMux I__12341 (
            .O(N__53240),
            .I(sweep_counter_5));
    Odrv4 I__12340 (
            .O(N__53237),
            .I(sweep_counter_5));
    InMux I__12339 (
            .O(N__53232),
            .I(n13057));
    InMux I__12338 (
            .O(N__53229),
            .I(N__53226));
    LocalMux I__12337 (
            .O(N__53226),
            .I(n1298));
    CascadeMux I__12336 (
            .O(N__53223),
            .I(N__53218));
    CascadeMux I__12335 (
            .O(N__53222),
            .I(N__53215));
    CascadeMux I__12334 (
            .O(N__53221),
            .I(N__53212));
    InMux I__12333 (
            .O(N__53218),
            .I(N__53209));
    InMux I__12332 (
            .O(N__53215),
            .I(N__53206));
    InMux I__12331 (
            .O(N__53212),
            .I(N__53203));
    LocalMux I__12330 (
            .O(N__53209),
            .I(N__53200));
    LocalMux I__12329 (
            .O(N__53206),
            .I(n1231));
    LocalMux I__12328 (
            .O(N__53203),
            .I(n1231));
    Odrv4 I__12327 (
            .O(N__53200),
            .I(n1231));
    CascadeMux I__12326 (
            .O(N__53193),
            .I(N__53190));
    InMux I__12325 (
            .O(N__53190),
            .I(N__53187));
    LocalMux I__12324 (
            .O(N__53187),
            .I(N__53184));
    Span4Mux_v I__12323 (
            .O(N__53184),
            .I(N__53181));
    Span4Mux_h I__12322 (
            .O(N__53181),
            .I(N__53176));
    CascadeMux I__12321 (
            .O(N__53180),
            .I(N__53168));
    CascadeMux I__12320 (
            .O(N__53179),
            .I(N__53163));
    Span4Mux_h I__12319 (
            .O(N__53176),
            .I(N__53159));
    InMux I__12318 (
            .O(N__53175),
            .I(N__53156));
    InMux I__12317 (
            .O(N__53174),
            .I(N__53153));
    InMux I__12316 (
            .O(N__53173),
            .I(N__53150));
    InMux I__12315 (
            .O(N__53172),
            .I(N__53145));
    InMux I__12314 (
            .O(N__53171),
            .I(N__53145));
    InMux I__12313 (
            .O(N__53168),
            .I(N__53134));
    InMux I__12312 (
            .O(N__53167),
            .I(N__53134));
    InMux I__12311 (
            .O(N__53166),
            .I(N__53134));
    InMux I__12310 (
            .O(N__53163),
            .I(N__53134));
    InMux I__12309 (
            .O(N__53162),
            .I(N__53134));
    Odrv4 I__12308 (
            .O(N__53159),
            .I(n1257));
    LocalMux I__12307 (
            .O(N__53156),
            .I(n1257));
    LocalMux I__12306 (
            .O(N__53153),
            .I(n1257));
    LocalMux I__12305 (
            .O(N__53150),
            .I(n1257));
    LocalMux I__12304 (
            .O(N__53145),
            .I(n1257));
    LocalMux I__12303 (
            .O(N__53134),
            .I(n1257));
    CascadeMux I__12302 (
            .O(N__53121),
            .I(N__53118));
    InMux I__12301 (
            .O(N__53118),
            .I(N__53115));
    LocalMux I__12300 (
            .O(N__53115),
            .I(N__53110));
    InMux I__12299 (
            .O(N__53114),
            .I(N__53107));
    InMux I__12298 (
            .O(N__53113),
            .I(N__53104));
    Span4Mux_h I__12297 (
            .O(N__53110),
            .I(N__53101));
    LocalMux I__12296 (
            .O(N__53107),
            .I(N__53096));
    LocalMux I__12295 (
            .O(N__53104),
            .I(N__53096));
    Odrv4 I__12294 (
            .O(N__53101),
            .I(n1330));
    Odrv4 I__12293 (
            .O(N__53096),
            .I(n1330));
    InMux I__12292 (
            .O(N__53091),
            .I(N__53088));
    LocalMux I__12291 (
            .O(N__53088),
            .I(N__53085));
    Span4Mux_v I__12290 (
            .O(N__53085),
            .I(N__53080));
    InMux I__12289 (
            .O(N__53084),
            .I(N__53075));
    InMux I__12288 (
            .O(N__53083),
            .I(N__53075));
    Odrv4 I__12287 (
            .O(N__53080),
            .I(n296));
    LocalMux I__12286 (
            .O(N__53075),
            .I(n296));
    InMux I__12285 (
            .O(N__53070),
            .I(N__53067));
    LocalMux I__12284 (
            .O(N__53067),
            .I(N__53064));
    Span4Mux_h I__12283 (
            .O(N__53064),
            .I(N__53061));
    Odrv4 I__12282 (
            .O(N__53061),
            .I(n1101));
    InMux I__12281 (
            .O(N__53058),
            .I(bfn_16_23_0_));
    CascadeMux I__12280 (
            .O(N__53055),
            .I(N__53052));
    InMux I__12279 (
            .O(N__53052),
            .I(N__53047));
    InMux I__12278 (
            .O(N__53051),
            .I(N__53042));
    InMux I__12277 (
            .O(N__53050),
            .I(N__53042));
    LocalMux I__12276 (
            .O(N__53047),
            .I(N__53039));
    LocalMux I__12275 (
            .O(N__53042),
            .I(n1033));
    Odrv12 I__12274 (
            .O(N__53039),
            .I(n1033));
    InMux I__12273 (
            .O(N__53034),
            .I(N__53031));
    LocalMux I__12272 (
            .O(N__53031),
            .I(N__53028));
    Odrv12 I__12271 (
            .O(N__53028),
            .I(n1100));
    InMux I__12270 (
            .O(N__53025),
            .I(n12514));
    CascadeMux I__12269 (
            .O(N__53022),
            .I(N__53018));
    CascadeMux I__12268 (
            .O(N__53021),
            .I(N__53014));
    InMux I__12267 (
            .O(N__53018),
            .I(N__53011));
    InMux I__12266 (
            .O(N__53017),
            .I(N__53008));
    InMux I__12265 (
            .O(N__53014),
            .I(N__53005));
    LocalMux I__12264 (
            .O(N__53011),
            .I(N__53002));
    LocalMux I__12263 (
            .O(N__53008),
            .I(n1032));
    LocalMux I__12262 (
            .O(N__53005),
            .I(n1032));
    Odrv12 I__12261 (
            .O(N__53002),
            .I(n1032));
    InMux I__12260 (
            .O(N__52995),
            .I(N__52992));
    LocalMux I__12259 (
            .O(N__52992),
            .I(N__52989));
    Span4Mux_h I__12258 (
            .O(N__52989),
            .I(N__52986));
    Odrv4 I__12257 (
            .O(N__52986),
            .I(n1099));
    InMux I__12256 (
            .O(N__52983),
            .I(n12515));
    CascadeMux I__12255 (
            .O(N__52980),
            .I(N__52976));
    CascadeMux I__12254 (
            .O(N__52979),
            .I(N__52973));
    InMux I__12253 (
            .O(N__52976),
            .I(N__52969));
    InMux I__12252 (
            .O(N__52973),
            .I(N__52966));
    InMux I__12251 (
            .O(N__52972),
            .I(N__52963));
    LocalMux I__12250 (
            .O(N__52969),
            .I(N__52960));
    LocalMux I__12249 (
            .O(N__52966),
            .I(n1031));
    LocalMux I__12248 (
            .O(N__52963),
            .I(n1031));
    Odrv12 I__12247 (
            .O(N__52960),
            .I(n1031));
    InMux I__12246 (
            .O(N__52953),
            .I(N__52950));
    LocalMux I__12245 (
            .O(N__52950),
            .I(N__52947));
    Span4Mux_h I__12244 (
            .O(N__52947),
            .I(N__52944));
    Odrv4 I__12243 (
            .O(N__52944),
            .I(n1098));
    InMux I__12242 (
            .O(N__52941),
            .I(n12516));
    CascadeMux I__12241 (
            .O(N__52938),
            .I(N__52934));
    CascadeMux I__12240 (
            .O(N__52937),
            .I(N__52931));
    InMux I__12239 (
            .O(N__52934),
            .I(N__52927));
    InMux I__12238 (
            .O(N__52931),
            .I(N__52924));
    InMux I__12237 (
            .O(N__52930),
            .I(N__52921));
    LocalMux I__12236 (
            .O(N__52927),
            .I(N__52918));
    LocalMux I__12235 (
            .O(N__52924),
            .I(n1030));
    LocalMux I__12234 (
            .O(N__52921),
            .I(n1030));
    Odrv4 I__12233 (
            .O(N__52918),
            .I(n1030));
    InMux I__12232 (
            .O(N__52911),
            .I(N__52908));
    LocalMux I__12231 (
            .O(N__52908),
            .I(N__52905));
    Span4Mux_h I__12230 (
            .O(N__52905),
            .I(N__52902));
    Odrv4 I__12229 (
            .O(N__52902),
            .I(n1097));
    InMux I__12228 (
            .O(N__52899),
            .I(n12517));
    CascadeMux I__12227 (
            .O(N__52896),
            .I(N__52892));
    InMux I__12226 (
            .O(N__52895),
            .I(N__52889));
    InMux I__12225 (
            .O(N__52892),
            .I(N__52886));
    LocalMux I__12224 (
            .O(N__52889),
            .I(N__52880));
    LocalMux I__12223 (
            .O(N__52886),
            .I(N__52880));
    InMux I__12222 (
            .O(N__52885),
            .I(N__52877));
    Span4Mux_h I__12221 (
            .O(N__52880),
            .I(N__52874));
    LocalMux I__12220 (
            .O(N__52877),
            .I(n1029));
    Odrv4 I__12219 (
            .O(N__52874),
            .I(n1029));
    InMux I__12218 (
            .O(N__52869),
            .I(N__52866));
    LocalMux I__12217 (
            .O(N__52866),
            .I(n1096));
    InMux I__12216 (
            .O(N__52863),
            .I(n12518));
    CascadeMux I__12215 (
            .O(N__52860),
            .I(N__52856));
    InMux I__12214 (
            .O(N__52859),
            .I(N__52853));
    InMux I__12213 (
            .O(N__52856),
            .I(N__52849));
    LocalMux I__12212 (
            .O(N__52853),
            .I(N__52846));
    InMux I__12211 (
            .O(N__52852),
            .I(N__52843));
    LocalMux I__12210 (
            .O(N__52849),
            .I(N__52840));
    Odrv4 I__12209 (
            .O(N__52846),
            .I(n1028));
    LocalMux I__12208 (
            .O(N__52843),
            .I(n1028));
    Odrv12 I__12207 (
            .O(N__52840),
            .I(n1028));
    InMux I__12206 (
            .O(N__52833),
            .I(N__52830));
    LocalMux I__12205 (
            .O(N__52830),
            .I(n1095));
    InMux I__12204 (
            .O(N__52827),
            .I(n12519));
    InMux I__12203 (
            .O(N__52824),
            .I(n12533));
    CascadeMux I__12202 (
            .O(N__52821),
            .I(N__52817));
    CascadeMux I__12201 (
            .O(N__52820),
            .I(N__52814));
    InMux I__12200 (
            .O(N__52817),
            .I(N__52810));
    InMux I__12199 (
            .O(N__52814),
            .I(N__52807));
    InMux I__12198 (
            .O(N__52813),
            .I(N__52804));
    LocalMux I__12197 (
            .O(N__52810),
            .I(N__52799));
    LocalMux I__12196 (
            .O(N__52807),
            .I(N__52799));
    LocalMux I__12195 (
            .O(N__52804),
            .I(n1230));
    Odrv4 I__12194 (
            .O(N__52799),
            .I(n1230));
    InMux I__12193 (
            .O(N__52794),
            .I(N__52791));
    LocalMux I__12192 (
            .O(N__52791),
            .I(n1297));
    InMux I__12191 (
            .O(N__52788),
            .I(n12534));
    CascadeMux I__12190 (
            .O(N__52785),
            .I(N__52782));
    InMux I__12189 (
            .O(N__52782),
            .I(N__52778));
    InMux I__12188 (
            .O(N__52781),
            .I(N__52775));
    LocalMux I__12187 (
            .O(N__52778),
            .I(N__52771));
    LocalMux I__12186 (
            .O(N__52775),
            .I(N__52768));
    InMux I__12185 (
            .O(N__52774),
            .I(N__52765));
    Span4Mux_h I__12184 (
            .O(N__52771),
            .I(N__52762));
    Odrv4 I__12183 (
            .O(N__52768),
            .I(n1229));
    LocalMux I__12182 (
            .O(N__52765),
            .I(n1229));
    Odrv4 I__12181 (
            .O(N__52762),
            .I(n1229));
    InMux I__12180 (
            .O(N__52755),
            .I(N__52752));
    LocalMux I__12179 (
            .O(N__52752),
            .I(n1296));
    InMux I__12178 (
            .O(N__52749),
            .I(n12535));
    CascadeMux I__12177 (
            .O(N__52746),
            .I(N__52742));
    CascadeMux I__12176 (
            .O(N__52745),
            .I(N__52739));
    InMux I__12175 (
            .O(N__52742),
            .I(N__52736));
    InMux I__12174 (
            .O(N__52739),
            .I(N__52733));
    LocalMux I__12173 (
            .O(N__52736),
            .I(N__52727));
    LocalMux I__12172 (
            .O(N__52733),
            .I(N__52727));
    InMux I__12171 (
            .O(N__52732),
            .I(N__52724));
    Odrv4 I__12170 (
            .O(N__52727),
            .I(n1228));
    LocalMux I__12169 (
            .O(N__52724),
            .I(n1228));
    InMux I__12168 (
            .O(N__52719),
            .I(N__52716));
    LocalMux I__12167 (
            .O(N__52716),
            .I(n1295));
    InMux I__12166 (
            .O(N__52713),
            .I(n12536));
    CascadeMux I__12165 (
            .O(N__52710),
            .I(N__52706));
    CascadeMux I__12164 (
            .O(N__52709),
            .I(N__52703));
    InMux I__12163 (
            .O(N__52706),
            .I(N__52700));
    InMux I__12162 (
            .O(N__52703),
            .I(N__52697));
    LocalMux I__12161 (
            .O(N__52700),
            .I(n1227));
    LocalMux I__12160 (
            .O(N__52697),
            .I(n1227));
    InMux I__12159 (
            .O(N__52692),
            .I(N__52689));
    LocalMux I__12158 (
            .O(N__52689),
            .I(n1294));
    InMux I__12157 (
            .O(N__52686),
            .I(n12537));
    CascadeMux I__12156 (
            .O(N__52683),
            .I(N__52680));
    InMux I__12155 (
            .O(N__52680),
            .I(N__52675));
    InMux I__12154 (
            .O(N__52679),
            .I(N__52670));
    InMux I__12153 (
            .O(N__52678),
            .I(N__52670));
    LocalMux I__12152 (
            .O(N__52675),
            .I(n1226));
    LocalMux I__12151 (
            .O(N__52670),
            .I(n1226));
    InMux I__12150 (
            .O(N__52665),
            .I(N__52662));
    LocalMux I__12149 (
            .O(N__52662),
            .I(n1293));
    InMux I__12148 (
            .O(N__52659),
            .I(bfn_16_22_0_));
    CascadeMux I__12147 (
            .O(N__52656),
            .I(N__52653));
    InMux I__12146 (
            .O(N__52653),
            .I(N__52649));
    InMux I__12145 (
            .O(N__52652),
            .I(N__52646));
    LocalMux I__12144 (
            .O(N__52649),
            .I(n1225));
    LocalMux I__12143 (
            .O(N__52646),
            .I(n1225));
    InMux I__12142 (
            .O(N__52641),
            .I(N__52638));
    LocalMux I__12141 (
            .O(N__52638),
            .I(n1292));
    InMux I__12140 (
            .O(N__52635),
            .I(n12539));
    InMux I__12139 (
            .O(N__52632),
            .I(N__52629));
    LocalMux I__12138 (
            .O(N__52629),
            .I(N__52626));
    Span4Mux_v I__12137 (
            .O(N__52626),
            .I(N__52623));
    Span4Mux_h I__12136 (
            .O(N__52623),
            .I(N__52620));
    Span4Mux_h I__12135 (
            .O(N__52620),
            .I(N__52616));
    InMux I__12134 (
            .O(N__52619),
            .I(N__52613));
    Odrv4 I__12133 (
            .O(N__52616),
            .I(n15537));
    LocalMux I__12132 (
            .O(N__52613),
            .I(n15537));
    CascadeMux I__12131 (
            .O(N__52608),
            .I(N__52605));
    InMux I__12130 (
            .O(N__52605),
            .I(N__52602));
    LocalMux I__12129 (
            .O(N__52602),
            .I(N__52598));
    InMux I__12128 (
            .O(N__52601),
            .I(N__52595));
    Span4Mux_h I__12127 (
            .O(N__52598),
            .I(N__52592));
    LocalMux I__12126 (
            .O(N__52595),
            .I(N__52589));
    Odrv4 I__12125 (
            .O(N__52592),
            .I(n1224));
    Odrv4 I__12124 (
            .O(N__52589),
            .I(n1224));
    InMux I__12123 (
            .O(N__52584),
            .I(n12540));
    CascadeMux I__12122 (
            .O(N__52581),
            .I(N__52578));
    InMux I__12121 (
            .O(N__52578),
            .I(N__52574));
    CascadeMux I__12120 (
            .O(N__52577),
            .I(N__52571));
    LocalMux I__12119 (
            .O(N__52574),
            .I(N__52568));
    InMux I__12118 (
            .O(N__52571),
            .I(N__52565));
    Span4Mux_h I__12117 (
            .O(N__52568),
            .I(N__52562));
    LocalMux I__12116 (
            .O(N__52565),
            .I(N__52559));
    Odrv4 I__12115 (
            .O(N__52562),
            .I(n1323));
    Odrv4 I__12114 (
            .O(N__52559),
            .I(n1323));
    InMux I__12113 (
            .O(N__52554),
            .I(N__52551));
    LocalMux I__12112 (
            .O(N__52551),
            .I(N__52548));
    Span4Mux_v I__12111 (
            .O(N__52548),
            .I(N__52545));
    Span4Mux_h I__12110 (
            .O(N__52545),
            .I(N__52542));
    Odrv4 I__12109 (
            .O(N__52542),
            .I(n1590));
    InMux I__12108 (
            .O(N__52539),
            .I(n12574));
    InMux I__12107 (
            .O(N__52536),
            .I(N__52533));
    LocalMux I__12106 (
            .O(N__52533),
            .I(N__52529));
    InMux I__12105 (
            .O(N__52532),
            .I(N__52526));
    Span4Mux_v I__12104 (
            .O(N__52529),
            .I(N__52522));
    LocalMux I__12103 (
            .O(N__52526),
            .I(N__52519));
    InMux I__12102 (
            .O(N__52525),
            .I(N__52516));
    Odrv4 I__12101 (
            .O(N__52522),
            .I(n1522));
    Odrv4 I__12100 (
            .O(N__52519),
            .I(n1522));
    LocalMux I__12099 (
            .O(N__52516),
            .I(n1522));
    InMux I__12098 (
            .O(N__52509),
            .I(N__52506));
    LocalMux I__12097 (
            .O(N__52506),
            .I(N__52503));
    Odrv4 I__12096 (
            .O(N__52503),
            .I(n1589));
    InMux I__12095 (
            .O(N__52500),
            .I(n12575));
    InMux I__12094 (
            .O(N__52497),
            .I(N__52493));
    InMux I__12093 (
            .O(N__52496),
            .I(N__52490));
    LocalMux I__12092 (
            .O(N__52493),
            .I(N__52487));
    LocalMux I__12091 (
            .O(N__52490),
            .I(N__52484));
    Odrv4 I__12090 (
            .O(N__52487),
            .I(n1521));
    Odrv4 I__12089 (
            .O(N__52484),
            .I(n1521));
    InMux I__12088 (
            .O(N__52479),
            .I(N__52476));
    LocalMux I__12087 (
            .O(N__52476),
            .I(N__52472));
    CascadeMux I__12086 (
            .O(N__52475),
            .I(N__52469));
    Span4Mux_v I__12085 (
            .O(N__52472),
            .I(N__52466));
    InMux I__12084 (
            .O(N__52469),
            .I(N__52463));
    Sp12to4 I__12083 (
            .O(N__52466),
            .I(N__52460));
    LocalMux I__12082 (
            .O(N__52463),
            .I(N__52457));
    Span12Mux_h I__12081 (
            .O(N__52460),
            .I(N__52454));
    Span4Mux_h I__12080 (
            .O(N__52457),
            .I(N__52451));
    Odrv12 I__12079 (
            .O(N__52454),
            .I(n15591));
    Odrv4 I__12078 (
            .O(N__52451),
            .I(n15591));
    InMux I__12077 (
            .O(N__52446),
            .I(n12576));
    CascadeMux I__12076 (
            .O(N__52443),
            .I(N__52440));
    InMux I__12075 (
            .O(N__52440),
            .I(N__52436));
    InMux I__12074 (
            .O(N__52439),
            .I(N__52433));
    LocalMux I__12073 (
            .O(N__52436),
            .I(N__52430));
    LocalMux I__12072 (
            .O(N__52433),
            .I(N__52427));
    Span4Mux_h I__12071 (
            .O(N__52430),
            .I(N__52424));
    Span4Mux_h I__12070 (
            .O(N__52427),
            .I(N__52421));
    Odrv4 I__12069 (
            .O(N__52424),
            .I(n1620_adj_600));
    Odrv4 I__12068 (
            .O(N__52421),
            .I(n1620_adj_600));
    InMux I__12067 (
            .O(N__52416),
            .I(N__52413));
    LocalMux I__12066 (
            .O(N__52413),
            .I(N__52410));
    Span4Mux_v I__12065 (
            .O(N__52410),
            .I(N__52405));
    InMux I__12064 (
            .O(N__52409),
            .I(N__52402));
    InMux I__12063 (
            .O(N__52408),
            .I(N__52399));
    Sp12to4 I__12062 (
            .O(N__52405),
            .I(N__52394));
    LocalMux I__12061 (
            .O(N__52402),
            .I(N__52394));
    LocalMux I__12060 (
            .O(N__52399),
            .I(encoder0_position_21));
    Odrv12 I__12059 (
            .O(N__52394),
            .I(encoder0_position_21));
    CascadeMux I__12058 (
            .O(N__52389),
            .I(N__52386));
    InMux I__12057 (
            .O(N__52386),
            .I(N__52383));
    LocalMux I__12056 (
            .O(N__52383),
            .I(N__52380));
    Span4Mux_v I__12055 (
            .O(N__52380),
            .I(N__52377));
    Span4Mux_h I__12054 (
            .O(N__52377),
            .I(N__52374));
    Odrv4 I__12053 (
            .O(N__52374),
            .I(n12_adj_630));
    CascadeMux I__12052 (
            .O(N__52371),
            .I(N__52368));
    InMux I__12051 (
            .O(N__52368),
            .I(N__52365));
    LocalMux I__12050 (
            .O(N__52365),
            .I(N__52362));
    Odrv12 I__12049 (
            .O(N__52362),
            .I(n1397));
    InMux I__12048 (
            .O(N__52359),
            .I(N__52356));
    LocalMux I__12047 (
            .O(N__52356),
            .I(N__52353));
    Span4Mux_h I__12046 (
            .O(N__52353),
            .I(N__52350));
    Span4Mux_h I__12045 (
            .O(N__52350),
            .I(N__52344));
    CascadeMux I__12044 (
            .O(N__52349),
            .I(N__52339));
    CascadeMux I__12043 (
            .O(N__52348),
            .I(N__52333));
    CascadeMux I__12042 (
            .O(N__52347),
            .I(N__52328));
    Span4Mux_v I__12041 (
            .O(N__52344),
            .I(N__52324));
    InMux I__12040 (
            .O(N__52343),
            .I(N__52319));
    InMux I__12039 (
            .O(N__52342),
            .I(N__52319));
    InMux I__12038 (
            .O(N__52339),
            .I(N__52314));
    InMux I__12037 (
            .O(N__52338),
            .I(N__52314));
    InMux I__12036 (
            .O(N__52337),
            .I(N__52311));
    InMux I__12035 (
            .O(N__52336),
            .I(N__52304));
    InMux I__12034 (
            .O(N__52333),
            .I(N__52304));
    InMux I__12033 (
            .O(N__52332),
            .I(N__52304));
    InMux I__12032 (
            .O(N__52331),
            .I(N__52301));
    InMux I__12031 (
            .O(N__52328),
            .I(N__52296));
    InMux I__12030 (
            .O(N__52327),
            .I(N__52296));
    Odrv4 I__12029 (
            .O(N__52324),
            .I(n1356));
    LocalMux I__12028 (
            .O(N__52319),
            .I(n1356));
    LocalMux I__12027 (
            .O(N__52314),
            .I(n1356));
    LocalMux I__12026 (
            .O(N__52311),
            .I(n1356));
    LocalMux I__12025 (
            .O(N__52304),
            .I(n1356));
    LocalMux I__12024 (
            .O(N__52301),
            .I(n1356));
    LocalMux I__12023 (
            .O(N__52296),
            .I(n1356));
    CascadeMux I__12022 (
            .O(N__52281),
            .I(N__52277));
    CascadeMux I__12021 (
            .O(N__52280),
            .I(N__52273));
    InMux I__12020 (
            .O(N__52277),
            .I(N__52270));
    InMux I__12019 (
            .O(N__52276),
            .I(N__52267));
    InMux I__12018 (
            .O(N__52273),
            .I(N__52264));
    LocalMux I__12017 (
            .O(N__52270),
            .I(N__52261));
    LocalMux I__12016 (
            .O(N__52267),
            .I(N__52258));
    LocalMux I__12015 (
            .O(N__52264),
            .I(N__52255));
    Odrv4 I__12014 (
            .O(N__52261),
            .I(n1429));
    Odrv4 I__12013 (
            .O(N__52258),
            .I(n1429));
    Odrv12 I__12012 (
            .O(N__52255),
            .I(n1429));
    InMux I__12011 (
            .O(N__52248),
            .I(N__52243));
    InMux I__12010 (
            .O(N__52247),
            .I(N__52240));
    InMux I__12009 (
            .O(N__52246),
            .I(N__52237));
    LocalMux I__12008 (
            .O(N__52243),
            .I(n298));
    LocalMux I__12007 (
            .O(N__52240),
            .I(n298));
    LocalMux I__12006 (
            .O(N__52237),
            .I(n298));
    InMux I__12005 (
            .O(N__52230),
            .I(N__52227));
    LocalMux I__12004 (
            .O(N__52227),
            .I(N__52224));
    Odrv4 I__12003 (
            .O(N__52224),
            .I(n1301));
    InMux I__12002 (
            .O(N__52221),
            .I(bfn_16_21_0_));
    CascadeMux I__12001 (
            .O(N__52218),
            .I(N__52215));
    InMux I__12000 (
            .O(N__52215),
            .I(N__52211));
    CascadeMux I__11999 (
            .O(N__52214),
            .I(N__52208));
    LocalMux I__11998 (
            .O(N__52211),
            .I(N__52205));
    InMux I__11997 (
            .O(N__52208),
            .I(N__52202));
    Span4Mux_h I__11996 (
            .O(N__52205),
            .I(N__52199));
    LocalMux I__11995 (
            .O(N__52202),
            .I(n1233));
    Odrv4 I__11994 (
            .O(N__52199),
            .I(n1233));
    InMux I__11993 (
            .O(N__52194),
            .I(N__52191));
    LocalMux I__11992 (
            .O(N__52191),
            .I(n1300));
    InMux I__11991 (
            .O(N__52188),
            .I(n12531));
    CascadeMux I__11990 (
            .O(N__52185),
            .I(N__52182));
    InMux I__11989 (
            .O(N__52182),
            .I(N__52179));
    LocalMux I__11988 (
            .O(N__52179),
            .I(N__52174));
    InMux I__11987 (
            .O(N__52178),
            .I(N__52171));
    InMux I__11986 (
            .O(N__52177),
            .I(N__52168));
    Span4Mux_h I__11985 (
            .O(N__52174),
            .I(N__52165));
    LocalMux I__11984 (
            .O(N__52171),
            .I(n1232));
    LocalMux I__11983 (
            .O(N__52168),
            .I(n1232));
    Odrv4 I__11982 (
            .O(N__52165),
            .I(n1232));
    InMux I__11981 (
            .O(N__52158),
            .I(N__52155));
    LocalMux I__11980 (
            .O(N__52155),
            .I(n1299));
    InMux I__11979 (
            .O(N__52152),
            .I(n12532));
    CascadeMux I__11978 (
            .O(N__52149),
            .I(N__52145));
    CascadeMux I__11977 (
            .O(N__52148),
            .I(N__52142));
    InMux I__11976 (
            .O(N__52145),
            .I(N__52138));
    InMux I__11975 (
            .O(N__52142),
            .I(N__52135));
    InMux I__11974 (
            .O(N__52141),
            .I(N__52132));
    LocalMux I__11973 (
            .O(N__52138),
            .I(n1530));
    LocalMux I__11972 (
            .O(N__52135),
            .I(n1530));
    LocalMux I__11971 (
            .O(N__52132),
            .I(n1530));
    InMux I__11970 (
            .O(N__52125),
            .I(N__52122));
    LocalMux I__11969 (
            .O(N__52122),
            .I(N__52119));
    Span4Mux_h I__11968 (
            .O(N__52119),
            .I(N__52116));
    Odrv4 I__11967 (
            .O(N__52116),
            .I(n1597));
    InMux I__11966 (
            .O(N__52113),
            .I(n12567));
    CascadeMux I__11965 (
            .O(N__52110),
            .I(N__52106));
    InMux I__11964 (
            .O(N__52109),
            .I(N__52102));
    InMux I__11963 (
            .O(N__52106),
            .I(N__52099));
    InMux I__11962 (
            .O(N__52105),
            .I(N__52096));
    LocalMux I__11961 (
            .O(N__52102),
            .I(n1529));
    LocalMux I__11960 (
            .O(N__52099),
            .I(n1529));
    LocalMux I__11959 (
            .O(N__52096),
            .I(n1529));
    InMux I__11958 (
            .O(N__52089),
            .I(N__52086));
    LocalMux I__11957 (
            .O(N__52086),
            .I(N__52083));
    Odrv4 I__11956 (
            .O(N__52083),
            .I(n1596));
    InMux I__11955 (
            .O(N__52080),
            .I(n12568));
    CascadeMux I__11954 (
            .O(N__52077),
            .I(N__52072));
    CascadeMux I__11953 (
            .O(N__52076),
            .I(N__52069));
    CascadeMux I__11952 (
            .O(N__52075),
            .I(N__52066));
    InMux I__11951 (
            .O(N__52072),
            .I(N__52063));
    InMux I__11950 (
            .O(N__52069),
            .I(N__52060));
    InMux I__11949 (
            .O(N__52066),
            .I(N__52057));
    LocalMux I__11948 (
            .O(N__52063),
            .I(n1528));
    LocalMux I__11947 (
            .O(N__52060),
            .I(n1528));
    LocalMux I__11946 (
            .O(N__52057),
            .I(n1528));
    InMux I__11945 (
            .O(N__52050),
            .I(N__52047));
    LocalMux I__11944 (
            .O(N__52047),
            .I(N__52044));
    Span4Mux_h I__11943 (
            .O(N__52044),
            .I(N__52041));
    Odrv4 I__11942 (
            .O(N__52041),
            .I(n1595));
    InMux I__11941 (
            .O(N__52038),
            .I(n12569));
    CascadeMux I__11940 (
            .O(N__52035),
            .I(N__52031));
    CascadeMux I__11939 (
            .O(N__52034),
            .I(N__52028));
    InMux I__11938 (
            .O(N__52031),
            .I(N__52024));
    InMux I__11937 (
            .O(N__52028),
            .I(N__52021));
    InMux I__11936 (
            .O(N__52027),
            .I(N__52018));
    LocalMux I__11935 (
            .O(N__52024),
            .I(n1527));
    LocalMux I__11934 (
            .O(N__52021),
            .I(n1527));
    LocalMux I__11933 (
            .O(N__52018),
            .I(n1527));
    InMux I__11932 (
            .O(N__52011),
            .I(N__52008));
    LocalMux I__11931 (
            .O(N__52008),
            .I(N__52005));
    Odrv12 I__11930 (
            .O(N__52005),
            .I(n1594));
    InMux I__11929 (
            .O(N__52002),
            .I(n12570));
    CascadeMux I__11928 (
            .O(N__51999),
            .I(N__51996));
    InMux I__11927 (
            .O(N__51996),
            .I(N__51993));
    LocalMux I__11926 (
            .O(N__51993),
            .I(N__51989));
    InMux I__11925 (
            .O(N__51992),
            .I(N__51986));
    Span4Mux_v I__11924 (
            .O(N__51989),
            .I(N__51982));
    LocalMux I__11923 (
            .O(N__51986),
            .I(N__51979));
    InMux I__11922 (
            .O(N__51985),
            .I(N__51976));
    Odrv4 I__11921 (
            .O(N__51982),
            .I(n1526));
    Odrv4 I__11920 (
            .O(N__51979),
            .I(n1526));
    LocalMux I__11919 (
            .O(N__51976),
            .I(n1526));
    InMux I__11918 (
            .O(N__51969),
            .I(N__51966));
    LocalMux I__11917 (
            .O(N__51966),
            .I(N__51963));
    Span4Mux_v I__11916 (
            .O(N__51963),
            .I(N__51960));
    Odrv4 I__11915 (
            .O(N__51960),
            .I(n1593));
    InMux I__11914 (
            .O(N__51957),
            .I(bfn_16_20_0_));
    CascadeMux I__11913 (
            .O(N__51954),
            .I(N__51950));
    CascadeMux I__11912 (
            .O(N__51953),
            .I(N__51947));
    InMux I__11911 (
            .O(N__51950),
            .I(N__51944));
    InMux I__11910 (
            .O(N__51947),
            .I(N__51940));
    LocalMux I__11909 (
            .O(N__51944),
            .I(N__51937));
    InMux I__11908 (
            .O(N__51943),
            .I(N__51934));
    LocalMux I__11907 (
            .O(N__51940),
            .I(n1525));
    Odrv4 I__11906 (
            .O(N__51937),
            .I(n1525));
    LocalMux I__11905 (
            .O(N__51934),
            .I(n1525));
    InMux I__11904 (
            .O(N__51927),
            .I(N__51924));
    LocalMux I__11903 (
            .O(N__51924),
            .I(N__51921));
    Span4Mux_h I__11902 (
            .O(N__51921),
            .I(N__51918));
    Odrv4 I__11901 (
            .O(N__51918),
            .I(n1592));
    InMux I__11900 (
            .O(N__51915),
            .I(n12572));
    CascadeMux I__11899 (
            .O(N__51912),
            .I(N__51909));
    InMux I__11898 (
            .O(N__51909),
            .I(N__51906));
    LocalMux I__11897 (
            .O(N__51906),
            .I(N__51901));
    InMux I__11896 (
            .O(N__51905),
            .I(N__51896));
    InMux I__11895 (
            .O(N__51904),
            .I(N__51896));
    Odrv4 I__11894 (
            .O(N__51901),
            .I(n1524));
    LocalMux I__11893 (
            .O(N__51896),
            .I(n1524));
    InMux I__11892 (
            .O(N__51891),
            .I(N__51888));
    LocalMux I__11891 (
            .O(N__51888),
            .I(N__51885));
    Span4Mux_h I__11890 (
            .O(N__51885),
            .I(N__51882));
    Odrv4 I__11889 (
            .O(N__51882),
            .I(n1591));
    InMux I__11888 (
            .O(N__51879),
            .I(n12573));
    CascadeMux I__11887 (
            .O(N__51876),
            .I(N__51873));
    InMux I__11886 (
            .O(N__51873),
            .I(N__51870));
    LocalMux I__11885 (
            .O(N__51870),
            .I(N__51867));
    Span4Mux_v I__11884 (
            .O(N__51867),
            .I(N__51863));
    InMux I__11883 (
            .O(N__51866),
            .I(N__51860));
    Odrv4 I__11882 (
            .O(N__51863),
            .I(n1523));
    LocalMux I__11881 (
            .O(N__51860),
            .I(n1523));
    InMux I__11880 (
            .O(N__51855),
            .I(N__51851));
    InMux I__11879 (
            .O(N__51854),
            .I(N__51848));
    LocalMux I__11878 (
            .O(N__51851),
            .I(n1425));
    LocalMux I__11877 (
            .O(N__51848),
            .I(n1425));
    InMux I__11876 (
            .O(N__51843),
            .I(N__51840));
    LocalMux I__11875 (
            .O(N__51840),
            .I(n1492));
    InMux I__11874 (
            .O(N__51837),
            .I(n12560));
    CascadeMux I__11873 (
            .O(N__51834),
            .I(N__51830));
    CascadeMux I__11872 (
            .O(N__51833),
            .I(N__51827));
    InMux I__11871 (
            .O(N__51830),
            .I(N__51824));
    InMux I__11870 (
            .O(N__51827),
            .I(N__51821));
    LocalMux I__11869 (
            .O(N__51824),
            .I(N__51816));
    LocalMux I__11868 (
            .O(N__51821),
            .I(N__51816));
    Span4Mux_h I__11867 (
            .O(N__51816),
            .I(N__51812));
    InMux I__11866 (
            .O(N__51815),
            .I(N__51809));
    Odrv4 I__11865 (
            .O(N__51812),
            .I(n1424));
    LocalMux I__11864 (
            .O(N__51809),
            .I(n1424));
    InMux I__11863 (
            .O(N__51804),
            .I(N__51801));
    LocalMux I__11862 (
            .O(N__51801),
            .I(N__51798));
    Odrv4 I__11861 (
            .O(N__51798),
            .I(n1491));
    InMux I__11860 (
            .O(N__51795),
            .I(n12561));
    CascadeMux I__11859 (
            .O(N__51792),
            .I(N__51788));
    InMux I__11858 (
            .O(N__51791),
            .I(N__51785));
    InMux I__11857 (
            .O(N__51788),
            .I(N__51782));
    LocalMux I__11856 (
            .O(N__51785),
            .I(N__51778));
    LocalMux I__11855 (
            .O(N__51782),
            .I(N__51775));
    InMux I__11854 (
            .O(N__51781),
            .I(N__51772));
    Odrv4 I__11853 (
            .O(N__51778),
            .I(n1423));
    Odrv4 I__11852 (
            .O(N__51775),
            .I(n1423));
    LocalMux I__11851 (
            .O(N__51772),
            .I(n1423));
    CascadeMux I__11850 (
            .O(N__51765),
            .I(N__51762));
    InMux I__11849 (
            .O(N__51762),
            .I(N__51759));
    LocalMux I__11848 (
            .O(N__51759),
            .I(n1490));
    InMux I__11847 (
            .O(N__51756),
            .I(n12562));
    InMux I__11846 (
            .O(N__51753),
            .I(N__51750));
    LocalMux I__11845 (
            .O(N__51750),
            .I(N__51747));
    Span12Mux_h I__11844 (
            .O(N__51747),
            .I(N__51743));
    InMux I__11843 (
            .O(N__51746),
            .I(N__51740));
    Odrv12 I__11842 (
            .O(N__51743),
            .I(n15572));
    LocalMux I__11841 (
            .O(N__51740),
            .I(n15572));
    CascadeMux I__11840 (
            .O(N__51735),
            .I(N__51732));
    InMux I__11839 (
            .O(N__51732),
            .I(N__51729));
    LocalMux I__11838 (
            .O(N__51729),
            .I(N__51725));
    InMux I__11837 (
            .O(N__51728),
            .I(N__51722));
    Span4Mux_h I__11836 (
            .O(N__51725),
            .I(N__51717));
    LocalMux I__11835 (
            .O(N__51722),
            .I(N__51717));
    Odrv4 I__11834 (
            .O(N__51717),
            .I(n1422));
    InMux I__11833 (
            .O(N__51714),
            .I(n12563));
    InMux I__11832 (
            .O(N__51711),
            .I(N__51707));
    InMux I__11831 (
            .O(N__51710),
            .I(N__51703));
    LocalMux I__11830 (
            .O(N__51707),
            .I(N__51700));
    InMux I__11829 (
            .O(N__51706),
            .I(N__51697));
    LocalMux I__11828 (
            .O(N__51703),
            .I(N__51694));
    Span4Mux_h I__11827 (
            .O(N__51700),
            .I(N__51689));
    LocalMux I__11826 (
            .O(N__51697),
            .I(N__51689));
    Span12Mux_v I__11825 (
            .O(N__51694),
            .I(N__51686));
    Span4Mux_h I__11824 (
            .O(N__51689),
            .I(N__51683));
    Odrv12 I__11823 (
            .O(N__51686),
            .I(n301));
    Odrv4 I__11822 (
            .O(N__51683),
            .I(n301));
    InMux I__11821 (
            .O(N__51678),
            .I(N__51675));
    LocalMux I__11820 (
            .O(N__51675),
            .I(N__51672));
    Span4Mux_h I__11819 (
            .O(N__51672),
            .I(N__51669));
    Odrv4 I__11818 (
            .O(N__51669),
            .I(n1601));
    InMux I__11817 (
            .O(N__51666),
            .I(bfn_16_19_0_));
    CascadeMux I__11816 (
            .O(N__51663),
            .I(N__51659));
    InMux I__11815 (
            .O(N__51662),
            .I(N__51655));
    InMux I__11814 (
            .O(N__51659),
            .I(N__51652));
    InMux I__11813 (
            .O(N__51658),
            .I(N__51649));
    LocalMux I__11812 (
            .O(N__51655),
            .I(n1533));
    LocalMux I__11811 (
            .O(N__51652),
            .I(n1533));
    LocalMux I__11810 (
            .O(N__51649),
            .I(n1533));
    CascadeMux I__11809 (
            .O(N__51642),
            .I(N__51639));
    InMux I__11808 (
            .O(N__51639),
            .I(N__51636));
    LocalMux I__11807 (
            .O(N__51636),
            .I(N__51633));
    Odrv4 I__11806 (
            .O(N__51633),
            .I(n1600));
    InMux I__11805 (
            .O(N__51630),
            .I(n12564));
    CascadeMux I__11804 (
            .O(N__51627),
            .I(N__51623));
    InMux I__11803 (
            .O(N__51626),
            .I(N__51619));
    InMux I__11802 (
            .O(N__51623),
            .I(N__51616));
    InMux I__11801 (
            .O(N__51622),
            .I(N__51613));
    LocalMux I__11800 (
            .O(N__51619),
            .I(n1532));
    LocalMux I__11799 (
            .O(N__51616),
            .I(n1532));
    LocalMux I__11798 (
            .O(N__51613),
            .I(n1532));
    InMux I__11797 (
            .O(N__51606),
            .I(N__51603));
    LocalMux I__11796 (
            .O(N__51603),
            .I(N__51600));
    Odrv4 I__11795 (
            .O(N__51600),
            .I(n1599));
    InMux I__11794 (
            .O(N__51597),
            .I(n12565));
    CascadeMux I__11793 (
            .O(N__51594),
            .I(N__51591));
    InMux I__11792 (
            .O(N__51591),
            .I(N__51587));
    CascadeMux I__11791 (
            .O(N__51590),
            .I(N__51584));
    LocalMux I__11790 (
            .O(N__51587),
            .I(N__51581));
    InMux I__11789 (
            .O(N__51584),
            .I(N__51578));
    Odrv4 I__11788 (
            .O(N__51581),
            .I(n1531));
    LocalMux I__11787 (
            .O(N__51578),
            .I(n1531));
    InMux I__11786 (
            .O(N__51573),
            .I(N__51570));
    LocalMux I__11785 (
            .O(N__51570),
            .I(N__51567));
    Span4Mux_v I__11784 (
            .O(N__51567),
            .I(N__51564));
    Odrv4 I__11783 (
            .O(N__51564),
            .I(n1598));
    InMux I__11782 (
            .O(N__51561),
            .I(n12566));
    CascadeMux I__11781 (
            .O(N__51558),
            .I(N__51554));
    CascadeMux I__11780 (
            .O(N__51557),
            .I(N__51551));
    InMux I__11779 (
            .O(N__51554),
            .I(N__51548));
    InMux I__11778 (
            .O(N__51551),
            .I(N__51545));
    LocalMux I__11777 (
            .O(N__51548),
            .I(N__51542));
    LocalMux I__11776 (
            .O(N__51545),
            .I(N__51539));
    Span4Mux_h I__11775 (
            .O(N__51542),
            .I(N__51535));
    Span4Mux_h I__11774 (
            .O(N__51539),
            .I(N__51532));
    InMux I__11773 (
            .O(N__51538),
            .I(N__51529));
    Span4Mux_v I__11772 (
            .O(N__51535),
            .I(N__51526));
    Odrv4 I__11771 (
            .O(N__51532),
            .I(n1433));
    LocalMux I__11770 (
            .O(N__51529),
            .I(n1433));
    Odrv4 I__11769 (
            .O(N__51526),
            .I(n1433));
    InMux I__11768 (
            .O(N__51519),
            .I(N__51516));
    LocalMux I__11767 (
            .O(N__51516),
            .I(n1500));
    InMux I__11766 (
            .O(N__51513),
            .I(n12552));
    CascadeMux I__11765 (
            .O(N__51510),
            .I(N__51507));
    InMux I__11764 (
            .O(N__51507),
            .I(N__51504));
    LocalMux I__11763 (
            .O(N__51504),
            .I(N__51500));
    InMux I__11762 (
            .O(N__51503),
            .I(N__51497));
    Span4Mux_v I__11761 (
            .O(N__51500),
            .I(N__51494));
    LocalMux I__11760 (
            .O(N__51497),
            .I(n1432));
    Odrv4 I__11759 (
            .O(N__51494),
            .I(n1432));
    InMux I__11758 (
            .O(N__51489),
            .I(N__51486));
    LocalMux I__11757 (
            .O(N__51486),
            .I(N__51483));
    Odrv4 I__11756 (
            .O(N__51483),
            .I(n1499));
    InMux I__11755 (
            .O(N__51480),
            .I(n12553));
    CascadeMux I__11754 (
            .O(N__51477),
            .I(N__51473));
    InMux I__11753 (
            .O(N__51476),
            .I(N__51470));
    InMux I__11752 (
            .O(N__51473),
            .I(N__51467));
    LocalMux I__11751 (
            .O(N__51470),
            .I(N__51461));
    LocalMux I__11750 (
            .O(N__51467),
            .I(N__51461));
    InMux I__11749 (
            .O(N__51466),
            .I(N__51458));
    Span4Mux_v I__11748 (
            .O(N__51461),
            .I(N__51455));
    LocalMux I__11747 (
            .O(N__51458),
            .I(n1431));
    Odrv4 I__11746 (
            .O(N__51455),
            .I(n1431));
    InMux I__11745 (
            .O(N__51450),
            .I(N__51447));
    LocalMux I__11744 (
            .O(N__51447),
            .I(n1498));
    InMux I__11743 (
            .O(N__51444),
            .I(n12554));
    CascadeMux I__11742 (
            .O(N__51441),
            .I(N__51437));
    CascadeMux I__11741 (
            .O(N__51440),
            .I(N__51434));
    InMux I__11740 (
            .O(N__51437),
            .I(N__51431));
    InMux I__11739 (
            .O(N__51434),
            .I(N__51428));
    LocalMux I__11738 (
            .O(N__51431),
            .I(N__51425));
    LocalMux I__11737 (
            .O(N__51428),
            .I(n1430));
    Odrv4 I__11736 (
            .O(N__51425),
            .I(n1430));
    InMux I__11735 (
            .O(N__51420),
            .I(N__51417));
    LocalMux I__11734 (
            .O(N__51417),
            .I(N__51414));
    Odrv4 I__11733 (
            .O(N__51414),
            .I(n1497));
    InMux I__11732 (
            .O(N__51411),
            .I(n12555));
    InMux I__11731 (
            .O(N__51408),
            .I(N__51405));
    LocalMux I__11730 (
            .O(N__51405),
            .I(n1496));
    InMux I__11729 (
            .O(N__51402),
            .I(n12556));
    CascadeMux I__11728 (
            .O(N__51399),
            .I(N__51396));
    InMux I__11727 (
            .O(N__51396),
            .I(N__51393));
    LocalMux I__11726 (
            .O(N__51393),
            .I(N__51389));
    InMux I__11725 (
            .O(N__51392),
            .I(N__51385));
    Span4Mux_h I__11724 (
            .O(N__51389),
            .I(N__51382));
    InMux I__11723 (
            .O(N__51388),
            .I(N__51379));
    LocalMux I__11722 (
            .O(N__51385),
            .I(n1428));
    Odrv4 I__11721 (
            .O(N__51382),
            .I(n1428));
    LocalMux I__11720 (
            .O(N__51379),
            .I(n1428));
    InMux I__11719 (
            .O(N__51372),
            .I(N__51369));
    LocalMux I__11718 (
            .O(N__51369),
            .I(n1495));
    InMux I__11717 (
            .O(N__51366),
            .I(n12557));
    CascadeMux I__11716 (
            .O(N__51363),
            .I(N__51360));
    InMux I__11715 (
            .O(N__51360),
            .I(N__51357));
    LocalMux I__11714 (
            .O(N__51357),
            .I(N__51353));
    InMux I__11713 (
            .O(N__51356),
            .I(N__51350));
    Span4Mux_h I__11712 (
            .O(N__51353),
            .I(N__51347));
    LocalMux I__11711 (
            .O(N__51350),
            .I(n1427));
    Odrv4 I__11710 (
            .O(N__51347),
            .I(n1427));
    InMux I__11709 (
            .O(N__51342),
            .I(N__51339));
    LocalMux I__11708 (
            .O(N__51339),
            .I(n1494));
    InMux I__11707 (
            .O(N__51336),
            .I(n12558));
    InMux I__11706 (
            .O(N__51333),
            .I(N__51329));
    CascadeMux I__11705 (
            .O(N__51332),
            .I(N__51326));
    LocalMux I__11704 (
            .O(N__51329),
            .I(N__51322));
    InMux I__11703 (
            .O(N__51326),
            .I(N__51319));
    InMux I__11702 (
            .O(N__51325),
            .I(N__51316));
    Odrv4 I__11701 (
            .O(N__51322),
            .I(n1426));
    LocalMux I__11700 (
            .O(N__51319),
            .I(n1426));
    LocalMux I__11699 (
            .O(N__51316),
            .I(n1426));
    InMux I__11698 (
            .O(N__51309),
            .I(N__51306));
    LocalMux I__11697 (
            .O(N__51306),
            .I(n1493));
    InMux I__11696 (
            .O(N__51303),
            .I(bfn_16_18_0_));
    CascadeMux I__11695 (
            .O(N__51300),
            .I(N__51297));
    InMux I__11694 (
            .O(N__51297),
            .I(N__51293));
    InMux I__11693 (
            .O(N__51296),
            .I(N__51288));
    LocalMux I__11692 (
            .O(N__51293),
            .I(N__51285));
    InMux I__11691 (
            .O(N__51292),
            .I(N__51280));
    InMux I__11690 (
            .O(N__51291),
            .I(N__51280));
    LocalMux I__11689 (
            .O(N__51288),
            .I(encoder0_position_target_20));
    Odrv4 I__11688 (
            .O(N__51285),
            .I(encoder0_position_target_20));
    LocalMux I__11687 (
            .O(N__51280),
            .I(encoder0_position_target_20));
    InMux I__11686 (
            .O(N__51273),
            .I(n12469));
    CascadeMux I__11685 (
            .O(N__51270),
            .I(N__51267));
    InMux I__11684 (
            .O(N__51267),
            .I(N__51261));
    InMux I__11683 (
            .O(N__51266),
            .I(N__51256));
    InMux I__11682 (
            .O(N__51265),
            .I(N__51256));
    CascadeMux I__11681 (
            .O(N__51264),
            .I(N__51253));
    LocalMux I__11680 (
            .O(N__51261),
            .I(N__51250));
    LocalMux I__11679 (
            .O(N__51256),
            .I(N__51247));
    InMux I__11678 (
            .O(N__51253),
            .I(N__51244));
    Span4Mux_h I__11677 (
            .O(N__51250),
            .I(N__51241));
    Span4Mux_h I__11676 (
            .O(N__51247),
            .I(N__51238));
    LocalMux I__11675 (
            .O(N__51244),
            .I(encoder0_position_target_21));
    Odrv4 I__11674 (
            .O(N__51241),
            .I(encoder0_position_target_21));
    Odrv4 I__11673 (
            .O(N__51238),
            .I(encoder0_position_target_21));
    InMux I__11672 (
            .O(N__51231),
            .I(n12470));
    CascadeMux I__11671 (
            .O(N__51228),
            .I(N__51224));
    InMux I__11670 (
            .O(N__51227),
            .I(N__51221));
    InMux I__11669 (
            .O(N__51224),
            .I(N__51217));
    LocalMux I__11668 (
            .O(N__51221),
            .I(N__51213));
    InMux I__11667 (
            .O(N__51220),
            .I(N__51210));
    LocalMux I__11666 (
            .O(N__51217),
            .I(N__51207));
    InMux I__11665 (
            .O(N__51216),
            .I(N__51204));
    Span4Mux_h I__11664 (
            .O(N__51213),
            .I(N__51201));
    LocalMux I__11663 (
            .O(N__51210),
            .I(encoder0_position_target_22));
    Odrv4 I__11662 (
            .O(N__51207),
            .I(encoder0_position_target_22));
    LocalMux I__11661 (
            .O(N__51204),
            .I(encoder0_position_target_22));
    Odrv4 I__11660 (
            .O(N__51201),
            .I(encoder0_position_target_22));
    InMux I__11659 (
            .O(N__51192),
            .I(n12471));
    CascadeMux I__11658 (
            .O(N__51189),
            .I(N__51182));
    CascadeMux I__11657 (
            .O(N__51188),
            .I(N__51178));
    CascadeMux I__11656 (
            .O(N__51187),
            .I(N__51174));
    CascadeMux I__11655 (
            .O(N__51186),
            .I(N__51170));
    InMux I__11654 (
            .O(N__51185),
            .I(N__51161));
    InMux I__11653 (
            .O(N__51182),
            .I(N__51144));
    InMux I__11652 (
            .O(N__51181),
            .I(N__51144));
    InMux I__11651 (
            .O(N__51178),
            .I(N__51144));
    InMux I__11650 (
            .O(N__51177),
            .I(N__51144));
    InMux I__11649 (
            .O(N__51174),
            .I(N__51144));
    InMux I__11648 (
            .O(N__51173),
            .I(N__51144));
    InMux I__11647 (
            .O(N__51170),
            .I(N__51144));
    InMux I__11646 (
            .O(N__51169),
            .I(N__51144));
    CascadeMux I__11645 (
            .O(N__51168),
            .I(N__51140));
    CascadeMux I__11644 (
            .O(N__51167),
            .I(N__51136));
    CascadeMux I__11643 (
            .O(N__51166),
            .I(N__51132));
    CascadeMux I__11642 (
            .O(N__51165),
            .I(N__51128));
    CascadeMux I__11641 (
            .O(N__51164),
            .I(N__51122));
    LocalMux I__11640 (
            .O(N__51161),
            .I(N__51110));
    LocalMux I__11639 (
            .O(N__51144),
            .I(N__51110));
    InMux I__11638 (
            .O(N__51143),
            .I(N__51093));
    InMux I__11637 (
            .O(N__51140),
            .I(N__51093));
    InMux I__11636 (
            .O(N__51139),
            .I(N__51093));
    InMux I__11635 (
            .O(N__51136),
            .I(N__51093));
    InMux I__11634 (
            .O(N__51135),
            .I(N__51093));
    InMux I__11633 (
            .O(N__51132),
            .I(N__51093));
    InMux I__11632 (
            .O(N__51131),
            .I(N__51093));
    InMux I__11631 (
            .O(N__51128),
            .I(N__51093));
    InMux I__11630 (
            .O(N__51127),
            .I(N__51084));
    InMux I__11629 (
            .O(N__51126),
            .I(N__51084));
    InMux I__11628 (
            .O(N__51125),
            .I(N__51084));
    InMux I__11627 (
            .O(N__51122),
            .I(N__51084));
    InMux I__11626 (
            .O(N__51121),
            .I(N__51075));
    InMux I__11625 (
            .O(N__51120),
            .I(N__51075));
    InMux I__11624 (
            .O(N__51119),
            .I(N__51075));
    InMux I__11623 (
            .O(N__51118),
            .I(N__51075));
    InMux I__11622 (
            .O(N__51117),
            .I(N__51068));
    InMux I__11621 (
            .O(N__51116),
            .I(N__51068));
    InMux I__11620 (
            .O(N__51115),
            .I(N__51068));
    Odrv4 I__11619 (
            .O(N__51110),
            .I(direction_c));
    LocalMux I__11618 (
            .O(N__51093),
            .I(direction_c));
    LocalMux I__11617 (
            .O(N__51084),
            .I(direction_c));
    LocalMux I__11616 (
            .O(N__51075),
            .I(direction_c));
    LocalMux I__11615 (
            .O(N__51068),
            .I(direction_c));
    InMux I__11614 (
            .O(N__51057),
            .I(bfn_15_28_0_));
    InMux I__11613 (
            .O(N__51054),
            .I(N__51051));
    LocalMux I__11612 (
            .O(N__51051),
            .I(N__51046));
    InMux I__11611 (
            .O(N__51050),
            .I(N__51043));
    CascadeMux I__11610 (
            .O(N__51049),
            .I(N__51040));
    Span4Mux_v I__11609 (
            .O(N__51046),
            .I(N__51034));
    LocalMux I__11608 (
            .O(N__51043),
            .I(N__51031));
    InMux I__11607 (
            .O(N__51040),
            .I(N__51028));
    InMux I__11606 (
            .O(N__51039),
            .I(N__51025));
    InMux I__11605 (
            .O(N__51038),
            .I(N__51022));
    InMux I__11604 (
            .O(N__51037),
            .I(N__51019));
    Span4Mux_h I__11603 (
            .O(N__51034),
            .I(N__51016));
    Span4Mux_h I__11602 (
            .O(N__51031),
            .I(N__51013));
    LocalMux I__11601 (
            .O(N__51028),
            .I(N__51006));
    LocalMux I__11600 (
            .O(N__51025),
            .I(N__51006));
    LocalMux I__11599 (
            .O(N__51022),
            .I(N__51006));
    LocalMux I__11598 (
            .O(N__51019),
            .I(encoder0_position_target_23));
    Odrv4 I__11597 (
            .O(N__51016),
            .I(encoder0_position_target_23));
    Odrv4 I__11596 (
            .O(N__51013),
            .I(encoder0_position_target_23));
    Odrv4 I__11595 (
            .O(N__51006),
            .I(encoder0_position_target_23));
    InMux I__11594 (
            .O(N__50997),
            .I(N__50994));
    LocalMux I__11593 (
            .O(N__50994),
            .I(N__50991));
    Span4Mux_h I__11592 (
            .O(N__50991),
            .I(N__50988));
    Span4Mux_h I__11591 (
            .O(N__50988),
            .I(N__50985));
    Odrv4 I__11590 (
            .O(N__50985),
            .I(pwm_setpoint_23));
    InMux I__11589 (
            .O(N__50982),
            .I(N__50977));
    InMux I__11588 (
            .O(N__50981),
            .I(N__50974));
    InMux I__11587 (
            .O(N__50980),
            .I(N__50971));
    LocalMux I__11586 (
            .O(N__50977),
            .I(pwm_counter_23));
    LocalMux I__11585 (
            .O(N__50974),
            .I(pwm_counter_23));
    LocalMux I__11584 (
            .O(N__50971),
            .I(pwm_counter_23));
    InMux I__11583 (
            .O(N__50964),
            .I(N__50961));
    LocalMux I__11582 (
            .O(N__50961),
            .I(N__50958));
    Span4Mux_h I__11581 (
            .O(N__50958),
            .I(N__50955));
    Odrv4 I__11580 (
            .O(N__50955),
            .I(n15245));
    InMux I__11579 (
            .O(N__50952),
            .I(N__50947));
    InMux I__11578 (
            .O(N__50951),
            .I(N__50944));
    InMux I__11577 (
            .O(N__50950),
            .I(N__50941));
    LocalMux I__11576 (
            .O(N__50947),
            .I(pwm_counter_31));
    LocalMux I__11575 (
            .O(N__50944),
            .I(pwm_counter_31));
    LocalMux I__11574 (
            .O(N__50941),
            .I(pwm_counter_31));
    InMux I__11573 (
            .O(N__50934),
            .I(N__50930));
    InMux I__11572 (
            .O(N__50933),
            .I(N__50927));
    LocalMux I__11571 (
            .O(N__50930),
            .I(N__50924));
    LocalMux I__11570 (
            .O(N__50927),
            .I(n5180));
    Odrv4 I__11569 (
            .O(N__50924),
            .I(n5180));
    SRMux I__11568 (
            .O(N__50919),
            .I(N__50916));
    LocalMux I__11567 (
            .O(N__50916),
            .I(N__50913));
    Odrv12 I__11566 (
            .O(N__50913),
            .I(n5182));
    InMux I__11565 (
            .O(N__50910),
            .I(N__50902));
    InMux I__11564 (
            .O(N__50909),
            .I(N__50896));
    InMux I__11563 (
            .O(N__50908),
            .I(N__50885));
    InMux I__11562 (
            .O(N__50907),
            .I(N__50885));
    InMux I__11561 (
            .O(N__50906),
            .I(N__50885));
    InMux I__11560 (
            .O(N__50905),
            .I(N__50882));
    LocalMux I__11559 (
            .O(N__50902),
            .I(N__50879));
    InMux I__11558 (
            .O(N__50901),
            .I(N__50874));
    InMux I__11557 (
            .O(N__50900),
            .I(N__50874));
    InMux I__11556 (
            .O(N__50899),
            .I(N__50870));
    LocalMux I__11555 (
            .O(N__50896),
            .I(N__50864));
    InMux I__11554 (
            .O(N__50895),
            .I(N__50858));
    InMux I__11553 (
            .O(N__50894),
            .I(N__50858));
    InMux I__11552 (
            .O(N__50893),
            .I(N__50853));
    InMux I__11551 (
            .O(N__50892),
            .I(N__50853));
    LocalMux I__11550 (
            .O(N__50885),
            .I(N__50850));
    LocalMux I__11549 (
            .O(N__50882),
            .I(N__50847));
    Span4Mux_s1_v I__11548 (
            .O(N__50879),
            .I(N__50842));
    LocalMux I__11547 (
            .O(N__50874),
            .I(N__50842));
    InMux I__11546 (
            .O(N__50873),
            .I(N__50839));
    LocalMux I__11545 (
            .O(N__50870),
            .I(N__50829));
    InMux I__11544 (
            .O(N__50869),
            .I(N__50822));
    InMux I__11543 (
            .O(N__50868),
            .I(N__50822));
    InMux I__11542 (
            .O(N__50867),
            .I(N__50822));
    Span4Mux_v I__11541 (
            .O(N__50864),
            .I(N__50819));
    InMux I__11540 (
            .O(N__50863),
            .I(N__50816));
    LocalMux I__11539 (
            .O(N__50858),
            .I(N__50811));
    LocalMux I__11538 (
            .O(N__50853),
            .I(N__50811));
    Span4Mux_v I__11537 (
            .O(N__50850),
            .I(N__50806));
    Span4Mux_v I__11536 (
            .O(N__50847),
            .I(N__50806));
    Sp12to4 I__11535 (
            .O(N__50842),
            .I(N__50801));
    LocalMux I__11534 (
            .O(N__50839),
            .I(N__50801));
    InMux I__11533 (
            .O(N__50838),
            .I(N__50798));
    InMux I__11532 (
            .O(N__50837),
            .I(N__50795));
    InMux I__11531 (
            .O(N__50836),
            .I(N__50792));
    InMux I__11530 (
            .O(N__50835),
            .I(N__50789));
    InMux I__11529 (
            .O(N__50834),
            .I(N__50782));
    InMux I__11528 (
            .O(N__50833),
            .I(N__50782));
    InMux I__11527 (
            .O(N__50832),
            .I(N__50782));
    Span12Mux_s5_v I__11526 (
            .O(N__50829),
            .I(N__50773));
    LocalMux I__11525 (
            .O(N__50822),
            .I(N__50773));
    Sp12to4 I__11524 (
            .O(N__50819),
            .I(N__50773));
    LocalMux I__11523 (
            .O(N__50816),
            .I(N__50773));
    Odrv4 I__11522 (
            .O(N__50811),
            .I(duty_23));
    Odrv4 I__11521 (
            .O(N__50806),
            .I(duty_23));
    Odrv12 I__11520 (
            .O(N__50801),
            .I(duty_23));
    LocalMux I__11519 (
            .O(N__50798),
            .I(duty_23));
    LocalMux I__11518 (
            .O(N__50795),
            .I(duty_23));
    LocalMux I__11517 (
            .O(N__50792),
            .I(duty_23));
    LocalMux I__11516 (
            .O(N__50789),
            .I(duty_23));
    LocalMux I__11515 (
            .O(N__50782),
            .I(duty_23));
    Odrv12 I__11514 (
            .O(N__50773),
            .I(duty_23));
    InMux I__11513 (
            .O(N__50754),
            .I(N__50751));
    LocalMux I__11512 (
            .O(N__50751),
            .I(N__50747));
    InMux I__11511 (
            .O(N__50750),
            .I(N__50744));
    Span4Mux_h I__11510 (
            .O(N__50747),
            .I(N__50740));
    LocalMux I__11509 (
            .O(N__50744),
            .I(N__50737));
    InMux I__11508 (
            .O(N__50743),
            .I(N__50734));
    Span4Mux_h I__11507 (
            .O(N__50740),
            .I(N__50731));
    Span12Mux_h I__11506 (
            .O(N__50737),
            .I(N__50728));
    LocalMux I__11505 (
            .O(N__50734),
            .I(N__50725));
    Odrv4 I__11504 (
            .O(N__50731),
            .I(n300));
    Odrv12 I__11503 (
            .O(N__50728),
            .I(n300));
    Odrv12 I__11502 (
            .O(N__50725),
            .I(n300));
    InMux I__11501 (
            .O(N__50718),
            .I(N__50715));
    LocalMux I__11500 (
            .O(N__50715),
            .I(n1501));
    InMux I__11499 (
            .O(N__50712),
            .I(bfn_16_17_0_));
    CascadeMux I__11498 (
            .O(N__50709),
            .I(N__50706));
    InMux I__11497 (
            .O(N__50706),
            .I(N__50701));
    CascadeMux I__11496 (
            .O(N__50705),
            .I(N__50697));
    InMux I__11495 (
            .O(N__50704),
            .I(N__50694));
    LocalMux I__11494 (
            .O(N__50701),
            .I(N__50691));
    InMux I__11493 (
            .O(N__50700),
            .I(N__50686));
    InMux I__11492 (
            .O(N__50697),
            .I(N__50686));
    LocalMux I__11491 (
            .O(N__50694),
            .I(encoder0_position_target_11));
    Odrv4 I__11490 (
            .O(N__50691),
            .I(encoder0_position_target_11));
    LocalMux I__11489 (
            .O(N__50686),
            .I(encoder0_position_target_11));
    InMux I__11488 (
            .O(N__50679),
            .I(n12460));
    CascadeMux I__11487 (
            .O(N__50676),
            .I(N__50671));
    CascadeMux I__11486 (
            .O(N__50675),
            .I(N__50667));
    InMux I__11485 (
            .O(N__50674),
            .I(N__50664));
    InMux I__11484 (
            .O(N__50671),
            .I(N__50661));
    InMux I__11483 (
            .O(N__50670),
            .I(N__50658));
    InMux I__11482 (
            .O(N__50667),
            .I(N__50655));
    LocalMux I__11481 (
            .O(N__50664),
            .I(N__50652));
    LocalMux I__11480 (
            .O(N__50661),
            .I(N__50647));
    LocalMux I__11479 (
            .O(N__50658),
            .I(N__50647));
    LocalMux I__11478 (
            .O(N__50655),
            .I(encoder0_position_target_12));
    Odrv4 I__11477 (
            .O(N__50652),
            .I(encoder0_position_target_12));
    Odrv4 I__11476 (
            .O(N__50647),
            .I(encoder0_position_target_12));
    InMux I__11475 (
            .O(N__50640),
            .I(n12461));
    CascadeMux I__11474 (
            .O(N__50637),
            .I(N__50634));
    InMux I__11473 (
            .O(N__50634),
            .I(N__50631));
    LocalMux I__11472 (
            .O(N__50631),
            .I(N__50626));
    InMux I__11471 (
            .O(N__50630),
            .I(N__50622));
    InMux I__11470 (
            .O(N__50629),
            .I(N__50619));
    Span4Mux_h I__11469 (
            .O(N__50626),
            .I(N__50616));
    InMux I__11468 (
            .O(N__50625),
            .I(N__50613));
    LocalMux I__11467 (
            .O(N__50622),
            .I(N__50610));
    LocalMux I__11466 (
            .O(N__50619),
            .I(encoder0_position_target_13));
    Odrv4 I__11465 (
            .O(N__50616),
            .I(encoder0_position_target_13));
    LocalMux I__11464 (
            .O(N__50613),
            .I(encoder0_position_target_13));
    Odrv12 I__11463 (
            .O(N__50610),
            .I(encoder0_position_target_13));
    InMux I__11462 (
            .O(N__50601),
            .I(n12462));
    CascadeMux I__11461 (
            .O(N__50598),
            .I(N__50594));
    CascadeMux I__11460 (
            .O(N__50597),
            .I(N__50591));
    InMux I__11459 (
            .O(N__50594),
            .I(N__50588));
    InMux I__11458 (
            .O(N__50591),
            .I(N__50583));
    LocalMux I__11457 (
            .O(N__50588),
            .I(N__50580));
    InMux I__11456 (
            .O(N__50587),
            .I(N__50575));
    InMux I__11455 (
            .O(N__50586),
            .I(N__50575));
    LocalMux I__11454 (
            .O(N__50583),
            .I(encoder0_position_target_14));
    Odrv12 I__11453 (
            .O(N__50580),
            .I(encoder0_position_target_14));
    LocalMux I__11452 (
            .O(N__50575),
            .I(encoder0_position_target_14));
    InMux I__11451 (
            .O(N__50568),
            .I(n12463));
    CascadeMux I__11450 (
            .O(N__50565),
            .I(N__50562));
    InMux I__11449 (
            .O(N__50562),
            .I(N__50559));
    LocalMux I__11448 (
            .O(N__50559),
            .I(N__50554));
    CascadeMux I__11447 (
            .O(N__50558),
            .I(N__50551));
    InMux I__11446 (
            .O(N__50557),
            .I(N__50548));
    Span4Mux_v I__11445 (
            .O(N__50554),
            .I(N__50545));
    InMux I__11444 (
            .O(N__50551),
            .I(N__50541));
    LocalMux I__11443 (
            .O(N__50548),
            .I(N__50538));
    Span4Mux_h I__11442 (
            .O(N__50545),
            .I(N__50535));
    InMux I__11441 (
            .O(N__50544),
            .I(N__50532));
    LocalMux I__11440 (
            .O(N__50541),
            .I(N__50527));
    Span4Mux_v I__11439 (
            .O(N__50538),
            .I(N__50527));
    Odrv4 I__11438 (
            .O(N__50535),
            .I(encoder0_position_target_15));
    LocalMux I__11437 (
            .O(N__50532),
            .I(encoder0_position_target_15));
    Odrv4 I__11436 (
            .O(N__50527),
            .I(encoder0_position_target_15));
    InMux I__11435 (
            .O(N__50520),
            .I(bfn_15_27_0_));
    CascadeMux I__11434 (
            .O(N__50517),
            .I(N__50514));
    InMux I__11433 (
            .O(N__50514),
            .I(N__50511));
    LocalMux I__11432 (
            .O(N__50511),
            .I(N__50506));
    CascadeMux I__11431 (
            .O(N__50510),
            .I(N__50502));
    InMux I__11430 (
            .O(N__50509),
            .I(N__50499));
    Span4Mux_h I__11429 (
            .O(N__50506),
            .I(N__50496));
    InMux I__11428 (
            .O(N__50505),
            .I(N__50491));
    InMux I__11427 (
            .O(N__50502),
            .I(N__50491));
    LocalMux I__11426 (
            .O(N__50499),
            .I(encoder0_position_target_16));
    Odrv4 I__11425 (
            .O(N__50496),
            .I(encoder0_position_target_16));
    LocalMux I__11424 (
            .O(N__50491),
            .I(encoder0_position_target_16));
    InMux I__11423 (
            .O(N__50484),
            .I(n12465));
    CascadeMux I__11422 (
            .O(N__50481),
            .I(N__50478));
    InMux I__11421 (
            .O(N__50478),
            .I(N__50473));
    CascadeMux I__11420 (
            .O(N__50477),
            .I(N__50470));
    InMux I__11419 (
            .O(N__50476),
            .I(N__50467));
    LocalMux I__11418 (
            .O(N__50473),
            .I(N__50464));
    InMux I__11417 (
            .O(N__50470),
            .I(N__50460));
    LocalMux I__11416 (
            .O(N__50467),
            .I(N__50457));
    Span4Mux_h I__11415 (
            .O(N__50464),
            .I(N__50454));
    InMux I__11414 (
            .O(N__50463),
            .I(N__50451));
    LocalMux I__11413 (
            .O(N__50460),
            .I(N__50446));
    Span4Mux_v I__11412 (
            .O(N__50457),
            .I(N__50446));
    Odrv4 I__11411 (
            .O(N__50454),
            .I(encoder0_position_target_17));
    LocalMux I__11410 (
            .O(N__50451),
            .I(encoder0_position_target_17));
    Odrv4 I__11409 (
            .O(N__50446),
            .I(encoder0_position_target_17));
    InMux I__11408 (
            .O(N__50439),
            .I(n12466));
    CascadeMux I__11407 (
            .O(N__50436),
            .I(N__50433));
    InMux I__11406 (
            .O(N__50433),
            .I(N__50430));
    LocalMux I__11405 (
            .O(N__50430),
            .I(N__50426));
    InMux I__11404 (
            .O(N__50429),
            .I(N__50423));
    Span4Mux_h I__11403 (
            .O(N__50426),
            .I(N__50420));
    LocalMux I__11402 (
            .O(N__50423),
            .I(N__50413));
    Span4Mux_v I__11401 (
            .O(N__50420),
            .I(N__50413));
    InMux I__11400 (
            .O(N__50419),
            .I(N__50410));
    InMux I__11399 (
            .O(N__50418),
            .I(N__50407));
    Odrv4 I__11398 (
            .O(N__50413),
            .I(encoder0_position_target_18));
    LocalMux I__11397 (
            .O(N__50410),
            .I(encoder0_position_target_18));
    LocalMux I__11396 (
            .O(N__50407),
            .I(encoder0_position_target_18));
    InMux I__11395 (
            .O(N__50400),
            .I(n12467));
    CascadeMux I__11394 (
            .O(N__50397),
            .I(N__50393));
    CascadeMux I__11393 (
            .O(N__50396),
            .I(N__50388));
    InMux I__11392 (
            .O(N__50393),
            .I(N__50385));
    InMux I__11391 (
            .O(N__50392),
            .I(N__50382));
    CascadeMux I__11390 (
            .O(N__50391),
            .I(N__50379));
    InMux I__11389 (
            .O(N__50388),
            .I(N__50376));
    LocalMux I__11388 (
            .O(N__50385),
            .I(N__50371));
    LocalMux I__11387 (
            .O(N__50382),
            .I(N__50371));
    InMux I__11386 (
            .O(N__50379),
            .I(N__50368));
    LocalMux I__11385 (
            .O(N__50376),
            .I(N__50365));
    Span4Mux_h I__11384 (
            .O(N__50371),
            .I(N__50362));
    LocalMux I__11383 (
            .O(N__50368),
            .I(encoder0_position_target_19));
    Odrv4 I__11382 (
            .O(N__50365),
            .I(encoder0_position_target_19));
    Odrv4 I__11381 (
            .O(N__50362),
            .I(encoder0_position_target_19));
    InMux I__11380 (
            .O(N__50355),
            .I(n12468));
    CascadeMux I__11379 (
            .O(N__50352),
            .I(N__50348));
    CascadeMux I__11378 (
            .O(N__50351),
            .I(N__50344));
    InMux I__11377 (
            .O(N__50348),
            .I(N__50341));
    InMux I__11376 (
            .O(N__50347),
            .I(N__50338));
    InMux I__11375 (
            .O(N__50344),
            .I(N__50335));
    LocalMux I__11374 (
            .O(N__50341),
            .I(N__50332));
    LocalMux I__11373 (
            .O(N__50338),
            .I(N__50329));
    LocalMux I__11372 (
            .O(N__50335),
            .I(encoder0_position_target_3));
    Odrv4 I__11371 (
            .O(N__50332),
            .I(encoder0_position_target_3));
    Odrv4 I__11370 (
            .O(N__50329),
            .I(encoder0_position_target_3));
    InMux I__11369 (
            .O(N__50322),
            .I(n12452));
    CascadeMux I__11368 (
            .O(N__50319),
            .I(N__50314));
    InMux I__11367 (
            .O(N__50318),
            .I(N__50311));
    CascadeMux I__11366 (
            .O(N__50317),
            .I(N__50307));
    InMux I__11365 (
            .O(N__50314),
            .I(N__50304));
    LocalMux I__11364 (
            .O(N__50311),
            .I(N__50301));
    InMux I__11363 (
            .O(N__50310),
            .I(N__50298));
    InMux I__11362 (
            .O(N__50307),
            .I(N__50295));
    LocalMux I__11361 (
            .O(N__50304),
            .I(N__50292));
    Span4Mux_h I__11360 (
            .O(N__50301),
            .I(N__50289));
    LocalMux I__11359 (
            .O(N__50298),
            .I(N__50286));
    LocalMux I__11358 (
            .O(N__50295),
            .I(encoder0_position_target_4));
    Odrv12 I__11357 (
            .O(N__50292),
            .I(encoder0_position_target_4));
    Odrv4 I__11356 (
            .O(N__50289),
            .I(encoder0_position_target_4));
    Odrv4 I__11355 (
            .O(N__50286),
            .I(encoder0_position_target_4));
    InMux I__11354 (
            .O(N__50277),
            .I(n12453));
    CascadeMux I__11353 (
            .O(N__50274),
            .I(N__50271));
    InMux I__11352 (
            .O(N__50271),
            .I(N__50267));
    CascadeMux I__11351 (
            .O(N__50270),
            .I(N__50262));
    LocalMux I__11350 (
            .O(N__50267),
            .I(N__50259));
    InMux I__11349 (
            .O(N__50266),
            .I(N__50254));
    InMux I__11348 (
            .O(N__50265),
            .I(N__50254));
    InMux I__11347 (
            .O(N__50262),
            .I(N__50251));
    Span4Mux_h I__11346 (
            .O(N__50259),
            .I(N__50246));
    LocalMux I__11345 (
            .O(N__50254),
            .I(N__50246));
    LocalMux I__11344 (
            .O(N__50251),
            .I(encoder0_position_target_5));
    Odrv4 I__11343 (
            .O(N__50246),
            .I(encoder0_position_target_5));
    InMux I__11342 (
            .O(N__50241),
            .I(n12454));
    CascadeMux I__11341 (
            .O(N__50238),
            .I(N__50234));
    CascadeMux I__11340 (
            .O(N__50237),
            .I(N__50229));
    InMux I__11339 (
            .O(N__50234),
            .I(N__50226));
    InMux I__11338 (
            .O(N__50233),
            .I(N__50221));
    InMux I__11337 (
            .O(N__50232),
            .I(N__50221));
    InMux I__11336 (
            .O(N__50229),
            .I(N__50218));
    LocalMux I__11335 (
            .O(N__50226),
            .I(N__50215));
    LocalMux I__11334 (
            .O(N__50221),
            .I(N__50212));
    LocalMux I__11333 (
            .O(N__50218),
            .I(encoder0_position_target_6));
    Odrv4 I__11332 (
            .O(N__50215),
            .I(encoder0_position_target_6));
    Odrv4 I__11331 (
            .O(N__50212),
            .I(encoder0_position_target_6));
    InMux I__11330 (
            .O(N__50205),
            .I(n12455));
    CascadeMux I__11329 (
            .O(N__50202),
            .I(N__50199));
    InMux I__11328 (
            .O(N__50199),
            .I(N__50195));
    CascadeMux I__11327 (
            .O(N__50198),
            .I(N__50192));
    LocalMux I__11326 (
            .O(N__50195),
            .I(N__50188));
    InMux I__11325 (
            .O(N__50192),
            .I(N__50185));
    InMux I__11324 (
            .O(N__50191),
            .I(N__50182));
    Span4Mux_v I__11323 (
            .O(N__50188),
            .I(N__50178));
    LocalMux I__11322 (
            .O(N__50185),
            .I(N__50173));
    LocalMux I__11321 (
            .O(N__50182),
            .I(N__50173));
    InMux I__11320 (
            .O(N__50181),
            .I(N__50170));
    Span4Mux_v I__11319 (
            .O(N__50178),
            .I(N__50165));
    Span4Mux_v I__11318 (
            .O(N__50173),
            .I(N__50165));
    LocalMux I__11317 (
            .O(N__50170),
            .I(encoder0_position_target_7));
    Odrv4 I__11316 (
            .O(N__50165),
            .I(encoder0_position_target_7));
    InMux I__11315 (
            .O(N__50160),
            .I(bfn_15_26_0_));
    CascadeMux I__11314 (
            .O(N__50157),
            .I(N__50154));
    InMux I__11313 (
            .O(N__50154),
            .I(N__50148));
    InMux I__11312 (
            .O(N__50153),
            .I(N__50145));
    CascadeMux I__11311 (
            .O(N__50152),
            .I(N__50142));
    InMux I__11310 (
            .O(N__50151),
            .I(N__50139));
    LocalMux I__11309 (
            .O(N__50148),
            .I(N__50134));
    LocalMux I__11308 (
            .O(N__50145),
            .I(N__50134));
    InMux I__11307 (
            .O(N__50142),
            .I(N__50131));
    LocalMux I__11306 (
            .O(N__50139),
            .I(N__50126));
    Span4Mux_v I__11305 (
            .O(N__50134),
            .I(N__50126));
    LocalMux I__11304 (
            .O(N__50131),
            .I(encoder0_position_target_8));
    Odrv4 I__11303 (
            .O(N__50126),
            .I(encoder0_position_target_8));
    InMux I__11302 (
            .O(N__50121),
            .I(n12457));
    CascadeMux I__11301 (
            .O(N__50118),
            .I(N__50114));
    InMux I__11300 (
            .O(N__50117),
            .I(N__50111));
    InMux I__11299 (
            .O(N__50114),
            .I(N__50108));
    LocalMux I__11298 (
            .O(N__50111),
            .I(N__50103));
    LocalMux I__11297 (
            .O(N__50108),
            .I(N__50100));
    InMux I__11296 (
            .O(N__50107),
            .I(N__50097));
    InMux I__11295 (
            .O(N__50106),
            .I(N__50094));
    Span4Mux_h I__11294 (
            .O(N__50103),
            .I(N__50091));
    Span4Mux_v I__11293 (
            .O(N__50100),
            .I(N__50086));
    LocalMux I__11292 (
            .O(N__50097),
            .I(N__50086));
    LocalMux I__11291 (
            .O(N__50094),
            .I(encoder0_position_target_9));
    Odrv4 I__11290 (
            .O(N__50091),
            .I(encoder0_position_target_9));
    Odrv4 I__11289 (
            .O(N__50086),
            .I(encoder0_position_target_9));
    InMux I__11288 (
            .O(N__50079),
            .I(n12458));
    CascadeMux I__11287 (
            .O(N__50076),
            .I(N__50073));
    InMux I__11286 (
            .O(N__50073),
            .I(N__50067));
    InMux I__11285 (
            .O(N__50072),
            .I(N__50062));
    InMux I__11284 (
            .O(N__50071),
            .I(N__50062));
    CascadeMux I__11283 (
            .O(N__50070),
            .I(N__50059));
    LocalMux I__11282 (
            .O(N__50067),
            .I(N__50056));
    LocalMux I__11281 (
            .O(N__50062),
            .I(N__50053));
    InMux I__11280 (
            .O(N__50059),
            .I(N__50050));
    Span4Mux_h I__11279 (
            .O(N__50056),
            .I(N__50047));
    Span4Mux_h I__11278 (
            .O(N__50053),
            .I(N__50044));
    LocalMux I__11277 (
            .O(N__50050),
            .I(encoder0_position_target_10));
    Odrv4 I__11276 (
            .O(N__50047),
            .I(encoder0_position_target_10));
    Odrv4 I__11275 (
            .O(N__50044),
            .I(encoder0_position_target_10));
    InMux I__11274 (
            .O(N__50037),
            .I(n12459));
    InMux I__11273 (
            .O(N__50034),
            .I(N__50030));
    CascadeMux I__11272 (
            .O(N__50033),
            .I(N__50027));
    LocalMux I__11271 (
            .O(N__50030),
            .I(N__50023));
    InMux I__11270 (
            .O(N__50027),
            .I(N__50020));
    InMux I__11269 (
            .O(N__50026),
            .I(N__50017));
    Odrv12 I__11268 (
            .O(N__50023),
            .I(n1126));
    LocalMux I__11267 (
            .O(N__50020),
            .I(n1126));
    LocalMux I__11266 (
            .O(N__50017),
            .I(n1126));
    InMux I__11265 (
            .O(N__50010),
            .I(N__50007));
    LocalMux I__11264 (
            .O(N__50007),
            .I(n1193));
    CascadeMux I__11263 (
            .O(N__50004),
            .I(n1225_cascade_));
    InMux I__11262 (
            .O(N__50001),
            .I(N__49996));
    InMux I__11261 (
            .O(N__50000),
            .I(N__49991));
    InMux I__11260 (
            .O(N__49999),
            .I(N__49991));
    LocalMux I__11259 (
            .O(N__49996),
            .I(N__49986));
    LocalMux I__11258 (
            .O(N__49991),
            .I(N__49986));
    Odrv4 I__11257 (
            .O(N__49986),
            .I(n1324));
    InMux I__11256 (
            .O(N__49983),
            .I(N__49980));
    LocalMux I__11255 (
            .O(N__49980),
            .I(N__49976));
    CascadeMux I__11254 (
            .O(N__49979),
            .I(N__49973));
    Span4Mux_v I__11253 (
            .O(N__49976),
            .I(N__49970));
    InMux I__11252 (
            .O(N__49973),
            .I(N__49967));
    Odrv4 I__11251 (
            .O(N__49970),
            .I(n1129));
    LocalMux I__11250 (
            .O(N__49967),
            .I(n1129));
    CascadeMux I__11249 (
            .O(N__49962),
            .I(N__49959));
    InMux I__11248 (
            .O(N__49959),
            .I(N__49956));
    LocalMux I__11247 (
            .O(N__49956),
            .I(n1196));
    InMux I__11246 (
            .O(N__49953),
            .I(N__49950));
    LocalMux I__11245 (
            .O(N__49950),
            .I(N__49947));
    Span4Mux_h I__11244 (
            .O(N__49947),
            .I(N__49944));
    Span4Mux_h I__11243 (
            .O(N__49944),
            .I(N__49938));
    CascadeMux I__11242 (
            .O(N__49943),
            .I(N__49935));
    CascadeMux I__11241 (
            .O(N__49942),
            .I(N__49931));
    InMux I__11240 (
            .O(N__49941),
            .I(N__49925));
    Span4Mux_v I__11239 (
            .O(N__49938),
            .I(N__49919));
    InMux I__11238 (
            .O(N__49935),
            .I(N__49916));
    InMux I__11237 (
            .O(N__49934),
            .I(N__49913));
    InMux I__11236 (
            .O(N__49931),
            .I(N__49904));
    InMux I__11235 (
            .O(N__49930),
            .I(N__49904));
    InMux I__11234 (
            .O(N__49929),
            .I(N__49904));
    InMux I__11233 (
            .O(N__49928),
            .I(N__49904));
    LocalMux I__11232 (
            .O(N__49925),
            .I(N__49901));
    InMux I__11231 (
            .O(N__49924),
            .I(N__49894));
    InMux I__11230 (
            .O(N__49923),
            .I(N__49894));
    InMux I__11229 (
            .O(N__49922),
            .I(N__49894));
    Odrv4 I__11228 (
            .O(N__49919),
            .I(n1158));
    LocalMux I__11227 (
            .O(N__49916),
            .I(n1158));
    LocalMux I__11226 (
            .O(N__49913),
            .I(n1158));
    LocalMux I__11225 (
            .O(N__49904),
            .I(n1158));
    Odrv4 I__11224 (
            .O(N__49901),
            .I(n1158));
    LocalMux I__11223 (
            .O(N__49894),
            .I(n1158));
    InMux I__11222 (
            .O(N__49881),
            .I(N__49878));
    LocalMux I__11221 (
            .O(N__49878),
            .I(N__49872));
    InMux I__11220 (
            .O(N__49877),
            .I(N__49869));
    CascadeMux I__11219 (
            .O(N__49876),
            .I(N__49864));
    CascadeMux I__11218 (
            .O(N__49875),
            .I(N__49861));
    Span4Mux_h I__11217 (
            .O(N__49872),
            .I(N__49855));
    LocalMux I__11216 (
            .O(N__49869),
            .I(N__49855));
    CascadeMux I__11215 (
            .O(N__49868),
            .I(N__49851));
    CascadeMux I__11214 (
            .O(N__49867),
            .I(N__49848));
    InMux I__11213 (
            .O(N__49864),
            .I(N__49843));
    InMux I__11212 (
            .O(N__49861),
            .I(N__49843));
    CascadeMux I__11211 (
            .O(N__49860),
            .I(N__49838));
    Span4Mux_v I__11210 (
            .O(N__49855),
            .I(N__49835));
    InMux I__11209 (
            .O(N__49854),
            .I(N__49832));
    InMux I__11208 (
            .O(N__49851),
            .I(N__49827));
    InMux I__11207 (
            .O(N__49848),
            .I(N__49827));
    LocalMux I__11206 (
            .O(N__49843),
            .I(N__49824));
    InMux I__11205 (
            .O(N__49842),
            .I(N__49817));
    InMux I__11204 (
            .O(N__49841),
            .I(N__49817));
    InMux I__11203 (
            .O(N__49838),
            .I(N__49817));
    Odrv4 I__11202 (
            .O(N__49835),
            .I(n1059));
    LocalMux I__11201 (
            .O(N__49832),
            .I(n1059));
    LocalMux I__11200 (
            .O(N__49827),
            .I(n1059));
    Odrv4 I__11199 (
            .O(N__49824),
            .I(n1059));
    LocalMux I__11198 (
            .O(N__49817),
            .I(n1059));
    InMux I__11197 (
            .O(N__49806),
            .I(N__49802));
    CascadeMux I__11196 (
            .O(N__49805),
            .I(N__49798));
    LocalMux I__11195 (
            .O(N__49802),
            .I(N__49795));
    InMux I__11194 (
            .O(N__49801),
            .I(N__49792));
    InMux I__11193 (
            .O(N__49798),
            .I(N__49789));
    Odrv4 I__11192 (
            .O(N__49795),
            .I(n1128));
    LocalMux I__11191 (
            .O(N__49792),
            .I(n1128));
    LocalMux I__11190 (
            .O(N__49789),
            .I(n1128));
    CascadeMux I__11189 (
            .O(N__49782),
            .I(N__49779));
    InMux I__11188 (
            .O(N__49779),
            .I(N__49776));
    LocalMux I__11187 (
            .O(N__49776),
            .I(N__49773));
    Odrv4 I__11186 (
            .O(N__49773),
            .I(n1693));
    CascadeMux I__11185 (
            .O(N__49770),
            .I(N__49767));
    InMux I__11184 (
            .O(N__49767),
            .I(N__49764));
    LocalMux I__11183 (
            .O(N__49764),
            .I(N__49759));
    InMux I__11182 (
            .O(N__49763),
            .I(N__49756));
    InMux I__11181 (
            .O(N__49762),
            .I(N__49753));
    Span4Mux_h I__11180 (
            .O(N__49759),
            .I(N__49748));
    LocalMux I__11179 (
            .O(N__49756),
            .I(N__49748));
    LocalMux I__11178 (
            .O(N__49753),
            .I(encoder0_position_target_0));
    Odrv4 I__11177 (
            .O(N__49748),
            .I(encoder0_position_target_0));
    InMux I__11176 (
            .O(N__49743),
            .I(n12449));
    CascadeMux I__11175 (
            .O(N__49740),
            .I(N__49737));
    InMux I__11174 (
            .O(N__49737),
            .I(N__49732));
    CascadeMux I__11173 (
            .O(N__49736),
            .I(N__49729));
    CascadeMux I__11172 (
            .O(N__49735),
            .I(N__49726));
    LocalMux I__11171 (
            .O(N__49732),
            .I(N__49723));
    InMux I__11170 (
            .O(N__49729),
            .I(N__49720));
    InMux I__11169 (
            .O(N__49726),
            .I(N__49717));
    Sp12to4 I__11168 (
            .O(N__49723),
            .I(N__49712));
    LocalMux I__11167 (
            .O(N__49720),
            .I(N__49712));
    LocalMux I__11166 (
            .O(N__49717),
            .I(encoder0_position_target_1));
    Odrv12 I__11165 (
            .O(N__49712),
            .I(encoder0_position_target_1));
    InMux I__11164 (
            .O(N__49707),
            .I(n12450));
    CascadeMux I__11163 (
            .O(N__49704),
            .I(N__49700));
    CascadeMux I__11162 (
            .O(N__49703),
            .I(N__49696));
    InMux I__11161 (
            .O(N__49700),
            .I(N__49693));
    InMux I__11160 (
            .O(N__49699),
            .I(N__49690));
    InMux I__11159 (
            .O(N__49696),
            .I(N__49687));
    LocalMux I__11158 (
            .O(N__49693),
            .I(N__49684));
    LocalMux I__11157 (
            .O(N__49690),
            .I(N__49681));
    LocalMux I__11156 (
            .O(N__49687),
            .I(encoder0_position_target_2));
    Odrv12 I__11155 (
            .O(N__49684),
            .I(encoder0_position_target_2));
    Odrv4 I__11154 (
            .O(N__49681),
            .I(encoder0_position_target_2));
    InMux I__11153 (
            .O(N__49674),
            .I(n12451));
    CascadeMux I__11152 (
            .O(N__49671),
            .I(n1257_cascade_));
    CascadeMux I__11151 (
            .O(N__49668),
            .I(N__49665));
    InMux I__11150 (
            .O(N__49665),
            .I(N__49661));
    CascadeMux I__11149 (
            .O(N__49664),
            .I(N__49658));
    LocalMux I__11148 (
            .O(N__49661),
            .I(N__49654));
    InMux I__11147 (
            .O(N__49658),
            .I(N__49651));
    InMux I__11146 (
            .O(N__49657),
            .I(N__49648));
    Odrv4 I__11145 (
            .O(N__49654),
            .I(n1325));
    LocalMux I__11144 (
            .O(N__49651),
            .I(n1325));
    LocalMux I__11143 (
            .O(N__49648),
            .I(n1325));
    InMux I__11142 (
            .O(N__49641),
            .I(N__49638));
    LocalMux I__11141 (
            .O(N__49638),
            .I(N__49635));
    Span4Mux_h I__11140 (
            .O(N__49635),
            .I(N__49632));
    Span4Mux_h I__11139 (
            .O(N__49632),
            .I(N__49629));
    Odrv4 I__11138 (
            .O(N__49629),
            .I(n12));
    InMux I__11137 (
            .O(N__49626),
            .I(N__49612));
    InMux I__11136 (
            .O(N__49625),
            .I(N__49612));
    InMux I__11135 (
            .O(N__49624),
            .I(N__49612));
    InMux I__11134 (
            .O(N__49623),
            .I(N__49612));
    InMux I__11133 (
            .O(N__49622),
            .I(N__49607));
    InMux I__11132 (
            .O(N__49621),
            .I(N__49594));
    LocalMux I__11131 (
            .O(N__49612),
            .I(N__49586));
    InMux I__11130 (
            .O(N__49611),
            .I(N__49581));
    InMux I__11129 (
            .O(N__49610),
            .I(N__49581));
    LocalMux I__11128 (
            .O(N__49607),
            .I(N__49577));
    InMux I__11127 (
            .O(N__49606),
            .I(N__49574));
    InMux I__11126 (
            .O(N__49605),
            .I(N__49569));
    InMux I__11125 (
            .O(N__49604),
            .I(N__49569));
    InMux I__11124 (
            .O(N__49603),
            .I(N__49566));
    InMux I__11123 (
            .O(N__49602),
            .I(N__49561));
    InMux I__11122 (
            .O(N__49601),
            .I(N__49561));
    InMux I__11121 (
            .O(N__49600),
            .I(N__49557));
    InMux I__11120 (
            .O(N__49599),
            .I(N__49554));
    CascadeMux I__11119 (
            .O(N__49598),
            .I(N__49549));
    CascadeMux I__11118 (
            .O(N__49597),
            .I(N__49543));
    LocalMux I__11117 (
            .O(N__49594),
            .I(N__49535));
    InMux I__11116 (
            .O(N__49593),
            .I(N__49528));
    InMux I__11115 (
            .O(N__49592),
            .I(N__49528));
    InMux I__11114 (
            .O(N__49591),
            .I(N__49528));
    InMux I__11113 (
            .O(N__49590),
            .I(N__49523));
    InMux I__11112 (
            .O(N__49589),
            .I(N__49523));
    Span4Mux_h I__11111 (
            .O(N__49586),
            .I(N__49518));
    LocalMux I__11110 (
            .O(N__49581),
            .I(N__49518));
    CascadeMux I__11109 (
            .O(N__49580),
            .I(N__49514));
    Span4Mux_v I__11108 (
            .O(N__49577),
            .I(N__49508));
    LocalMux I__11107 (
            .O(N__49574),
            .I(N__49508));
    LocalMux I__11106 (
            .O(N__49569),
            .I(N__49505));
    LocalMux I__11105 (
            .O(N__49566),
            .I(N__49500));
    LocalMux I__11104 (
            .O(N__49561),
            .I(N__49500));
    InMux I__11103 (
            .O(N__49560),
            .I(N__49497));
    LocalMux I__11102 (
            .O(N__49557),
            .I(N__49488));
    LocalMux I__11101 (
            .O(N__49554),
            .I(N__49488));
    CascadeMux I__11100 (
            .O(N__49553),
            .I(N__49485));
    CascadeMux I__11099 (
            .O(N__49552),
            .I(N__49482));
    InMux I__11098 (
            .O(N__49549),
            .I(N__49469));
    InMux I__11097 (
            .O(N__49548),
            .I(N__49469));
    InMux I__11096 (
            .O(N__49547),
            .I(N__49469));
    InMux I__11095 (
            .O(N__49546),
            .I(N__49469));
    InMux I__11094 (
            .O(N__49543),
            .I(N__49469));
    InMux I__11093 (
            .O(N__49542),
            .I(N__49469));
    InMux I__11092 (
            .O(N__49541),
            .I(N__49466));
    InMux I__11091 (
            .O(N__49540),
            .I(N__49463));
    InMux I__11090 (
            .O(N__49539),
            .I(N__49460));
    InMux I__11089 (
            .O(N__49538),
            .I(N__49457));
    Span4Mux_v I__11088 (
            .O(N__49535),
            .I(N__49452));
    LocalMux I__11087 (
            .O(N__49528),
            .I(N__49452));
    LocalMux I__11086 (
            .O(N__49523),
            .I(N__49447));
    Span4Mux_h I__11085 (
            .O(N__49518),
            .I(N__49447));
    InMux I__11084 (
            .O(N__49517),
            .I(N__49440));
    InMux I__11083 (
            .O(N__49514),
            .I(N__49440));
    InMux I__11082 (
            .O(N__49513),
            .I(N__49440));
    Span4Mux_h I__11081 (
            .O(N__49508),
            .I(N__49437));
    Span4Mux_h I__11080 (
            .O(N__49505),
            .I(N__49430));
    Span4Mux_h I__11079 (
            .O(N__49500),
            .I(N__49430));
    LocalMux I__11078 (
            .O(N__49497),
            .I(N__49430));
    InMux I__11077 (
            .O(N__49496),
            .I(N__49427));
    InMux I__11076 (
            .O(N__49495),
            .I(N__49420));
    InMux I__11075 (
            .O(N__49494),
            .I(N__49420));
    InMux I__11074 (
            .O(N__49493),
            .I(N__49420));
    Span4Mux_h I__11073 (
            .O(N__49488),
            .I(N__49417));
    InMux I__11072 (
            .O(N__49485),
            .I(N__49412));
    InMux I__11071 (
            .O(N__49482),
            .I(N__49412));
    LocalMux I__11070 (
            .O(N__49469),
            .I(N__49407));
    LocalMux I__11069 (
            .O(N__49466),
            .I(N__49407));
    LocalMux I__11068 (
            .O(N__49463),
            .I(encoder0_position_31));
    LocalMux I__11067 (
            .O(N__49460),
            .I(encoder0_position_31));
    LocalMux I__11066 (
            .O(N__49457),
            .I(encoder0_position_31));
    Odrv4 I__11065 (
            .O(N__49452),
            .I(encoder0_position_31));
    Odrv4 I__11064 (
            .O(N__49447),
            .I(encoder0_position_31));
    LocalMux I__11063 (
            .O(N__49440),
            .I(encoder0_position_31));
    Odrv4 I__11062 (
            .O(N__49437),
            .I(encoder0_position_31));
    Odrv4 I__11061 (
            .O(N__49430),
            .I(encoder0_position_31));
    LocalMux I__11060 (
            .O(N__49427),
            .I(encoder0_position_31));
    LocalMux I__11059 (
            .O(N__49420),
            .I(encoder0_position_31));
    Odrv4 I__11058 (
            .O(N__49417),
            .I(encoder0_position_31));
    LocalMux I__11057 (
            .O(N__49412),
            .I(encoder0_position_31));
    Odrv12 I__11056 (
            .O(N__49407),
            .I(encoder0_position_31));
    CascadeMux I__11055 (
            .O(N__49380),
            .I(N__49377));
    InMux I__11054 (
            .O(N__49377),
            .I(N__49373));
    CascadeMux I__11053 (
            .O(N__49376),
            .I(N__49370));
    LocalMux I__11052 (
            .O(N__49373),
            .I(N__49366));
    InMux I__11051 (
            .O(N__49370),
            .I(N__49363));
    InMux I__11050 (
            .O(N__49369),
            .I(N__49360));
    Odrv4 I__11049 (
            .O(N__49366),
            .I(n1326));
    LocalMux I__11048 (
            .O(N__49363),
            .I(n1326));
    LocalMux I__11047 (
            .O(N__49360),
            .I(n1326));
    InMux I__11046 (
            .O(N__49353),
            .I(N__49350));
    LocalMux I__11045 (
            .O(N__49350),
            .I(n1195));
    CascadeMux I__11044 (
            .O(N__49347),
            .I(n1227_cascade_));
    InMux I__11043 (
            .O(N__49344),
            .I(N__49341));
    LocalMux I__11042 (
            .O(N__49341),
            .I(n14476));
    InMux I__11041 (
            .O(N__49338),
            .I(N__49335));
    LocalMux I__11040 (
            .O(N__49335),
            .I(n1199));
    CascadeMux I__11039 (
            .O(N__49332),
            .I(N__49329));
    InMux I__11038 (
            .O(N__49329),
            .I(N__49325));
    CascadeMux I__11037 (
            .O(N__49328),
            .I(N__49322));
    LocalMux I__11036 (
            .O(N__49325),
            .I(N__49319));
    InMux I__11035 (
            .O(N__49322),
            .I(N__49316));
    Odrv4 I__11034 (
            .O(N__49319),
            .I(n1132));
    LocalMux I__11033 (
            .O(N__49316),
            .I(n1132));
    CascadeMux I__11032 (
            .O(N__49311),
            .I(N__49308));
    InMux I__11031 (
            .O(N__49308),
            .I(N__49304));
    InMux I__11030 (
            .O(N__49307),
            .I(N__49301));
    LocalMux I__11029 (
            .O(N__49304),
            .I(n1127));
    LocalMux I__11028 (
            .O(N__49301),
            .I(n1127));
    InMux I__11027 (
            .O(N__49296),
            .I(N__49293));
    LocalMux I__11026 (
            .O(N__49293),
            .I(n1194));
    CascadeMux I__11025 (
            .O(N__49290),
            .I(n1127_cascade_));
    InMux I__11024 (
            .O(N__49287),
            .I(N__49283));
    CascadeMux I__11023 (
            .O(N__49286),
            .I(N__49280));
    LocalMux I__11022 (
            .O(N__49283),
            .I(N__49277));
    InMux I__11021 (
            .O(N__49280),
            .I(N__49274));
    Odrv4 I__11020 (
            .O(N__49277),
            .I(n1328));
    LocalMux I__11019 (
            .O(N__49274),
            .I(n1328));
    CascadeMux I__11018 (
            .O(N__49269),
            .I(n1328_cascade_));
    InMux I__11017 (
            .O(N__49266),
            .I(N__49263));
    LocalMux I__11016 (
            .O(N__49263),
            .I(n14414));
    CascadeMux I__11015 (
            .O(N__49260),
            .I(N__49257));
    InMux I__11014 (
            .O(N__49257),
            .I(N__49253));
    CascadeMux I__11013 (
            .O(N__49256),
            .I(N__49250));
    LocalMux I__11012 (
            .O(N__49253),
            .I(N__49246));
    InMux I__11011 (
            .O(N__49250),
            .I(N__49243));
    InMux I__11010 (
            .O(N__49249),
            .I(N__49240));
    Odrv4 I__11009 (
            .O(N__49246),
            .I(n1327));
    LocalMux I__11008 (
            .O(N__49243),
            .I(n1327));
    LocalMux I__11007 (
            .O(N__49240),
            .I(n1327));
    CascadeMux I__11006 (
            .O(N__49233),
            .I(N__49229));
    CascadeMux I__11005 (
            .O(N__49232),
            .I(N__49226));
    InMux I__11004 (
            .O(N__49229),
            .I(N__49222));
    InMux I__11003 (
            .O(N__49226),
            .I(N__49217));
    InMux I__11002 (
            .O(N__49225),
            .I(N__49217));
    LocalMux I__11001 (
            .O(N__49222),
            .I(n1331));
    LocalMux I__11000 (
            .O(N__49217),
            .I(n1331));
    CascadeMux I__10999 (
            .O(N__49212),
            .I(N__49209));
    InMux I__10998 (
            .O(N__49209),
            .I(N__49205));
    InMux I__10997 (
            .O(N__49208),
            .I(N__49202));
    LocalMux I__10996 (
            .O(N__49205),
            .I(n1332));
    LocalMux I__10995 (
            .O(N__49202),
            .I(n1332));
    InMux I__10994 (
            .O(N__49197),
            .I(N__49194));
    LocalMux I__10993 (
            .O(N__49194),
            .I(n1399));
    CascadeMux I__10992 (
            .O(N__49191),
            .I(n1332_cascade_));
    CascadeMux I__10991 (
            .O(N__49188),
            .I(N__49185));
    InMux I__10990 (
            .O(N__49185),
            .I(N__49181));
    CascadeMux I__10989 (
            .O(N__49184),
            .I(N__49178));
    LocalMux I__10988 (
            .O(N__49181),
            .I(N__49174));
    InMux I__10987 (
            .O(N__49178),
            .I(N__49171));
    InMux I__10986 (
            .O(N__49177),
            .I(N__49168));
    Odrv4 I__10985 (
            .O(N__49174),
            .I(n1329));
    LocalMux I__10984 (
            .O(N__49171),
            .I(n1329));
    LocalMux I__10983 (
            .O(N__49168),
            .I(n1329));
    InMux I__10982 (
            .O(N__49161),
            .I(N__49158));
    LocalMux I__10981 (
            .O(N__49158),
            .I(n11927));
    CascadeMux I__10980 (
            .O(N__49155),
            .I(n13723_cascade_));
    InMux I__10979 (
            .O(N__49152),
            .I(N__49149));
    LocalMux I__10978 (
            .O(N__49149),
            .I(n1394));
    InMux I__10977 (
            .O(N__49146),
            .I(N__49143));
    LocalMux I__10976 (
            .O(N__49143),
            .I(n1391));
    InMux I__10975 (
            .O(N__49140),
            .I(N__49135));
    InMux I__10974 (
            .O(N__49139),
            .I(N__49132));
    InMux I__10973 (
            .O(N__49138),
            .I(N__49129));
    LocalMux I__10972 (
            .O(N__49135),
            .I(N__49126));
    LocalMux I__10971 (
            .O(N__49132),
            .I(N__49121));
    LocalMux I__10970 (
            .O(N__49129),
            .I(N__49121));
    Span4Mux_h I__10969 (
            .O(N__49126),
            .I(N__49118));
    Odrv12 I__10968 (
            .O(N__49121),
            .I(n299));
    Odrv4 I__10967 (
            .O(N__49118),
            .I(n299));
    CascadeMux I__10966 (
            .O(N__49113),
            .I(n11925_cascade_));
    InMux I__10965 (
            .O(N__49110),
            .I(N__49107));
    LocalMux I__10964 (
            .O(N__49107),
            .I(n1398));
    CascadeMux I__10963 (
            .O(N__49104),
            .I(n1430_cascade_));
    InMux I__10962 (
            .O(N__49101),
            .I(N__49098));
    LocalMux I__10961 (
            .O(N__49098),
            .I(n13739));
    InMux I__10960 (
            .O(N__49095),
            .I(N__49092));
    LocalMux I__10959 (
            .O(N__49092),
            .I(n13720));
    InMux I__10958 (
            .O(N__49089),
            .I(N__49086));
    LocalMux I__10957 (
            .O(N__49086),
            .I(n1400));
    CascadeMux I__10956 (
            .O(N__49083),
            .I(n1356_cascade_));
    CascadeMux I__10955 (
            .O(N__49080),
            .I(N__49076));
    CascadeMux I__10954 (
            .O(N__49079),
            .I(N__49072));
    InMux I__10953 (
            .O(N__49076),
            .I(N__49069));
    InMux I__10952 (
            .O(N__49075),
            .I(N__49064));
    InMux I__10951 (
            .O(N__49072),
            .I(N__49064));
    LocalMux I__10950 (
            .O(N__49069),
            .I(n1333));
    LocalMux I__10949 (
            .O(N__49064),
            .I(n1333));
    CascadeMux I__10948 (
            .O(N__49059),
            .I(n1432_cascade_));
    InMux I__10947 (
            .O(N__49056),
            .I(N__49053));
    LocalMux I__10946 (
            .O(N__49053),
            .I(n11923));
    InMux I__10945 (
            .O(N__49050),
            .I(N__49047));
    LocalMux I__10944 (
            .O(N__49047),
            .I(N__49044));
    Odrv4 I__10943 (
            .O(N__49044),
            .I(n1393));
    CascadeMux I__10942 (
            .O(N__49041),
            .I(n1425_cascade_));
    InMux I__10941 (
            .O(N__49038),
            .I(N__49035));
    LocalMux I__10940 (
            .O(N__49035),
            .I(n14484));
    CascadeMux I__10939 (
            .O(N__49032),
            .I(n14490_cascade_));
    CascadeMux I__10938 (
            .O(N__49029),
            .I(n1455_cascade_));
    CascadeMux I__10937 (
            .O(N__49026),
            .I(n1531_cascade_));
    CascadeMux I__10936 (
            .O(N__49023),
            .I(N__49020));
    InMux I__10935 (
            .O(N__49020),
            .I(N__49017));
    LocalMux I__10934 (
            .O(N__49017),
            .I(n11997));
    CascadeMux I__10933 (
            .O(N__49014),
            .I(N__49011));
    InMux I__10932 (
            .O(N__49011),
            .I(N__49008));
    LocalMux I__10931 (
            .O(N__49008),
            .I(N__49004));
    CascadeMux I__10930 (
            .O(N__49007),
            .I(N__49001));
    Sp12to4 I__10929 (
            .O(N__49004),
            .I(N__48994));
    InMux I__10928 (
            .O(N__49001),
            .I(N__48988));
    CascadeMux I__10927 (
            .O(N__49000),
            .I(N__48984));
    CascadeMux I__10926 (
            .O(N__48999),
            .I(N__48981));
    CascadeMux I__10925 (
            .O(N__48998),
            .I(N__48977));
    CascadeMux I__10924 (
            .O(N__48997),
            .I(N__48973));
    Span12Mux_v I__10923 (
            .O(N__48994),
            .I(N__48969));
    InMux I__10922 (
            .O(N__48993),
            .I(N__48966));
    InMux I__10921 (
            .O(N__48992),
            .I(N__48961));
    InMux I__10920 (
            .O(N__48991),
            .I(N__48961));
    LocalMux I__10919 (
            .O(N__48988),
            .I(N__48958));
    InMux I__10918 (
            .O(N__48987),
            .I(N__48941));
    InMux I__10917 (
            .O(N__48984),
            .I(N__48941));
    InMux I__10916 (
            .O(N__48981),
            .I(N__48941));
    InMux I__10915 (
            .O(N__48980),
            .I(N__48941));
    InMux I__10914 (
            .O(N__48977),
            .I(N__48941));
    InMux I__10913 (
            .O(N__48976),
            .I(N__48941));
    InMux I__10912 (
            .O(N__48973),
            .I(N__48941));
    InMux I__10911 (
            .O(N__48972),
            .I(N__48941));
    Odrv12 I__10910 (
            .O(N__48969),
            .I(n1455));
    LocalMux I__10909 (
            .O(N__48966),
            .I(n1455));
    LocalMux I__10908 (
            .O(N__48961),
            .I(n1455));
    Odrv4 I__10907 (
            .O(N__48958),
            .I(n1455));
    LocalMux I__10906 (
            .O(N__48941),
            .I(n1455));
    CascadeMux I__10905 (
            .O(N__48930),
            .I(N__48927));
    InMux I__10904 (
            .O(N__48927),
            .I(N__48923));
    CascadeMux I__10903 (
            .O(N__48926),
            .I(N__48920));
    LocalMux I__10902 (
            .O(N__48923),
            .I(N__48917));
    InMux I__10901 (
            .O(N__48920),
            .I(N__48914));
    Span4Mux_v I__10900 (
            .O(N__48917),
            .I(N__48908));
    LocalMux I__10899 (
            .O(N__48914),
            .I(N__48908));
    InMux I__10898 (
            .O(N__48913),
            .I(N__48905));
    Odrv4 I__10897 (
            .O(N__48908),
            .I(n1631_adj_611));
    LocalMux I__10896 (
            .O(N__48905),
            .I(n1631_adj_611));
    InMux I__10895 (
            .O(N__48900),
            .I(N__48897));
    LocalMux I__10894 (
            .O(N__48897),
            .I(N__48894));
    Span4Mux_v I__10893 (
            .O(N__48894),
            .I(N__48890));
    CascadeMux I__10892 (
            .O(N__48893),
            .I(N__48887));
    Sp12to4 I__10891 (
            .O(N__48890),
            .I(N__48881));
    InMux I__10890 (
            .O(N__48887),
            .I(N__48878));
    CascadeMux I__10889 (
            .O(N__48886),
            .I(N__48871));
    CascadeMux I__10888 (
            .O(N__48885),
            .I(N__48867));
    CascadeMux I__10887 (
            .O(N__48884),
            .I(N__48863));
    Span12Mux_h I__10886 (
            .O(N__48881),
            .I(N__48857));
    LocalMux I__10885 (
            .O(N__48878),
            .I(N__48854));
    InMux I__10884 (
            .O(N__48877),
            .I(N__48851));
    InMux I__10883 (
            .O(N__48876),
            .I(N__48844));
    InMux I__10882 (
            .O(N__48875),
            .I(N__48844));
    InMux I__10881 (
            .O(N__48874),
            .I(N__48844));
    InMux I__10880 (
            .O(N__48871),
            .I(N__48839));
    InMux I__10879 (
            .O(N__48870),
            .I(N__48839));
    InMux I__10878 (
            .O(N__48867),
            .I(N__48834));
    InMux I__10877 (
            .O(N__48866),
            .I(N__48834));
    InMux I__10876 (
            .O(N__48863),
            .I(N__48825));
    InMux I__10875 (
            .O(N__48862),
            .I(N__48825));
    InMux I__10874 (
            .O(N__48861),
            .I(N__48825));
    InMux I__10873 (
            .O(N__48860),
            .I(N__48825));
    Odrv12 I__10872 (
            .O(N__48857),
            .I(n1554));
    Odrv4 I__10871 (
            .O(N__48854),
            .I(n1554));
    LocalMux I__10870 (
            .O(N__48851),
            .I(n1554));
    LocalMux I__10869 (
            .O(N__48844),
            .I(n1554));
    LocalMux I__10868 (
            .O(N__48839),
            .I(n1554));
    LocalMux I__10867 (
            .O(N__48834),
            .I(n1554));
    LocalMux I__10866 (
            .O(N__48825),
            .I(n1554));
    InMux I__10865 (
            .O(N__48810),
            .I(N__48806));
    CascadeMux I__10864 (
            .O(N__48809),
            .I(N__48803));
    LocalMux I__10863 (
            .O(N__48806),
            .I(N__48800));
    InMux I__10862 (
            .O(N__48803),
            .I(N__48797));
    Span4Mux_v I__10861 (
            .O(N__48800),
            .I(N__48792));
    LocalMux I__10860 (
            .O(N__48797),
            .I(N__48792));
    Odrv4 I__10859 (
            .O(N__48792),
            .I(n1632_adj_612));
    InMux I__10858 (
            .O(N__48789),
            .I(N__48784));
    InMux I__10857 (
            .O(N__48788),
            .I(N__48781));
    InMux I__10856 (
            .O(N__48787),
            .I(N__48778));
    LocalMux I__10855 (
            .O(N__48784),
            .I(N__48775));
    LocalMux I__10854 (
            .O(N__48781),
            .I(N__48770));
    LocalMux I__10853 (
            .O(N__48778),
            .I(N__48770));
    Span4Mux_h I__10852 (
            .O(N__48775),
            .I(N__48767));
    Span4Mux_h I__10851 (
            .O(N__48770),
            .I(N__48764));
    Odrv4 I__10850 (
            .O(N__48767),
            .I(n302));
    Odrv4 I__10849 (
            .O(N__48764),
            .I(n302));
    CascadeMux I__10848 (
            .O(N__48759),
            .I(n1632_adj_612_cascade_));
    CascadeMux I__10847 (
            .O(N__48756),
            .I(N__48753));
    InMux I__10846 (
            .O(N__48753),
            .I(N__48750));
    LocalMux I__10845 (
            .O(N__48750),
            .I(N__48746));
    CascadeMux I__10844 (
            .O(N__48749),
            .I(N__48743));
    Span4Mux_h I__10843 (
            .O(N__48746),
            .I(N__48739));
    InMux I__10842 (
            .O(N__48743),
            .I(N__48736));
    InMux I__10841 (
            .O(N__48742),
            .I(N__48733));
    Odrv4 I__10840 (
            .O(N__48739),
            .I(n1633_adj_613));
    LocalMux I__10839 (
            .O(N__48736),
            .I(n1633_adj_613));
    LocalMux I__10838 (
            .O(N__48733),
            .I(n1633_adj_613));
    InMux I__10837 (
            .O(N__48726),
            .I(N__48723));
    LocalMux I__10836 (
            .O(N__48723),
            .I(n11919));
    InMux I__10835 (
            .O(N__48720),
            .I(\PWM.n13047 ));
    InMux I__10834 (
            .O(N__48717),
            .I(\PWM.n13048 ));
    InMux I__10833 (
            .O(N__48714),
            .I(\PWM.n13049 ));
    InMux I__10832 (
            .O(N__48711),
            .I(\PWM.n13050 ));
    InMux I__10831 (
            .O(N__48708),
            .I(\PWM.n13051 ));
    InMux I__10830 (
            .O(N__48705),
            .I(\PWM.n13052 ));
    SRMux I__10829 (
            .O(N__48702),
            .I(N__48699));
    LocalMux I__10828 (
            .O(N__48699),
            .I(N__48696));
    Span4Mux_h I__10827 (
            .O(N__48696),
            .I(N__48690));
    SRMux I__10826 (
            .O(N__48695),
            .I(N__48687));
    SRMux I__10825 (
            .O(N__48694),
            .I(N__48684));
    SRMux I__10824 (
            .O(N__48693),
            .I(N__48681));
    Odrv4 I__10823 (
            .O(N__48690),
            .I(\PWM.pwm_counter_31__N_407 ));
    LocalMux I__10822 (
            .O(N__48687),
            .I(\PWM.pwm_counter_31__N_407 ));
    LocalMux I__10821 (
            .O(N__48684),
            .I(\PWM.pwm_counter_31__N_407 ));
    LocalMux I__10820 (
            .O(N__48681),
            .I(\PWM.pwm_counter_31__N_407 ));
    InMux I__10819 (
            .O(N__48672),
            .I(N__48668));
    InMux I__10818 (
            .O(N__48671),
            .I(N__48665));
    LocalMux I__10817 (
            .O(N__48668),
            .I(pwm_counter_24));
    LocalMux I__10816 (
            .O(N__48665),
            .I(pwm_counter_24));
    InMux I__10815 (
            .O(N__48660),
            .I(N__48656));
    InMux I__10814 (
            .O(N__48659),
            .I(N__48653));
    LocalMux I__10813 (
            .O(N__48656),
            .I(pwm_counter_29));
    LocalMux I__10812 (
            .O(N__48653),
            .I(pwm_counter_29));
    CascadeMux I__10811 (
            .O(N__48648),
            .I(N__48644));
    InMux I__10810 (
            .O(N__48647),
            .I(N__48641));
    InMux I__10809 (
            .O(N__48644),
            .I(N__48638));
    LocalMux I__10808 (
            .O(N__48641),
            .I(pwm_counter_27));
    LocalMux I__10807 (
            .O(N__48638),
            .I(pwm_counter_27));
    InMux I__10806 (
            .O(N__48633),
            .I(N__48629));
    InMux I__10805 (
            .O(N__48632),
            .I(N__48626));
    LocalMux I__10804 (
            .O(N__48629),
            .I(pwm_counter_26));
    LocalMux I__10803 (
            .O(N__48626),
            .I(pwm_counter_26));
    InMux I__10802 (
            .O(N__48621),
            .I(N__48617));
    InMux I__10801 (
            .O(N__48620),
            .I(N__48614));
    LocalMux I__10800 (
            .O(N__48617),
            .I(pwm_counter_30));
    LocalMux I__10799 (
            .O(N__48614),
            .I(pwm_counter_30));
    InMux I__10798 (
            .O(N__48609),
            .I(N__48605));
    InMux I__10797 (
            .O(N__48608),
            .I(N__48602));
    LocalMux I__10796 (
            .O(N__48605),
            .I(pwm_counter_25));
    LocalMux I__10795 (
            .O(N__48602),
            .I(pwm_counter_25));
    CascadeMux I__10794 (
            .O(N__48597),
            .I(n12_adj_615_cascade_));
    InMux I__10793 (
            .O(N__48594),
            .I(N__48590));
    InMux I__10792 (
            .O(N__48593),
            .I(N__48587));
    LocalMux I__10791 (
            .O(N__48590),
            .I(pwm_counter_28));
    LocalMux I__10790 (
            .O(N__48587),
            .I(pwm_counter_28));
    InMux I__10789 (
            .O(N__48582),
            .I(N__48579));
    LocalMux I__10788 (
            .O(N__48579),
            .I(N__48574));
    InMux I__10787 (
            .O(N__48578),
            .I(N__48571));
    InMux I__10786 (
            .O(N__48577),
            .I(N__48568));
    Span4Mux_s2_v I__10785 (
            .O(N__48574),
            .I(N__48565));
    LocalMux I__10784 (
            .O(N__48571),
            .I(pwm_counter_17));
    LocalMux I__10783 (
            .O(N__48568),
            .I(pwm_counter_17));
    Odrv4 I__10782 (
            .O(N__48565),
            .I(pwm_counter_17));
    InMux I__10781 (
            .O(N__48558),
            .I(\PWM.n13038 ));
    InMux I__10780 (
            .O(N__48555),
            .I(N__48551));
    InMux I__10779 (
            .O(N__48554),
            .I(N__48547));
    LocalMux I__10778 (
            .O(N__48551),
            .I(N__48544));
    InMux I__10777 (
            .O(N__48550),
            .I(N__48541));
    LocalMux I__10776 (
            .O(N__48547),
            .I(N__48536));
    Span4Mux_s2_v I__10775 (
            .O(N__48544),
            .I(N__48536));
    LocalMux I__10774 (
            .O(N__48541),
            .I(pwm_counter_18));
    Odrv4 I__10773 (
            .O(N__48536),
            .I(pwm_counter_18));
    InMux I__10772 (
            .O(N__48531),
            .I(\PWM.n13039 ));
    InMux I__10771 (
            .O(N__48528),
            .I(N__48523));
    InMux I__10770 (
            .O(N__48527),
            .I(N__48520));
    InMux I__10769 (
            .O(N__48526),
            .I(N__48517));
    LocalMux I__10768 (
            .O(N__48523),
            .I(N__48514));
    LocalMux I__10767 (
            .O(N__48520),
            .I(pwm_counter_19));
    LocalMux I__10766 (
            .O(N__48517),
            .I(pwm_counter_19));
    Odrv4 I__10765 (
            .O(N__48514),
            .I(pwm_counter_19));
    InMux I__10764 (
            .O(N__48507),
            .I(\PWM.n13040 ));
    InMux I__10763 (
            .O(N__48504),
            .I(N__48501));
    LocalMux I__10762 (
            .O(N__48501),
            .I(N__48496));
    InMux I__10761 (
            .O(N__48500),
            .I(N__48493));
    InMux I__10760 (
            .O(N__48499),
            .I(N__48490));
    Span4Mux_h I__10759 (
            .O(N__48496),
            .I(N__48487));
    LocalMux I__10758 (
            .O(N__48493),
            .I(pwm_counter_20));
    LocalMux I__10757 (
            .O(N__48490),
            .I(pwm_counter_20));
    Odrv4 I__10756 (
            .O(N__48487),
            .I(pwm_counter_20));
    InMux I__10755 (
            .O(N__48480),
            .I(\PWM.n13041 ));
    CascadeMux I__10754 (
            .O(N__48477),
            .I(N__48472));
    InMux I__10753 (
            .O(N__48476),
            .I(N__48469));
    InMux I__10752 (
            .O(N__48475),
            .I(N__48464));
    InMux I__10751 (
            .O(N__48472),
            .I(N__48464));
    LocalMux I__10750 (
            .O(N__48469),
            .I(N__48459));
    LocalMux I__10749 (
            .O(N__48464),
            .I(N__48456));
    InMux I__10748 (
            .O(N__48463),
            .I(N__48453));
    InMux I__10747 (
            .O(N__48462),
            .I(N__48450));
    Span4Mux_h I__10746 (
            .O(N__48459),
            .I(N__48447));
    Span4Mux_h I__10745 (
            .O(N__48456),
            .I(N__48444));
    LocalMux I__10744 (
            .O(N__48453),
            .I(pwm_counter_21));
    LocalMux I__10743 (
            .O(N__48450),
            .I(pwm_counter_21));
    Odrv4 I__10742 (
            .O(N__48447),
            .I(pwm_counter_21));
    Odrv4 I__10741 (
            .O(N__48444),
            .I(pwm_counter_21));
    InMux I__10740 (
            .O(N__48435),
            .I(\PWM.n13042 ));
    InMux I__10739 (
            .O(N__48432),
            .I(N__48429));
    LocalMux I__10738 (
            .O(N__48429),
            .I(N__48424));
    InMux I__10737 (
            .O(N__48428),
            .I(N__48421));
    InMux I__10736 (
            .O(N__48427),
            .I(N__48418));
    Span4Mux_h I__10735 (
            .O(N__48424),
            .I(N__48415));
    LocalMux I__10734 (
            .O(N__48421),
            .I(pwm_counter_22));
    LocalMux I__10733 (
            .O(N__48418),
            .I(pwm_counter_22));
    Odrv4 I__10732 (
            .O(N__48415),
            .I(pwm_counter_22));
    InMux I__10731 (
            .O(N__48408),
            .I(\PWM.n13043 ));
    InMux I__10730 (
            .O(N__48405),
            .I(\PWM.n13044 ));
    InMux I__10729 (
            .O(N__48402),
            .I(bfn_14_31_0_));
    InMux I__10728 (
            .O(N__48399),
            .I(\PWM.n13046 ));
    InMux I__10727 (
            .O(N__48396),
            .I(N__48388));
    InMux I__10726 (
            .O(N__48395),
            .I(N__48388));
    InMux I__10725 (
            .O(N__48394),
            .I(N__48385));
    InMux I__10724 (
            .O(N__48393),
            .I(N__48382));
    LocalMux I__10723 (
            .O(N__48388),
            .I(N__48379));
    LocalMux I__10722 (
            .O(N__48385),
            .I(pwm_counter_9));
    LocalMux I__10721 (
            .O(N__48382),
            .I(pwm_counter_9));
    Odrv12 I__10720 (
            .O(N__48379),
            .I(pwm_counter_9));
    InMux I__10719 (
            .O(N__48372),
            .I(\PWM.n13030 ));
    InMux I__10718 (
            .O(N__48369),
            .I(N__48364));
    InMux I__10717 (
            .O(N__48368),
            .I(N__48361));
    InMux I__10716 (
            .O(N__48367),
            .I(N__48358));
    LocalMux I__10715 (
            .O(N__48364),
            .I(N__48355));
    LocalMux I__10714 (
            .O(N__48361),
            .I(pwm_counter_10));
    LocalMux I__10713 (
            .O(N__48358),
            .I(pwm_counter_10));
    Odrv4 I__10712 (
            .O(N__48355),
            .I(pwm_counter_10));
    InMux I__10711 (
            .O(N__48348),
            .I(\PWM.n13031 ));
    InMux I__10710 (
            .O(N__48345),
            .I(N__48341));
    InMux I__10709 (
            .O(N__48344),
            .I(N__48337));
    LocalMux I__10708 (
            .O(N__48341),
            .I(N__48334));
    InMux I__10707 (
            .O(N__48340),
            .I(N__48331));
    LocalMux I__10706 (
            .O(N__48337),
            .I(N__48328));
    Odrv4 I__10705 (
            .O(N__48334),
            .I(pwm_counter_11));
    LocalMux I__10704 (
            .O(N__48331),
            .I(pwm_counter_11));
    Odrv4 I__10703 (
            .O(N__48328),
            .I(pwm_counter_11));
    InMux I__10702 (
            .O(N__48321),
            .I(\PWM.n13032 ));
    InMux I__10701 (
            .O(N__48318),
            .I(N__48315));
    LocalMux I__10700 (
            .O(N__48315),
            .I(N__48310));
    InMux I__10699 (
            .O(N__48314),
            .I(N__48307));
    InMux I__10698 (
            .O(N__48313),
            .I(N__48304));
    Span4Mux_s3_v I__10697 (
            .O(N__48310),
            .I(N__48301));
    LocalMux I__10696 (
            .O(N__48307),
            .I(pwm_counter_12));
    LocalMux I__10695 (
            .O(N__48304),
            .I(pwm_counter_12));
    Odrv4 I__10694 (
            .O(N__48301),
            .I(pwm_counter_12));
    InMux I__10693 (
            .O(N__48294),
            .I(\PWM.n13033 ));
    InMux I__10692 (
            .O(N__48291),
            .I(N__48286));
    InMux I__10691 (
            .O(N__48290),
            .I(N__48283));
    InMux I__10690 (
            .O(N__48289),
            .I(N__48280));
    LocalMux I__10689 (
            .O(N__48286),
            .I(pwm_counter_13));
    LocalMux I__10688 (
            .O(N__48283),
            .I(pwm_counter_13));
    LocalMux I__10687 (
            .O(N__48280),
            .I(pwm_counter_13));
    InMux I__10686 (
            .O(N__48273),
            .I(\PWM.n13034 ));
    CascadeMux I__10685 (
            .O(N__48270),
            .I(N__48267));
    InMux I__10684 (
            .O(N__48267),
            .I(N__48262));
    InMux I__10683 (
            .O(N__48266),
            .I(N__48259));
    InMux I__10682 (
            .O(N__48265),
            .I(N__48256));
    LocalMux I__10681 (
            .O(N__48262),
            .I(N__48251));
    LocalMux I__10680 (
            .O(N__48259),
            .I(N__48251));
    LocalMux I__10679 (
            .O(N__48256),
            .I(pwm_counter_14));
    Odrv4 I__10678 (
            .O(N__48251),
            .I(pwm_counter_14));
    InMux I__10677 (
            .O(N__48246),
            .I(\PWM.n13035 ));
    CascadeMux I__10676 (
            .O(N__48243),
            .I(N__48239));
    InMux I__10675 (
            .O(N__48242),
            .I(N__48236));
    InMux I__10674 (
            .O(N__48239),
            .I(N__48232));
    LocalMux I__10673 (
            .O(N__48236),
            .I(N__48229));
    InMux I__10672 (
            .O(N__48235),
            .I(N__48226));
    LocalMux I__10671 (
            .O(N__48232),
            .I(N__48221));
    Span4Mux_h I__10670 (
            .O(N__48229),
            .I(N__48221));
    LocalMux I__10669 (
            .O(N__48226),
            .I(pwm_counter_15));
    Odrv4 I__10668 (
            .O(N__48221),
            .I(pwm_counter_15));
    InMux I__10667 (
            .O(N__48216),
            .I(\PWM.n13036 ));
    InMux I__10666 (
            .O(N__48213),
            .I(N__48203));
    InMux I__10665 (
            .O(N__48212),
            .I(N__48203));
    InMux I__10664 (
            .O(N__48211),
            .I(N__48203));
    CascadeMux I__10663 (
            .O(N__48210),
            .I(N__48199));
    LocalMux I__10662 (
            .O(N__48203),
            .I(N__48196));
    InMux I__10661 (
            .O(N__48202),
            .I(N__48193));
    InMux I__10660 (
            .O(N__48199),
            .I(N__48190));
    Span4Mux_s2_v I__10659 (
            .O(N__48196),
            .I(N__48187));
    LocalMux I__10658 (
            .O(N__48193),
            .I(pwm_counter_16));
    LocalMux I__10657 (
            .O(N__48190),
            .I(pwm_counter_16));
    Odrv4 I__10656 (
            .O(N__48187),
            .I(pwm_counter_16));
    InMux I__10655 (
            .O(N__48180),
            .I(bfn_14_30_0_));
    CascadeMux I__10654 (
            .O(N__48177),
            .I(N__48174));
    InMux I__10653 (
            .O(N__48174),
            .I(N__48170));
    InMux I__10652 (
            .O(N__48173),
            .I(N__48167));
    LocalMux I__10651 (
            .O(N__48170),
            .I(N__48164));
    LocalMux I__10650 (
            .O(N__48167),
            .I(pwm_counter_0));
    Odrv4 I__10649 (
            .O(N__48164),
            .I(pwm_counter_0));
    InMux I__10648 (
            .O(N__48159),
            .I(bfn_14_28_0_));
    InMux I__10647 (
            .O(N__48156),
            .I(N__48152));
    InMux I__10646 (
            .O(N__48155),
            .I(N__48149));
    LocalMux I__10645 (
            .O(N__48152),
            .I(N__48146));
    LocalMux I__10644 (
            .O(N__48149),
            .I(pwm_counter_1));
    Odrv4 I__10643 (
            .O(N__48146),
            .I(pwm_counter_1));
    InMux I__10642 (
            .O(N__48141),
            .I(\PWM.n13022 ));
    CascadeMux I__10641 (
            .O(N__48138),
            .I(N__48134));
    InMux I__10640 (
            .O(N__48137),
            .I(N__48131));
    InMux I__10639 (
            .O(N__48134),
            .I(N__48128));
    LocalMux I__10638 (
            .O(N__48131),
            .I(pwm_counter_2));
    LocalMux I__10637 (
            .O(N__48128),
            .I(pwm_counter_2));
    InMux I__10636 (
            .O(N__48123),
            .I(\PWM.n13023 ));
    InMux I__10635 (
            .O(N__48120),
            .I(N__48115));
    InMux I__10634 (
            .O(N__48119),
            .I(N__48110));
    InMux I__10633 (
            .O(N__48118),
            .I(N__48110));
    LocalMux I__10632 (
            .O(N__48115),
            .I(pwm_counter_3));
    LocalMux I__10631 (
            .O(N__48110),
            .I(pwm_counter_3));
    InMux I__10630 (
            .O(N__48105),
            .I(\PWM.n13024 ));
    InMux I__10629 (
            .O(N__48102),
            .I(N__48099));
    LocalMux I__10628 (
            .O(N__48099),
            .I(N__48095));
    InMux I__10627 (
            .O(N__48098),
            .I(N__48092));
    Span4Mux_h I__10626 (
            .O(N__48095),
            .I(N__48089));
    LocalMux I__10625 (
            .O(N__48092),
            .I(pwm_counter_4));
    Odrv4 I__10624 (
            .O(N__48089),
            .I(pwm_counter_4));
    InMux I__10623 (
            .O(N__48084),
            .I(\PWM.n13025 ));
    InMux I__10622 (
            .O(N__48081),
            .I(N__48076));
    InMux I__10621 (
            .O(N__48080),
            .I(N__48073));
    InMux I__10620 (
            .O(N__48079),
            .I(N__48070));
    LocalMux I__10619 (
            .O(N__48076),
            .I(N__48067));
    LocalMux I__10618 (
            .O(N__48073),
            .I(pwm_counter_5));
    LocalMux I__10617 (
            .O(N__48070),
            .I(pwm_counter_5));
    Odrv4 I__10616 (
            .O(N__48067),
            .I(pwm_counter_5));
    InMux I__10615 (
            .O(N__48060),
            .I(\PWM.n13026 ));
    InMux I__10614 (
            .O(N__48057),
            .I(N__48053));
    InMux I__10613 (
            .O(N__48056),
            .I(N__48050));
    LocalMux I__10612 (
            .O(N__48053),
            .I(N__48045));
    LocalMux I__10611 (
            .O(N__48050),
            .I(N__48042));
    InMux I__10610 (
            .O(N__48049),
            .I(N__48039));
    InMux I__10609 (
            .O(N__48048),
            .I(N__48036));
    Span4Mux_h I__10608 (
            .O(N__48045),
            .I(N__48033));
    Span4Mux_h I__10607 (
            .O(N__48042),
            .I(N__48030));
    LocalMux I__10606 (
            .O(N__48039),
            .I(pwm_counter_6));
    LocalMux I__10605 (
            .O(N__48036),
            .I(pwm_counter_6));
    Odrv4 I__10604 (
            .O(N__48033),
            .I(pwm_counter_6));
    Odrv4 I__10603 (
            .O(N__48030),
            .I(pwm_counter_6));
    InMux I__10602 (
            .O(N__48021),
            .I(\PWM.n13027 ));
    InMux I__10601 (
            .O(N__48018),
            .I(N__48014));
    InMux I__10600 (
            .O(N__48017),
            .I(N__48011));
    LocalMux I__10599 (
            .O(N__48014),
            .I(N__48006));
    LocalMux I__10598 (
            .O(N__48011),
            .I(N__48003));
    InMux I__10597 (
            .O(N__48010),
            .I(N__48000));
    InMux I__10596 (
            .O(N__48009),
            .I(N__47997));
    Span4Mux_h I__10595 (
            .O(N__48006),
            .I(N__47994));
    Span4Mux_h I__10594 (
            .O(N__48003),
            .I(N__47991));
    LocalMux I__10593 (
            .O(N__48000),
            .I(pwm_counter_7));
    LocalMux I__10592 (
            .O(N__47997),
            .I(pwm_counter_7));
    Odrv4 I__10591 (
            .O(N__47994),
            .I(pwm_counter_7));
    Odrv4 I__10590 (
            .O(N__47991),
            .I(pwm_counter_7));
    InMux I__10589 (
            .O(N__47982),
            .I(\PWM.n13028 ));
    InMux I__10588 (
            .O(N__47979),
            .I(N__47974));
    InMux I__10587 (
            .O(N__47978),
            .I(N__47971));
    CascadeMux I__10586 (
            .O(N__47977),
            .I(N__47968));
    LocalMux I__10585 (
            .O(N__47974),
            .I(N__47964));
    LocalMux I__10584 (
            .O(N__47971),
            .I(N__47961));
    InMux I__10583 (
            .O(N__47968),
            .I(N__47958));
    InMux I__10582 (
            .O(N__47967),
            .I(N__47955));
    Span4Mux_h I__10581 (
            .O(N__47964),
            .I(N__47950));
    Span4Mux_h I__10580 (
            .O(N__47961),
            .I(N__47950));
    LocalMux I__10579 (
            .O(N__47958),
            .I(pwm_counter_8));
    LocalMux I__10578 (
            .O(N__47955),
            .I(pwm_counter_8));
    Odrv4 I__10577 (
            .O(N__47950),
            .I(pwm_counter_8));
    InMux I__10576 (
            .O(N__47943),
            .I(bfn_14_29_0_));
    InMux I__10575 (
            .O(N__47940),
            .I(N__47937));
    LocalMux I__10574 (
            .O(N__47937),
            .I(N__47934));
    Span4Mux_h I__10573 (
            .O(N__47934),
            .I(N__47931));
    Odrv4 I__10572 (
            .O(N__47931),
            .I(pwm_setpoint_1));
    CascadeMux I__10571 (
            .O(N__47928),
            .I(n16_adj_679_cascade_));
    InMux I__10570 (
            .O(N__47925),
            .I(N__47922));
    LocalMux I__10569 (
            .O(N__47922),
            .I(n15_adj_680));
    InMux I__10568 (
            .O(N__47919),
            .I(N__47916));
    LocalMux I__10567 (
            .O(N__47916),
            .I(n25_adj_652));
    CascadeMux I__10566 (
            .O(N__47913),
            .I(n16_adj_619_cascade_));
    InMux I__10565 (
            .O(N__47910),
            .I(N__47907));
    LocalMux I__10564 (
            .O(N__47907),
            .I(n22_adj_617));
    InMux I__10563 (
            .O(N__47904),
            .I(N__47901));
    LocalMux I__10562 (
            .O(N__47901),
            .I(N__47898));
    Odrv4 I__10561 (
            .O(N__47898),
            .I(n24_adj_616));
    InMux I__10560 (
            .O(N__47895),
            .I(N__47892));
    LocalMux I__10559 (
            .O(N__47892),
            .I(N__47889));
    Span4Mux_h I__10558 (
            .O(N__47889),
            .I(N__47886));
    Odrv4 I__10557 (
            .O(N__47886),
            .I(encoder0_position_scaled_16));
    InMux I__10556 (
            .O(N__47883),
            .I(N__47880));
    LocalMux I__10555 (
            .O(N__47880),
            .I(N__47877));
    Odrv4 I__10554 (
            .O(N__47877),
            .I(n9_adj_567));
    InMux I__10553 (
            .O(N__47874),
            .I(N__47870));
    InMux I__10552 (
            .O(N__47873),
            .I(N__47867));
    LocalMux I__10551 (
            .O(N__47870),
            .I(N__47864));
    LocalMux I__10550 (
            .O(N__47867),
            .I(N__47861));
    Span4Mux_h I__10549 (
            .O(N__47864),
            .I(N__47858));
    Span4Mux_h I__10548 (
            .O(N__47861),
            .I(N__47855));
    Odrv4 I__10547 (
            .O(N__47858),
            .I(duty_1));
    Odrv4 I__10546 (
            .O(N__47855),
            .I(duty_1));
    InMux I__10545 (
            .O(N__47850),
            .I(N__47847));
    LocalMux I__10544 (
            .O(N__47847),
            .I(N__47844));
    Span4Mux_h I__10543 (
            .O(N__47844),
            .I(N__47841));
    Odrv4 I__10542 (
            .O(N__47841),
            .I(n24_adj_596));
    SRMux I__10541 (
            .O(N__47838),
            .I(N__47832));
    InMux I__10540 (
            .O(N__47837),
            .I(N__47832));
    LocalMux I__10539 (
            .O(N__47832),
            .I(N__47829));
    Span4Mux_h I__10538 (
            .O(N__47829),
            .I(N__47826));
    Odrv4 I__10537 (
            .O(N__47826),
            .I(pwm_setpoint_23__N_195));
    CascadeMux I__10536 (
            .O(N__47823),
            .I(n13197_cascade_));
    InMux I__10535 (
            .O(N__47820),
            .I(N__47817));
    LocalMux I__10534 (
            .O(N__47817),
            .I(n24_adj_653));
    CascadeMux I__10533 (
            .O(N__47814),
            .I(direction_N_342_cascade_));
    InMux I__10532 (
            .O(N__47811),
            .I(N__47808));
    LocalMux I__10531 (
            .O(N__47808),
            .I(direction_N_342));
    InMux I__10530 (
            .O(N__47805),
            .I(N__47802));
    LocalMux I__10529 (
            .O(N__47802),
            .I(n13675));
    CascadeMux I__10528 (
            .O(N__47799),
            .I(n23_adj_709_cascade_));
    InMux I__10527 (
            .O(N__47796),
            .I(N__47793));
    LocalMux I__10526 (
            .O(N__47793),
            .I(n25_adj_707));
    InMux I__10525 (
            .O(N__47790),
            .I(N__47786));
    InMux I__10524 (
            .O(N__47789),
            .I(N__47783));
    LocalMux I__10523 (
            .O(N__47786),
            .I(direction_N_340));
    LocalMux I__10522 (
            .O(N__47783),
            .I(direction_N_340));
    InMux I__10521 (
            .O(N__47778),
            .I(N__47775));
    LocalMux I__10520 (
            .O(N__47775),
            .I(n24_adj_708));
    InMux I__10519 (
            .O(N__47772),
            .I(N__47769));
    LocalMux I__10518 (
            .O(N__47769),
            .I(n23_adj_654));
    InMux I__10517 (
            .O(N__47766),
            .I(N__47763));
    LocalMux I__10516 (
            .O(N__47763),
            .I(N__47760));
    Odrv12 I__10515 (
            .O(N__47760),
            .I(pwm_setpoint_23_N_171_1));
    InMux I__10514 (
            .O(N__47757),
            .I(n12527));
    InMux I__10513 (
            .O(N__47754),
            .I(n12528));
    InMux I__10512 (
            .O(N__47751),
            .I(bfn_14_24_0_));
    InMux I__10511 (
            .O(N__47748),
            .I(n12530));
    InMux I__10510 (
            .O(N__47745),
            .I(N__47742));
    LocalMux I__10509 (
            .O(N__47742),
            .I(N__47739));
    Span12Mux_s8_v I__10508 (
            .O(N__47739),
            .I(N__47735));
    InMux I__10507 (
            .O(N__47738),
            .I(N__47732));
    Odrv12 I__10506 (
            .O(N__47735),
            .I(n15522));
    LocalMux I__10505 (
            .O(N__47732),
            .I(n15522));
    InMux I__10504 (
            .O(N__47727),
            .I(N__47724));
    LocalMux I__10503 (
            .O(N__47724),
            .I(N__47721));
    Span4Mux_h I__10502 (
            .O(N__47721),
            .I(N__47718));
    Odrv4 I__10501 (
            .O(N__47718),
            .I(n13));
    CascadeMux I__10500 (
            .O(N__47715),
            .I(N__47712));
    InMux I__10499 (
            .O(N__47712),
            .I(N__47708));
    CascadeMux I__10498 (
            .O(N__47711),
            .I(N__47704));
    LocalMux I__10497 (
            .O(N__47708),
            .I(N__47701));
    InMux I__10496 (
            .O(N__47707),
            .I(N__47698));
    InMux I__10495 (
            .O(N__47704),
            .I(N__47695));
    Span4Mux_v I__10494 (
            .O(N__47701),
            .I(N__47692));
    LocalMux I__10493 (
            .O(N__47698),
            .I(N__47689));
    LocalMux I__10492 (
            .O(N__47695),
            .I(encoder0_position_20));
    Odrv4 I__10491 (
            .O(N__47692),
            .I(encoder0_position_20));
    Odrv4 I__10490 (
            .O(N__47689),
            .I(encoder0_position_20));
    CascadeMux I__10489 (
            .O(N__47682),
            .I(N__47678));
    InMux I__10488 (
            .O(N__47681),
            .I(N__47675));
    InMux I__10487 (
            .O(N__47678),
            .I(N__47672));
    LocalMux I__10486 (
            .O(N__47675),
            .I(N__47669));
    LocalMux I__10485 (
            .O(N__47672),
            .I(n1125));
    Odrv4 I__10484 (
            .O(N__47669),
            .I(n1125));
    CascadeMux I__10483 (
            .O(N__47664),
            .I(n20_adj_618_cascade_));
    InMux I__10482 (
            .O(N__47661),
            .I(N__47658));
    LocalMux I__10481 (
            .O(N__47658),
            .I(N__47655));
    Odrv4 I__10480 (
            .O(N__47655),
            .I(n13197));
    CascadeMux I__10479 (
            .O(N__47652),
            .I(n1233_cascade_));
    InMux I__10478 (
            .O(N__47649),
            .I(N__47644));
    InMux I__10477 (
            .O(N__47648),
            .I(N__47641));
    InMux I__10476 (
            .O(N__47647),
            .I(N__47638));
    LocalMux I__10475 (
            .O(N__47644),
            .I(N__47631));
    LocalMux I__10474 (
            .O(N__47641),
            .I(N__47631));
    LocalMux I__10473 (
            .O(N__47638),
            .I(N__47631));
    Span4Mux_v I__10472 (
            .O(N__47631),
            .I(N__47628));
    Odrv4 I__10471 (
            .O(N__47628),
            .I(n297));
    InMux I__10470 (
            .O(N__47625),
            .I(N__47622));
    LocalMux I__10469 (
            .O(N__47622),
            .I(n1201));
    InMux I__10468 (
            .O(N__47619),
            .I(bfn_14_23_0_));
    CascadeMux I__10467 (
            .O(N__47616),
            .I(N__47612));
    InMux I__10466 (
            .O(N__47615),
            .I(N__47608));
    InMux I__10465 (
            .O(N__47612),
            .I(N__47605));
    InMux I__10464 (
            .O(N__47611),
            .I(N__47602));
    LocalMux I__10463 (
            .O(N__47608),
            .I(n1133));
    LocalMux I__10462 (
            .O(N__47605),
            .I(n1133));
    LocalMux I__10461 (
            .O(N__47602),
            .I(n1133));
    CascadeMux I__10460 (
            .O(N__47595),
            .I(N__47592));
    InMux I__10459 (
            .O(N__47592),
            .I(N__47589));
    LocalMux I__10458 (
            .O(N__47589),
            .I(n1200));
    InMux I__10457 (
            .O(N__47586),
            .I(n12522));
    InMux I__10456 (
            .O(N__47583),
            .I(n12523));
    CascadeMux I__10455 (
            .O(N__47580),
            .I(N__47576));
    CascadeMux I__10454 (
            .O(N__47579),
            .I(N__47573));
    InMux I__10453 (
            .O(N__47576),
            .I(N__47569));
    InMux I__10452 (
            .O(N__47573),
            .I(N__47566));
    InMux I__10451 (
            .O(N__47572),
            .I(N__47563));
    LocalMux I__10450 (
            .O(N__47569),
            .I(n1131));
    LocalMux I__10449 (
            .O(N__47566),
            .I(n1131));
    LocalMux I__10448 (
            .O(N__47563),
            .I(n1131));
    InMux I__10447 (
            .O(N__47556),
            .I(N__47553));
    LocalMux I__10446 (
            .O(N__47553),
            .I(N__47550));
    Odrv4 I__10445 (
            .O(N__47550),
            .I(n1198));
    InMux I__10444 (
            .O(N__47547),
            .I(n12524));
    CascadeMux I__10443 (
            .O(N__47544),
            .I(N__47540));
    CascadeMux I__10442 (
            .O(N__47543),
            .I(N__47537));
    InMux I__10441 (
            .O(N__47540),
            .I(N__47533));
    InMux I__10440 (
            .O(N__47537),
            .I(N__47530));
    InMux I__10439 (
            .O(N__47536),
            .I(N__47527));
    LocalMux I__10438 (
            .O(N__47533),
            .I(n1130));
    LocalMux I__10437 (
            .O(N__47530),
            .I(n1130));
    LocalMux I__10436 (
            .O(N__47527),
            .I(n1130));
    InMux I__10435 (
            .O(N__47520),
            .I(N__47517));
    LocalMux I__10434 (
            .O(N__47517),
            .I(n1197));
    InMux I__10433 (
            .O(N__47514),
            .I(n12525));
    InMux I__10432 (
            .O(N__47511),
            .I(n12526));
    InMux I__10431 (
            .O(N__47508),
            .I(n12550));
    InMux I__10430 (
            .O(N__47505),
            .I(n12551));
    InMux I__10429 (
            .O(N__47502),
            .I(N__47499));
    LocalMux I__10428 (
            .O(N__47499),
            .I(N__47496));
    Span4Mux_h I__10427 (
            .O(N__47496),
            .I(N__47493));
    Span4Mux_h I__10426 (
            .O(N__47493),
            .I(N__47490));
    Span4Mux_v I__10425 (
            .O(N__47490),
            .I(N__47486));
    InMux I__10424 (
            .O(N__47489),
            .I(N__47483));
    Odrv4 I__10423 (
            .O(N__47486),
            .I(n15553));
    LocalMux I__10422 (
            .O(N__47483),
            .I(n15553));
    CascadeMux I__10421 (
            .O(N__47478),
            .I(N__47475));
    InMux I__10420 (
            .O(N__47475),
            .I(N__47472));
    LocalMux I__10419 (
            .O(N__47472),
            .I(n1401));
    InMux I__10418 (
            .O(N__47469),
            .I(N__47466));
    LocalMux I__10417 (
            .O(N__47466),
            .I(n12019));
    CascadeMux I__10416 (
            .O(N__47463),
            .I(n14406_cascade_));
    InMux I__10415 (
            .O(N__47460),
            .I(N__47457));
    LocalMux I__10414 (
            .O(N__47457),
            .I(n14464));
    InMux I__10413 (
            .O(N__47454),
            .I(n12542));
    InMux I__10412 (
            .O(N__47451),
            .I(n12543));
    InMux I__10411 (
            .O(N__47448),
            .I(n12544));
    InMux I__10410 (
            .O(N__47445),
            .I(N__47442));
    LocalMux I__10409 (
            .O(N__47442),
            .I(n1396));
    InMux I__10408 (
            .O(N__47439),
            .I(n12545));
    InMux I__10407 (
            .O(N__47436),
            .I(N__47433));
    LocalMux I__10406 (
            .O(N__47433),
            .I(n1395));
    InMux I__10405 (
            .O(N__47430),
            .I(n12546));
    InMux I__10404 (
            .O(N__47427),
            .I(n12547));
    InMux I__10403 (
            .O(N__47424),
            .I(bfn_14_21_0_));
    InMux I__10402 (
            .O(N__47421),
            .I(N__47418));
    LocalMux I__10401 (
            .O(N__47418),
            .I(N__47415));
    Odrv4 I__10400 (
            .O(N__47415),
            .I(n1392));
    InMux I__10399 (
            .O(N__47412),
            .I(n12549));
    CascadeMux I__10398 (
            .O(N__47409),
            .I(n1427_cascade_));
    InMux I__10397 (
            .O(N__47406),
            .I(N__47402));
    InMux I__10396 (
            .O(N__47405),
            .I(N__47398));
    LocalMux I__10395 (
            .O(N__47402),
            .I(N__47395));
    InMux I__10394 (
            .O(N__47401),
            .I(N__47392));
    LocalMux I__10393 (
            .O(N__47398),
            .I(n1628_adj_608));
    Odrv4 I__10392 (
            .O(N__47395),
            .I(n1628_adj_608));
    LocalMux I__10391 (
            .O(N__47392),
            .I(n1628_adj_608));
    InMux I__10390 (
            .O(N__47385),
            .I(N__47382));
    LocalMux I__10389 (
            .O(N__47382),
            .I(N__47379));
    Span4Mux_v I__10388 (
            .O(N__47379),
            .I(N__47376));
    Span4Mux_h I__10387 (
            .O(N__47376),
            .I(N__47373));
    Odrv4 I__10386 (
            .O(N__47373),
            .I(n11));
    InMux I__10385 (
            .O(N__47370),
            .I(N__47366));
    CascadeMux I__10384 (
            .O(N__47369),
            .I(N__47362));
    LocalMux I__10383 (
            .O(N__47366),
            .I(N__47359));
    InMux I__10382 (
            .O(N__47365),
            .I(N__47356));
    InMux I__10381 (
            .O(N__47362),
            .I(N__47353));
    Span4Mux_h I__10380 (
            .O(N__47359),
            .I(N__47350));
    LocalMux I__10379 (
            .O(N__47356),
            .I(N__47347));
    LocalMux I__10378 (
            .O(N__47353),
            .I(encoder0_position_22));
    Odrv4 I__10377 (
            .O(N__47350),
            .I(encoder0_position_22));
    Odrv12 I__10376 (
            .O(N__47347),
            .I(encoder0_position_22));
    CascadeMux I__10375 (
            .O(N__47340),
            .I(N__47337));
    InMux I__10374 (
            .O(N__47337),
            .I(N__47332));
    InMux I__10373 (
            .O(N__47336),
            .I(N__47327));
    InMux I__10372 (
            .O(N__47335),
            .I(N__47327));
    LocalMux I__10371 (
            .O(N__47332),
            .I(n1626_adj_606));
    LocalMux I__10370 (
            .O(N__47327),
            .I(n1626_adj_606));
    InMux I__10369 (
            .O(N__47322),
            .I(N__47318));
    InMux I__10368 (
            .O(N__47321),
            .I(N__47315));
    LocalMux I__10367 (
            .O(N__47318),
            .I(N__47312));
    LocalMux I__10366 (
            .O(N__47315),
            .I(N__47309));
    Span12Mux_h I__10365 (
            .O(N__47312),
            .I(N__47306));
    Odrv4 I__10364 (
            .O(N__47309),
            .I(duty_6));
    Odrv12 I__10363 (
            .O(N__47306),
            .I(duty_6));
    InMux I__10362 (
            .O(N__47301),
            .I(N__47298));
    LocalMux I__10361 (
            .O(N__47298),
            .I(N__47295));
    Span12Mux_h I__10360 (
            .O(N__47295),
            .I(N__47292));
    Odrv12 I__10359 (
            .O(N__47292),
            .I(n19_adj_591));
    InMux I__10358 (
            .O(N__47289),
            .I(bfn_14_20_0_));
    InMux I__10357 (
            .O(N__47286),
            .I(n12541));
    CascadeMux I__10356 (
            .O(N__47283),
            .I(N__47280));
    InMux I__10355 (
            .O(N__47280),
            .I(N__47277));
    LocalMux I__10354 (
            .O(N__47277),
            .I(N__47273));
    CascadeMux I__10353 (
            .O(N__47276),
            .I(N__47270));
    Span4Mux_h I__10352 (
            .O(N__47273),
            .I(N__47267));
    InMux I__10351 (
            .O(N__47270),
            .I(N__47264));
    Odrv4 I__10350 (
            .O(N__47267),
            .I(n1624_adj_604));
    LocalMux I__10349 (
            .O(N__47264),
            .I(n1624_adj_604));
    InMux I__10348 (
            .O(N__47259),
            .I(N__47256));
    LocalMux I__10347 (
            .O(N__47256),
            .I(n14502));
    InMux I__10346 (
            .O(N__47253),
            .I(N__47250));
    LocalMux I__10345 (
            .O(N__47250),
            .I(N__47247));
    Span4Mux_h I__10344 (
            .O(N__47247),
            .I(N__47242));
    InMux I__10343 (
            .O(N__47246),
            .I(N__47239));
    InMux I__10342 (
            .O(N__47245),
            .I(N__47236));
    Odrv4 I__10341 (
            .O(N__47242),
            .I(n1623_adj_603));
    LocalMux I__10340 (
            .O(N__47239),
            .I(n1623_adj_603));
    LocalMux I__10339 (
            .O(N__47236),
            .I(n1623_adj_603));
    CascadeMux I__10338 (
            .O(N__47229),
            .I(n1624_adj_604_cascade_));
    InMux I__10337 (
            .O(N__47226),
            .I(N__47223));
    LocalMux I__10336 (
            .O(N__47223),
            .I(n13748));
    CascadeMux I__10335 (
            .O(N__47220),
            .I(N__47217));
    InMux I__10334 (
            .O(N__47217),
            .I(N__47214));
    LocalMux I__10333 (
            .O(N__47214),
            .I(n14508));
    CascadeMux I__10332 (
            .O(N__47211),
            .I(N__47208));
    InMux I__10331 (
            .O(N__47208),
            .I(N__47204));
    CascadeMux I__10330 (
            .O(N__47207),
            .I(N__47201));
    LocalMux I__10329 (
            .O(N__47204),
            .I(N__47197));
    InMux I__10328 (
            .O(N__47201),
            .I(N__47194));
    InMux I__10327 (
            .O(N__47200),
            .I(N__47191));
    Odrv4 I__10326 (
            .O(N__47197),
            .I(n1627_adj_607));
    LocalMux I__10325 (
            .O(N__47194),
            .I(n1627_adj_607));
    LocalMux I__10324 (
            .O(N__47191),
            .I(n1627_adj_607));
    CascadeMux I__10323 (
            .O(N__47184),
            .I(n1523_cascade_));
    InMux I__10322 (
            .O(N__47181),
            .I(N__47177));
    CascadeMux I__10321 (
            .O(N__47180),
            .I(N__47174));
    LocalMux I__10320 (
            .O(N__47177),
            .I(N__47170));
    InMux I__10319 (
            .O(N__47174),
            .I(N__47167));
    InMux I__10318 (
            .O(N__47173),
            .I(N__47164));
    Odrv4 I__10317 (
            .O(N__47170),
            .I(n1622_adj_602));
    LocalMux I__10316 (
            .O(N__47167),
            .I(n1622_adj_602));
    LocalMux I__10315 (
            .O(N__47164),
            .I(n1622_adj_602));
    InMux I__10314 (
            .O(N__47157),
            .I(N__47154));
    LocalMux I__10313 (
            .O(N__47154),
            .I(n14426));
    CascadeMux I__10312 (
            .O(N__47151),
            .I(n14428_cascade_));
    CascadeMux I__10311 (
            .O(N__47148),
            .I(n1554_cascade_));
    CascadeMux I__10310 (
            .O(N__47145),
            .I(N__47141));
    InMux I__10309 (
            .O(N__47144),
            .I(N__47138));
    InMux I__10308 (
            .O(N__47141),
            .I(N__47135));
    LocalMux I__10307 (
            .O(N__47138),
            .I(N__47132));
    LocalMux I__10306 (
            .O(N__47135),
            .I(N__47129));
    Span4Mux_h I__10305 (
            .O(N__47132),
            .I(N__47126));
    Span4Mux_h I__10304 (
            .O(N__47129),
            .I(N__47123));
    Odrv4 I__10303 (
            .O(N__47126),
            .I(n21_adj_667));
    Odrv4 I__10302 (
            .O(N__47123),
            .I(n21_adj_667));
    InMux I__10301 (
            .O(N__47118),
            .I(N__47112));
    InMux I__10300 (
            .O(N__47117),
            .I(N__47112));
    LocalMux I__10299 (
            .O(N__47112),
            .I(N__47109));
    Odrv4 I__10298 (
            .O(N__47109),
            .I(pwm_setpoint_10));
    CascadeMux I__10297 (
            .O(N__47106),
            .I(n21_adj_667_cascade_));
    InMux I__10296 (
            .O(N__47103),
            .I(N__47100));
    LocalMux I__10295 (
            .O(N__47100),
            .I(N__47097));
    Odrv12 I__10294 (
            .O(N__47097),
            .I(n6_adj_656));
    InMux I__10293 (
            .O(N__47094),
            .I(N__47091));
    LocalMux I__10292 (
            .O(N__47091),
            .I(N__47088));
    Odrv4 I__10291 (
            .O(N__47088),
            .I(n15203));
    CascadeMux I__10290 (
            .O(N__47085),
            .I(n14420_cascade_));
    InMux I__10289 (
            .O(N__47082),
            .I(N__47078));
    CascadeMux I__10288 (
            .O(N__47081),
            .I(N__47075));
    LocalMux I__10287 (
            .O(N__47078),
            .I(N__47072));
    InMux I__10286 (
            .O(N__47075),
            .I(N__47069));
    Odrv4 I__10285 (
            .O(N__47072),
            .I(n1630_adj_610));
    LocalMux I__10284 (
            .O(N__47069),
            .I(n1630_adj_610));
    InMux I__10283 (
            .O(N__47064),
            .I(N__47060));
    CascadeMux I__10282 (
            .O(N__47063),
            .I(N__47057));
    LocalMux I__10281 (
            .O(N__47060),
            .I(N__47053));
    InMux I__10280 (
            .O(N__47057),
            .I(N__47050));
    InMux I__10279 (
            .O(N__47056),
            .I(N__47047));
    Odrv4 I__10278 (
            .O(N__47053),
            .I(n1629_adj_609));
    LocalMux I__10277 (
            .O(N__47050),
            .I(n1629_adj_609));
    LocalMux I__10276 (
            .O(N__47047),
            .I(n1629_adj_609));
    CascadeMux I__10275 (
            .O(N__47040),
            .I(n1630_adj_610_cascade_));
    InMux I__10274 (
            .O(N__47037),
            .I(N__47034));
    LocalMux I__10273 (
            .O(N__47034),
            .I(\PWM.n17 ));
    CascadeMux I__10272 (
            .O(N__47031),
            .I(\PWM.n26_cascade_ ));
    InMux I__10271 (
            .O(N__47028),
            .I(N__47025));
    LocalMux I__10270 (
            .O(N__47025),
            .I(\PWM.n27 ));
    CascadeMux I__10269 (
            .O(N__47022),
            .I(\PWM.n29_cascade_ ));
    InMux I__10268 (
            .O(N__47019),
            .I(N__47016));
    LocalMux I__10267 (
            .O(N__47016),
            .I(\PWM.n28 ));
    InMux I__10266 (
            .O(N__47013),
            .I(N__47010));
    LocalMux I__10265 (
            .O(N__47010),
            .I(commutation_state_prev_2));
    InMux I__10264 (
            .O(N__47007),
            .I(N__47001));
    InMux I__10263 (
            .O(N__47006),
            .I(N__46997));
    InMux I__10262 (
            .O(N__47005),
            .I(N__46992));
    InMux I__10261 (
            .O(N__47004),
            .I(N__46992));
    LocalMux I__10260 (
            .O(N__47001),
            .I(N__46989));
    InMux I__10259 (
            .O(N__47000),
            .I(N__46985));
    LocalMux I__10258 (
            .O(N__46997),
            .I(N__46980));
    LocalMux I__10257 (
            .O(N__46992),
            .I(N__46980));
    Span4Mux_h I__10256 (
            .O(N__46989),
            .I(N__46977));
    InMux I__10255 (
            .O(N__46988),
            .I(N__46974));
    LocalMux I__10254 (
            .O(N__46985),
            .I(N__46971));
    Span4Mux_h I__10253 (
            .O(N__46980),
            .I(N__46968));
    Odrv4 I__10252 (
            .O(N__46977),
            .I(h2));
    LocalMux I__10251 (
            .O(N__46974),
            .I(h2));
    Odrv4 I__10250 (
            .O(N__46971),
            .I(h2));
    Odrv4 I__10249 (
            .O(N__46968),
            .I(h2));
    InMux I__10248 (
            .O(N__46959),
            .I(N__46952));
    InMux I__10247 (
            .O(N__46958),
            .I(N__46949));
    InMux I__10246 (
            .O(N__46957),
            .I(N__46944));
    InMux I__10245 (
            .O(N__46956),
            .I(N__46944));
    InMux I__10244 (
            .O(N__46955),
            .I(N__46941));
    LocalMux I__10243 (
            .O(N__46952),
            .I(N__46934));
    LocalMux I__10242 (
            .O(N__46949),
            .I(N__46934));
    LocalMux I__10241 (
            .O(N__46944),
            .I(N__46934));
    LocalMux I__10240 (
            .O(N__46941),
            .I(N__46931));
    Sp12to4 I__10239 (
            .O(N__46934),
            .I(N__46928));
    Sp12to4 I__10238 (
            .O(N__46931),
            .I(N__46924));
    Span12Mux_s10_v I__10237 (
            .O(N__46928),
            .I(N__46921));
    InMux I__10236 (
            .O(N__46927),
            .I(N__46918));
    Span12Mux_s6_v I__10235 (
            .O(N__46924),
            .I(N__46915));
    Span12Mux_h I__10234 (
            .O(N__46921),
            .I(N__46912));
    LocalMux I__10233 (
            .O(N__46918),
            .I(h3));
    Odrv12 I__10232 (
            .O(N__46915),
            .I(h3));
    Odrv12 I__10231 (
            .O(N__46912),
            .I(h3));
    CascadeMux I__10230 (
            .O(N__46905),
            .I(N__46900));
    CascadeMux I__10229 (
            .O(N__46904),
            .I(N__46896));
    InMux I__10228 (
            .O(N__46903),
            .I(N__46893));
    InMux I__10227 (
            .O(N__46900),
            .I(N__46887));
    InMux I__10226 (
            .O(N__46899),
            .I(N__46887));
    InMux I__10225 (
            .O(N__46896),
            .I(N__46884));
    LocalMux I__10224 (
            .O(N__46893),
            .I(N__46881));
    InMux I__10223 (
            .O(N__46892),
            .I(N__46878));
    LocalMux I__10222 (
            .O(N__46887),
            .I(N__46875));
    LocalMux I__10221 (
            .O(N__46884),
            .I(N__46870));
    Span4Mux_s2_v I__10220 (
            .O(N__46881),
            .I(N__46870));
    LocalMux I__10219 (
            .O(N__46878),
            .I(N__46867));
    Span4Mux_s2_v I__10218 (
            .O(N__46875),
            .I(N__46863));
    Span4Mux_h I__10217 (
            .O(N__46870),
            .I(N__46858));
    Span4Mux_s2_v I__10216 (
            .O(N__46867),
            .I(N__46858));
    InMux I__10215 (
            .O(N__46866),
            .I(N__46855));
    Sp12to4 I__10214 (
            .O(N__46863),
            .I(N__46850));
    Sp12to4 I__10213 (
            .O(N__46858),
            .I(N__46850));
    LocalMux I__10212 (
            .O(N__46855),
            .I(h1));
    Odrv12 I__10211 (
            .O(N__46850),
            .I(h1));
    CEMux I__10210 (
            .O(N__46845),
            .I(N__46842));
    LocalMux I__10209 (
            .O(N__46842),
            .I(N__46839));
    Odrv12 I__10208 (
            .O(N__46839),
            .I(n6_adj_721));
    SRMux I__10207 (
            .O(N__46836),
            .I(N__46833));
    LocalMux I__10206 (
            .O(N__46833),
            .I(commutation_state_7__N_261));
    InMux I__10205 (
            .O(N__46830),
            .I(N__46826));
    InMux I__10204 (
            .O(N__46829),
            .I(N__46823));
    LocalMux I__10203 (
            .O(N__46826),
            .I(N__46818));
    LocalMux I__10202 (
            .O(N__46823),
            .I(N__46818));
    Span4Mux_s2_v I__10201 (
            .O(N__46818),
            .I(N__46815));
    Span4Mux_v I__10200 (
            .O(N__46815),
            .I(N__46812));
    Odrv4 I__10199 (
            .O(N__46812),
            .I(pwm_setpoint_5));
    InMux I__10198 (
            .O(N__46809),
            .I(N__46806));
    LocalMux I__10197 (
            .O(N__46806),
            .I(N__46802));
    CascadeMux I__10196 (
            .O(N__46805),
            .I(N__46799));
    Span4Mux_v I__10195 (
            .O(N__46802),
            .I(N__46796));
    InMux I__10194 (
            .O(N__46799),
            .I(N__46793));
    Odrv4 I__10193 (
            .O(N__46796),
            .I(n11_adj_660));
    LocalMux I__10192 (
            .O(N__46793),
            .I(n11_adj_660));
    InMux I__10191 (
            .O(N__46788),
            .I(N__46785));
    LocalMux I__10190 (
            .O(N__46785),
            .I(N__46781));
    InMux I__10189 (
            .O(N__46784),
            .I(N__46778));
    Span4Mux_s2_v I__10188 (
            .O(N__46781),
            .I(N__46775));
    LocalMux I__10187 (
            .O(N__46778),
            .I(pwm_setpoint_14));
    Odrv4 I__10186 (
            .O(N__46775),
            .I(pwm_setpoint_14));
    CascadeMux I__10185 (
            .O(N__46770),
            .I(N__46767));
    InMux I__10184 (
            .O(N__46767),
            .I(N__46760));
    InMux I__10183 (
            .O(N__46766),
            .I(N__46760));
    InMux I__10182 (
            .O(N__46765),
            .I(N__46757));
    LocalMux I__10181 (
            .O(N__46760),
            .I(n29_adj_672));
    LocalMux I__10180 (
            .O(N__46757),
            .I(n29_adj_672));
    CascadeMux I__10179 (
            .O(N__46752),
            .I(N__46749));
    InMux I__10178 (
            .O(N__46749),
            .I(N__46745));
    InMux I__10177 (
            .O(N__46748),
            .I(N__46742));
    LocalMux I__10176 (
            .O(N__46745),
            .I(duty_19));
    LocalMux I__10175 (
            .O(N__46742),
            .I(duty_19));
    InMux I__10174 (
            .O(N__46737),
            .I(N__46734));
    LocalMux I__10173 (
            .O(N__46734),
            .I(N__46731));
    Odrv4 I__10172 (
            .O(N__46731),
            .I(n6_adj_578));
    InMux I__10171 (
            .O(N__46728),
            .I(N__46725));
    LocalMux I__10170 (
            .O(N__46725),
            .I(\PWM.n13991 ));
    CascadeMux I__10169 (
            .O(N__46722),
            .I(N__46715));
    CascadeMux I__10168 (
            .O(N__46721),
            .I(N__46712));
    InMux I__10167 (
            .O(N__46720),
            .I(N__46699));
    InMux I__10166 (
            .O(N__46719),
            .I(N__46699));
    InMux I__10165 (
            .O(N__46718),
            .I(N__46699));
    InMux I__10164 (
            .O(N__46715),
            .I(N__46699));
    InMux I__10163 (
            .O(N__46712),
            .I(N__46699));
    InMux I__10162 (
            .O(N__46711),
            .I(N__46694));
    InMux I__10161 (
            .O(N__46710),
            .I(N__46694));
    LocalMux I__10160 (
            .O(N__46699),
            .I(N__46687));
    LocalMux I__10159 (
            .O(N__46694),
            .I(N__46687));
    InMux I__10158 (
            .O(N__46693),
            .I(N__46682));
    InMux I__10157 (
            .O(N__46692),
            .I(N__46682));
    Span4Mux_v I__10156 (
            .O(N__46687),
            .I(N__46677));
    LocalMux I__10155 (
            .O(N__46682),
            .I(N__46677));
    Span4Mux_h I__10154 (
            .O(N__46677),
            .I(N__46674));
    Odrv4 I__10153 (
            .O(N__46674),
            .I(n4_adj_599));
    InMux I__10152 (
            .O(N__46671),
            .I(N__46668));
    LocalMux I__10151 (
            .O(N__46668),
            .I(commutation_state_prev_1));
    InMux I__10150 (
            .O(N__46665),
            .I(N__46661));
    InMux I__10149 (
            .O(N__46664),
            .I(N__46655));
    LocalMux I__10148 (
            .O(N__46661),
            .I(N__46652));
    InMux I__10147 (
            .O(N__46660),
            .I(N__46649));
    InMux I__10146 (
            .O(N__46659),
            .I(N__46644));
    InMux I__10145 (
            .O(N__46658),
            .I(N__46644));
    LocalMux I__10144 (
            .O(N__46655),
            .I(N__46641));
    Span4Mux_v I__10143 (
            .O(N__46652),
            .I(N__46638));
    LocalMux I__10142 (
            .O(N__46649),
            .I(N__46633));
    LocalMux I__10141 (
            .O(N__46644),
            .I(N__46633));
    Span4Mux_v I__10140 (
            .O(N__46641),
            .I(N__46630));
    Odrv4 I__10139 (
            .O(N__46638),
            .I(n5137));
    Odrv4 I__10138 (
            .O(N__46633),
            .I(n5137));
    Odrv4 I__10137 (
            .O(N__46630),
            .I(n5137));
    InMux I__10136 (
            .O(N__46623),
            .I(N__46617));
    InMux I__10135 (
            .O(N__46622),
            .I(N__46617));
    LocalMux I__10134 (
            .O(N__46617),
            .I(N__46611));
    InMux I__10133 (
            .O(N__46616),
            .I(N__46608));
    InMux I__10132 (
            .O(N__46615),
            .I(N__46605));
    InMux I__10131 (
            .O(N__46614),
            .I(N__46602));
    Span4Mux_v I__10130 (
            .O(N__46611),
            .I(N__46598));
    LocalMux I__10129 (
            .O(N__46608),
            .I(N__46591));
    LocalMux I__10128 (
            .O(N__46605),
            .I(N__46591));
    LocalMux I__10127 (
            .O(N__46602),
            .I(N__46591));
    InMux I__10126 (
            .O(N__46601),
            .I(N__46588));
    Span4Mux_v I__10125 (
            .O(N__46598),
            .I(N__46583));
    Span4Mux_v I__10124 (
            .O(N__46591),
            .I(N__46583));
    LocalMux I__10123 (
            .O(N__46588),
            .I(dti));
    Odrv4 I__10122 (
            .O(N__46583),
            .I(dti));
    CascadeMux I__10121 (
            .O(N__46578),
            .I(n5201_cascade_));
    InMux I__10120 (
            .O(N__46575),
            .I(N__46572));
    LocalMux I__10119 (
            .O(N__46572),
            .I(N__46568));
    InMux I__10118 (
            .O(N__46571),
            .I(N__46565));
    Span4Mux_v I__10117 (
            .O(N__46568),
            .I(N__46562));
    LocalMux I__10116 (
            .O(N__46565),
            .I(N__46559));
    Sp12to4 I__10115 (
            .O(N__46562),
            .I(N__46556));
    Span4Mux_h I__10114 (
            .O(N__46559),
            .I(N__46553));
    Odrv12 I__10113 (
            .O(N__46556),
            .I(pwm_setpoint_13));
    Odrv4 I__10112 (
            .O(N__46553),
            .I(pwm_setpoint_13));
    InMux I__10111 (
            .O(N__46548),
            .I(N__46544));
    InMux I__10110 (
            .O(N__46547),
            .I(N__46541));
    LocalMux I__10109 (
            .O(N__46544),
            .I(N__46535));
    LocalMux I__10108 (
            .O(N__46541),
            .I(N__46535));
    InMux I__10107 (
            .O(N__46540),
            .I(N__46532));
    Odrv4 I__10106 (
            .O(N__46535),
            .I(n27_adj_671));
    LocalMux I__10105 (
            .O(N__46532),
            .I(n27_adj_671));
    InMux I__10104 (
            .O(N__46527),
            .I(N__46523));
    InMux I__10103 (
            .O(N__46526),
            .I(N__46520));
    LocalMux I__10102 (
            .O(N__46523),
            .I(N__46517));
    LocalMux I__10101 (
            .O(N__46520),
            .I(duty_2));
    Odrv4 I__10100 (
            .O(N__46517),
            .I(duty_2));
    InMux I__10099 (
            .O(N__46512),
            .I(N__46509));
    LocalMux I__10098 (
            .O(N__46509),
            .I(N__46506));
    Span4Mux_v I__10097 (
            .O(N__46506),
            .I(N__46503));
    Odrv4 I__10096 (
            .O(N__46503),
            .I(n23_adj_595));
    InMux I__10095 (
            .O(N__46500),
            .I(N__46496));
    InMux I__10094 (
            .O(N__46499),
            .I(N__46493));
    LocalMux I__10093 (
            .O(N__46496),
            .I(N__46490));
    LocalMux I__10092 (
            .O(N__46493),
            .I(duty_15));
    Odrv12 I__10091 (
            .O(N__46490),
            .I(duty_15));
    InMux I__10090 (
            .O(N__46485),
            .I(N__46482));
    LocalMux I__10089 (
            .O(N__46482),
            .I(N__46479));
    Odrv12 I__10088 (
            .O(N__46479),
            .I(pwm_setpoint_23_N_171_15));
    InMux I__10087 (
            .O(N__46476),
            .I(N__46470));
    InMux I__10086 (
            .O(N__46475),
            .I(N__46470));
    LocalMux I__10085 (
            .O(N__46470),
            .I(N__46467));
    Span4Mux_s2_v I__10084 (
            .O(N__46467),
            .I(N__46464));
    Odrv4 I__10083 (
            .O(N__46464),
            .I(pwm_setpoint_15));
    InMux I__10082 (
            .O(N__46461),
            .I(N__46458));
    LocalMux I__10081 (
            .O(N__46458),
            .I(N__46453));
    InMux I__10080 (
            .O(N__46457),
            .I(N__46450));
    InMux I__10079 (
            .O(N__46456),
            .I(N__46447));
    Span4Mux_v I__10078 (
            .O(N__46453),
            .I(N__46442));
    LocalMux I__10077 (
            .O(N__46450),
            .I(N__46442));
    LocalMux I__10076 (
            .O(N__46447),
            .I(N__46439));
    Span4Mux_h I__10075 (
            .O(N__46442),
            .I(N__46434));
    Span4Mux_h I__10074 (
            .O(N__46439),
            .I(N__46434));
    Span4Mux_h I__10073 (
            .O(N__46434),
            .I(N__46431));
    Odrv4 I__10072 (
            .O(N__46431),
            .I(\quad_counter0.a_new_0 ));
    InMux I__10071 (
            .O(N__46428),
            .I(N__46425));
    LocalMux I__10070 (
            .O(N__46425),
            .I(N__46421));
    InMux I__10069 (
            .O(N__46424),
            .I(N__46418));
    Span4Mux_h I__10068 (
            .O(N__46421),
            .I(N__46412));
    LocalMux I__10067 (
            .O(N__46418),
            .I(N__46412));
    InMux I__10066 (
            .O(N__46417),
            .I(N__46409));
    Span4Mux_v I__10065 (
            .O(N__46412),
            .I(N__46406));
    LocalMux I__10064 (
            .O(N__46409),
            .I(\quad_counter0.b_new_0 ));
    Odrv4 I__10063 (
            .O(N__46406),
            .I(\quad_counter0.b_new_0 ));
    CascadeMux I__10062 (
            .O(N__46401),
            .I(N__46397));
    InMux I__10061 (
            .O(N__46400),
            .I(N__46390));
    InMux I__10060 (
            .O(N__46397),
            .I(N__46387));
    InMux I__10059 (
            .O(N__46396),
            .I(N__46380));
    InMux I__10058 (
            .O(N__46395),
            .I(N__46380));
    InMux I__10057 (
            .O(N__46394),
            .I(N__46380));
    CascadeMux I__10056 (
            .O(N__46393),
            .I(N__46377));
    LocalMux I__10055 (
            .O(N__46390),
            .I(N__46372));
    LocalMux I__10054 (
            .O(N__46387),
            .I(N__46372));
    LocalMux I__10053 (
            .O(N__46380),
            .I(N__46369));
    InMux I__10052 (
            .O(N__46377),
            .I(N__46366));
    Span4Mux_v I__10051 (
            .O(N__46372),
            .I(N__46361));
    Span4Mux_v I__10050 (
            .O(N__46369),
            .I(N__46361));
    LocalMux I__10049 (
            .O(N__46366),
            .I(a_new_1));
    Odrv4 I__10048 (
            .O(N__46361),
            .I(a_new_1));
    InMux I__10047 (
            .O(N__46356),
            .I(N__46353));
    LocalMux I__10046 (
            .O(N__46353),
            .I(N__46350));
    Odrv12 I__10045 (
            .O(N__46350),
            .I(\quad_counter0.a_prev_N_543 ));
    CascadeMux I__10044 (
            .O(N__46347),
            .I(N__46344));
    InMux I__10043 (
            .O(N__46344),
            .I(N__46341));
    LocalMux I__10042 (
            .O(N__46341),
            .I(N__46337));
    InMux I__10041 (
            .O(N__46340),
            .I(N__46334));
    Span4Mux_v I__10040 (
            .O(N__46337),
            .I(N__46327));
    LocalMux I__10039 (
            .O(N__46334),
            .I(N__46327));
    InMux I__10038 (
            .O(N__46333),
            .I(N__46322));
    InMux I__10037 (
            .O(N__46332),
            .I(N__46322));
    Span4Mux_v I__10036 (
            .O(N__46327),
            .I(N__46319));
    LocalMux I__10035 (
            .O(N__46322),
            .I(N__46316));
    Span4Mux_h I__10034 (
            .O(N__46319),
            .I(N__46313));
    Odrv12 I__10033 (
            .O(N__46316),
            .I(\quad_counter0.b_new_1 ));
    Odrv4 I__10032 (
            .O(N__46313),
            .I(\quad_counter0.b_new_1 ));
    CascadeMux I__10031 (
            .O(N__46308),
            .I(N__46303));
    InMux I__10030 (
            .O(N__46307),
            .I(N__46300));
    InMux I__10029 (
            .O(N__46306),
            .I(N__46297));
    InMux I__10028 (
            .O(N__46303),
            .I(N__46294));
    LocalMux I__10027 (
            .O(N__46300),
            .I(N__46291));
    LocalMux I__10026 (
            .O(N__46297),
            .I(N__46288));
    LocalMux I__10025 (
            .O(N__46294),
            .I(\quad_counter0.debounce_cnt ));
    Odrv12 I__10024 (
            .O(N__46291),
            .I(\quad_counter0.debounce_cnt ));
    Odrv12 I__10023 (
            .O(N__46288),
            .I(\quad_counter0.debounce_cnt ));
    CascadeMux I__10022 (
            .O(N__46281),
            .I(\quad_counter0.a_prev_N_543_cascade_ ));
    InMux I__10021 (
            .O(N__46278),
            .I(N__46274));
    InMux I__10020 (
            .O(N__46277),
            .I(N__46271));
    LocalMux I__10019 (
            .O(N__46274),
            .I(N__46266));
    LocalMux I__10018 (
            .O(N__46271),
            .I(N__46263));
    InMux I__10017 (
            .O(N__46270),
            .I(N__46260));
    InMux I__10016 (
            .O(N__46269),
            .I(N__46257));
    Span4Mux_h I__10015 (
            .O(N__46266),
            .I(N__46254));
    Span4Mux_h I__10014 (
            .O(N__46263),
            .I(N__46251));
    LocalMux I__10013 (
            .O(N__46260),
            .I(N__46248));
    LocalMux I__10012 (
            .O(N__46257),
            .I(b_prev));
    Odrv4 I__10011 (
            .O(N__46254),
            .I(b_prev));
    Odrv4 I__10010 (
            .O(N__46251),
            .I(b_prev));
    Odrv12 I__10009 (
            .O(N__46248),
            .I(b_prev));
    CascadeMux I__10008 (
            .O(N__46239),
            .I(N__46236));
    InMux I__10007 (
            .O(N__46236),
            .I(N__46233));
    LocalMux I__10006 (
            .O(N__46233),
            .I(N__46230));
    Span4Mux_v I__10005 (
            .O(N__46230),
            .I(N__46227));
    Odrv4 I__10004 (
            .O(N__46227),
            .I(n15121));
    InMux I__10003 (
            .O(N__46224),
            .I(N__46221));
    LocalMux I__10002 (
            .O(N__46221),
            .I(N__46218));
    Span4Mux_h I__10001 (
            .O(N__46218),
            .I(N__46215));
    Odrv4 I__10000 (
            .O(N__46215),
            .I(pwm_setpoint_23_N_171_6));
    InMux I__9999 (
            .O(N__46212),
            .I(N__46209));
    LocalMux I__9998 (
            .O(N__46209),
            .I(N__46205));
    InMux I__9997 (
            .O(N__46208),
            .I(N__46202));
    Odrv4 I__9996 (
            .O(N__46205),
            .I(pwm_setpoint_6));
    LocalMux I__9995 (
            .O(N__46202),
            .I(pwm_setpoint_6));
    InMux I__9994 (
            .O(N__46197),
            .I(N__46191));
    InMux I__9993 (
            .O(N__46196),
            .I(N__46191));
    LocalMux I__9992 (
            .O(N__46191),
            .I(N__46188));
    Odrv4 I__9991 (
            .O(N__46188),
            .I(pwm_setpoint_2));
    InMux I__9990 (
            .O(N__46185),
            .I(N__46179));
    InMux I__9989 (
            .O(N__46184),
            .I(N__46179));
    LocalMux I__9988 (
            .O(N__46179),
            .I(N__46176));
    Odrv4 I__9987 (
            .O(N__46176),
            .I(pwm_setpoint_3));
    CascadeMux I__9986 (
            .O(N__46173),
            .I(n14034_cascade_));
    CascadeMux I__9985 (
            .O(N__46170),
            .I(n14116_cascade_));
    InMux I__9984 (
            .O(N__46167),
            .I(N__46164));
    LocalMux I__9983 (
            .O(N__46164),
            .I(n10_adj_598));
    InMux I__9982 (
            .O(N__46161),
            .I(N__46158));
    LocalMux I__9981 (
            .O(N__46158),
            .I(N__46155));
    Odrv4 I__9980 (
            .O(N__46155),
            .I(pwm_setpoint_23_N_171_2));
    InMux I__9979 (
            .O(N__46152),
            .I(N__46149));
    LocalMux I__9978 (
            .O(N__46149),
            .I(N__46146));
    Odrv4 I__9977 (
            .O(N__46146),
            .I(pwm_setpoint_23_N_171_3));
    InMux I__9976 (
            .O(N__46143),
            .I(N__46139));
    InMux I__9975 (
            .O(N__46142),
            .I(N__46136));
    LocalMux I__9974 (
            .O(N__46139),
            .I(duty_3));
    LocalMux I__9973 (
            .O(N__46136),
            .I(duty_3));
    CascadeMux I__9972 (
            .O(N__46131),
            .I(N__46128));
    InMux I__9971 (
            .O(N__46128),
            .I(N__46125));
    LocalMux I__9970 (
            .O(N__46125),
            .I(n10_adj_681));
    CascadeMux I__9969 (
            .O(N__46122),
            .I(n16_adj_710_cascade_));
    InMux I__9968 (
            .O(N__46119),
            .I(N__46116));
    LocalMux I__9967 (
            .O(N__46116),
            .I(N__46113));
    Odrv4 I__9966 (
            .O(N__46113),
            .I(n15_adj_711));
    InMux I__9965 (
            .O(N__46110),
            .I(n12509));
    CascadeMux I__9964 (
            .O(N__46107),
            .I(N__46104));
    InMux I__9963 (
            .O(N__46104),
            .I(N__46101));
    LocalMux I__9962 (
            .O(N__46101),
            .I(N__46097));
    InMux I__9961 (
            .O(N__46100),
            .I(N__46093));
    Span4Mux_v I__9960 (
            .O(N__46097),
            .I(N__46090));
    InMux I__9959 (
            .O(N__46096),
            .I(N__46087));
    LocalMux I__9958 (
            .O(N__46093),
            .I(n930));
    Odrv4 I__9957 (
            .O(N__46090),
            .I(n930));
    LocalMux I__9956 (
            .O(N__46087),
            .I(n930));
    InMux I__9955 (
            .O(N__46080),
            .I(N__46077));
    LocalMux I__9954 (
            .O(N__46077),
            .I(n997));
    InMux I__9953 (
            .O(N__46074),
            .I(n12510));
    CascadeMux I__9952 (
            .O(N__46071),
            .I(N__46068));
    InMux I__9951 (
            .O(N__46068),
            .I(N__46065));
    LocalMux I__9950 (
            .O(N__46065),
            .I(N__46061));
    InMux I__9949 (
            .O(N__46064),
            .I(N__46058));
    Span4Mux_h I__9948 (
            .O(N__46061),
            .I(N__46055));
    LocalMux I__9947 (
            .O(N__46058),
            .I(n929));
    Odrv4 I__9946 (
            .O(N__46055),
            .I(n929));
    InMux I__9945 (
            .O(N__46050),
            .I(N__46047));
    LocalMux I__9944 (
            .O(N__46047),
            .I(n996));
    InMux I__9943 (
            .O(N__46044),
            .I(n12511));
    CascadeMux I__9942 (
            .O(N__46041),
            .I(N__46038));
    InMux I__9941 (
            .O(N__46038),
            .I(N__46033));
    InMux I__9940 (
            .O(N__46037),
            .I(N__46028));
    InMux I__9939 (
            .O(N__46036),
            .I(N__46028));
    LocalMux I__9938 (
            .O(N__46033),
            .I(n928));
    LocalMux I__9937 (
            .O(N__46028),
            .I(n928));
    InMux I__9936 (
            .O(N__46023),
            .I(N__46020));
    LocalMux I__9935 (
            .O(N__46020),
            .I(n995));
    InMux I__9934 (
            .O(N__46017),
            .I(n12512));
    CascadeMux I__9933 (
            .O(N__46014),
            .I(N__46009));
    CascadeMux I__9932 (
            .O(N__46013),
            .I(N__46005));
    InMux I__9931 (
            .O(N__46012),
            .I(N__45999));
    InMux I__9930 (
            .O(N__46009),
            .I(N__45996));
    InMux I__9929 (
            .O(N__46008),
            .I(N__45993));
    InMux I__9928 (
            .O(N__46005),
            .I(N__45984));
    InMux I__9927 (
            .O(N__46004),
            .I(N__45984));
    InMux I__9926 (
            .O(N__46003),
            .I(N__45984));
    InMux I__9925 (
            .O(N__46002),
            .I(N__45984));
    LocalMux I__9924 (
            .O(N__45999),
            .I(n960));
    LocalMux I__9923 (
            .O(N__45996),
            .I(n960));
    LocalMux I__9922 (
            .O(N__45993),
            .I(n960));
    LocalMux I__9921 (
            .O(N__45984),
            .I(n960));
    CascadeMux I__9920 (
            .O(N__45975),
            .I(N__45972));
    InMux I__9919 (
            .O(N__45972),
            .I(N__45969));
    LocalMux I__9918 (
            .O(N__45969),
            .I(N__45965));
    InMux I__9917 (
            .O(N__45968),
            .I(N__45962));
    Odrv4 I__9916 (
            .O(N__45965),
            .I(n927));
    LocalMux I__9915 (
            .O(N__45962),
            .I(n927));
    InMux I__9914 (
            .O(N__45957),
            .I(n12513));
    InMux I__9913 (
            .O(N__45954),
            .I(N__45951));
    LocalMux I__9912 (
            .O(N__45951),
            .I(N__45948));
    Odrv12 I__9911 (
            .O(N__45948),
            .I(encoder0_position_scaled_0));
    InMux I__9910 (
            .O(N__45945),
            .I(N__45942));
    LocalMux I__9909 (
            .O(N__45942),
            .I(n25_adj_551));
    CascadeMux I__9908 (
            .O(N__45939),
            .I(n11872_cascade_));
    CascadeMux I__9907 (
            .O(N__45936),
            .I(n11933_cascade_));
    CascadeMux I__9906 (
            .O(N__45933),
            .I(n13728_cascade_));
    CascadeMux I__9905 (
            .O(N__45930),
            .I(n1059_cascade_));
    CascadeMux I__9904 (
            .O(N__45927),
            .I(n1132_cascade_));
    InMux I__9903 (
            .O(N__45924),
            .I(N__45920));
    InMux I__9902 (
            .O(N__45923),
            .I(N__45917));
    LocalMux I__9901 (
            .O(N__45920),
            .I(n295));
    LocalMux I__9900 (
            .O(N__45917),
            .I(n295));
    InMux I__9899 (
            .O(N__45912),
            .I(N__45909));
    LocalMux I__9898 (
            .O(N__45909),
            .I(n1001));
    InMux I__9897 (
            .O(N__45906),
            .I(bfn_13_24_0_));
    CascadeMux I__9896 (
            .O(N__45903),
            .I(N__45900));
    InMux I__9895 (
            .O(N__45900),
            .I(N__45896));
    InMux I__9894 (
            .O(N__45899),
            .I(N__45893));
    LocalMux I__9893 (
            .O(N__45896),
            .I(n933));
    LocalMux I__9892 (
            .O(N__45893),
            .I(n933));
    InMux I__9891 (
            .O(N__45888),
            .I(N__45885));
    LocalMux I__9890 (
            .O(N__45885),
            .I(n1000));
    InMux I__9889 (
            .O(N__45882),
            .I(n12507));
    CascadeMux I__9888 (
            .O(N__45879),
            .I(N__45876));
    InMux I__9887 (
            .O(N__45876),
            .I(N__45872));
    InMux I__9886 (
            .O(N__45875),
            .I(N__45869));
    LocalMux I__9885 (
            .O(N__45872),
            .I(n932));
    LocalMux I__9884 (
            .O(N__45869),
            .I(n932));
    InMux I__9883 (
            .O(N__45864),
            .I(N__45861));
    LocalMux I__9882 (
            .O(N__45861),
            .I(n999));
    InMux I__9881 (
            .O(N__45858),
            .I(n12508));
    CascadeMux I__9880 (
            .O(N__45855),
            .I(N__45851));
    InMux I__9879 (
            .O(N__45854),
            .I(N__45847));
    InMux I__9878 (
            .O(N__45851),
            .I(N__45844));
    InMux I__9877 (
            .O(N__45850),
            .I(N__45841));
    LocalMux I__9876 (
            .O(N__45847),
            .I(n931));
    LocalMux I__9875 (
            .O(N__45844),
            .I(n931));
    LocalMux I__9874 (
            .O(N__45841),
            .I(n931));
    CascadeMux I__9873 (
            .O(N__45834),
            .I(N__45831));
    InMux I__9872 (
            .O(N__45831),
            .I(N__45828));
    LocalMux I__9871 (
            .O(N__45828),
            .I(N__45825));
    Odrv4 I__9870 (
            .O(N__45825),
            .I(n998));
    InMux I__9869 (
            .O(N__45822),
            .I(N__45819));
    LocalMux I__9868 (
            .O(N__45819),
            .I(N__45816));
    Span4Mux_v I__9867 (
            .O(N__45816),
            .I(N__45813));
    Span4Mux_h I__9866 (
            .O(N__45813),
            .I(N__45810));
    Sp12to4 I__9865 (
            .O(N__45810),
            .I(N__45807));
    Odrv12 I__9864 (
            .O(N__45807),
            .I(ENCODER0_B_N));
    InMux I__9863 (
            .O(N__45804),
            .I(N__45801));
    LocalMux I__9862 (
            .O(N__45801),
            .I(N__45796));
    InMux I__9861 (
            .O(N__45800),
            .I(N__45793));
    CascadeMux I__9860 (
            .O(N__45799),
            .I(N__45790));
    Span4Mux_h I__9859 (
            .O(N__45796),
            .I(N__45787));
    LocalMux I__9858 (
            .O(N__45793),
            .I(N__45784));
    InMux I__9857 (
            .O(N__45790),
            .I(N__45781));
    Span4Mux_v I__9856 (
            .O(N__45787),
            .I(N__45776));
    Span4Mux_v I__9855 (
            .O(N__45784),
            .I(N__45776));
    LocalMux I__9854 (
            .O(N__45781),
            .I(encoder0_position_1));
    Odrv4 I__9853 (
            .O(N__45776),
            .I(encoder0_position_1));
    CascadeMux I__9852 (
            .O(N__45771),
            .I(N__45768));
    InMux I__9851 (
            .O(N__45768),
            .I(N__45765));
    LocalMux I__9850 (
            .O(N__45765),
            .I(N__45762));
    Odrv12 I__9849 (
            .O(N__45762),
            .I(n32_adj_650));
    InMux I__9848 (
            .O(N__45759),
            .I(N__45754));
    InMux I__9847 (
            .O(N__45758),
            .I(N__45751));
    CascadeMux I__9846 (
            .O(N__45757),
            .I(N__45748));
    LocalMux I__9845 (
            .O(N__45754),
            .I(N__45743));
    LocalMux I__9844 (
            .O(N__45751),
            .I(N__45743));
    InMux I__9843 (
            .O(N__45748),
            .I(N__45740));
    Span4Mux_h I__9842 (
            .O(N__45743),
            .I(N__45737));
    LocalMux I__9841 (
            .O(N__45740),
            .I(encoder0_position_16));
    Odrv4 I__9840 (
            .O(N__45737),
            .I(encoder0_position_16));
    CascadeMux I__9839 (
            .O(N__45732),
            .I(N__45729));
    InMux I__9838 (
            .O(N__45729),
            .I(N__45726));
    LocalMux I__9837 (
            .O(N__45726),
            .I(N__45723));
    Span4Mux_v I__9836 (
            .O(N__45723),
            .I(N__45720));
    Odrv4 I__9835 (
            .O(N__45720),
            .I(n17_adj_635));
    CascadeMux I__9834 (
            .O(N__45717),
            .I(n1129_cascade_));
    CascadeMux I__9833 (
            .O(N__45714),
            .I(n1625_adj_605_cascade_));
    InMux I__9832 (
            .O(N__45711),
            .I(N__45708));
    LocalMux I__9831 (
            .O(N__45708),
            .I(N__45705));
    Odrv4 I__9830 (
            .O(N__45705),
            .I(n1698));
    InMux I__9829 (
            .O(N__45702),
            .I(N__45698));
    CascadeMux I__9828 (
            .O(N__45701),
            .I(N__45695));
    LocalMux I__9827 (
            .O(N__45698),
            .I(N__45692));
    InMux I__9826 (
            .O(N__45695),
            .I(N__45689));
    Odrv4 I__9825 (
            .O(N__45692),
            .I(n1730));
    LocalMux I__9824 (
            .O(N__45689),
            .I(n1730));
    CascadeMux I__9823 (
            .O(N__45684),
            .I(n1730_cascade_));
    CascadeMux I__9822 (
            .O(N__45681),
            .I(N__45678));
    InMux I__9821 (
            .O(N__45678),
            .I(N__45674));
    CascadeMux I__9820 (
            .O(N__45677),
            .I(N__45671));
    LocalMux I__9819 (
            .O(N__45674),
            .I(N__45667));
    InMux I__9818 (
            .O(N__45671),
            .I(N__45664));
    InMux I__9817 (
            .O(N__45670),
            .I(N__45661));
    Odrv4 I__9816 (
            .O(N__45667),
            .I(n1729));
    LocalMux I__9815 (
            .O(N__45664),
            .I(n1729));
    LocalMux I__9814 (
            .O(N__45661),
            .I(n1729));
    InMux I__9813 (
            .O(N__45654),
            .I(N__45651));
    LocalMux I__9812 (
            .O(N__45651),
            .I(N__45648));
    Odrv4 I__9811 (
            .O(N__45648),
            .I(n14514));
    CascadeMux I__9810 (
            .O(N__45645),
            .I(N__45642));
    InMux I__9809 (
            .O(N__45642),
            .I(N__45639));
    LocalMux I__9808 (
            .O(N__45639),
            .I(N__45636));
    Span4Mux_v I__9807 (
            .O(N__45636),
            .I(N__45633));
    Odrv4 I__9806 (
            .O(N__45633),
            .I(n11_adj_629));
    InMux I__9805 (
            .O(N__45630),
            .I(N__45627));
    LocalMux I__9804 (
            .O(N__45627),
            .I(N__45624));
    Odrv12 I__9803 (
            .O(N__45624),
            .I(n1701));
    InMux I__9802 (
            .O(N__45621),
            .I(N__45618));
    LocalMux I__9801 (
            .O(N__45618),
            .I(N__45610));
    CascadeMux I__9800 (
            .O(N__45617),
            .I(N__45605));
    CascadeMux I__9799 (
            .O(N__45616),
            .I(N__45599));
    CascadeMux I__9798 (
            .O(N__45615),
            .I(N__45594));
    CascadeMux I__9797 (
            .O(N__45614),
            .I(N__45591));
    CascadeMux I__9796 (
            .O(N__45613),
            .I(N__45588));
    Span12Mux_h I__9795 (
            .O(N__45610),
            .I(N__45583));
    InMux I__9794 (
            .O(N__45609),
            .I(N__45578));
    InMux I__9793 (
            .O(N__45608),
            .I(N__45578));
    InMux I__9792 (
            .O(N__45605),
            .I(N__45575));
    InMux I__9791 (
            .O(N__45604),
            .I(N__45564));
    InMux I__9790 (
            .O(N__45603),
            .I(N__45564));
    InMux I__9789 (
            .O(N__45602),
            .I(N__45564));
    InMux I__9788 (
            .O(N__45599),
            .I(N__45564));
    InMux I__9787 (
            .O(N__45598),
            .I(N__45564));
    InMux I__9786 (
            .O(N__45597),
            .I(N__45559));
    InMux I__9785 (
            .O(N__45594),
            .I(N__45559));
    InMux I__9784 (
            .O(N__45591),
            .I(N__45550));
    InMux I__9783 (
            .O(N__45588),
            .I(N__45550));
    InMux I__9782 (
            .O(N__45587),
            .I(N__45550));
    InMux I__9781 (
            .O(N__45586),
            .I(N__45550));
    Odrv12 I__9780 (
            .O(N__45583),
            .I(n1653));
    LocalMux I__9779 (
            .O(N__45578),
            .I(n1653));
    LocalMux I__9778 (
            .O(N__45575),
            .I(n1653));
    LocalMux I__9777 (
            .O(N__45564),
            .I(n1653));
    LocalMux I__9776 (
            .O(N__45559),
            .I(n1653));
    LocalMux I__9775 (
            .O(N__45550),
            .I(n1653));
    InMux I__9774 (
            .O(N__45537),
            .I(N__45534));
    LocalMux I__9773 (
            .O(N__45534),
            .I(N__45530));
    CascadeMux I__9772 (
            .O(N__45533),
            .I(N__45527));
    Span4Mux_h I__9771 (
            .O(N__45530),
            .I(N__45523));
    InMux I__9770 (
            .O(N__45527),
            .I(N__45520));
    InMux I__9769 (
            .O(N__45526),
            .I(N__45517));
    Odrv4 I__9768 (
            .O(N__45523),
            .I(n1733));
    LocalMux I__9767 (
            .O(N__45520),
            .I(n1733));
    LocalMux I__9766 (
            .O(N__45517),
            .I(n1733));
    InMux I__9765 (
            .O(N__45510),
            .I(N__45507));
    LocalMux I__9764 (
            .O(N__45507),
            .I(N__45503));
    CascadeMux I__9763 (
            .O(N__45506),
            .I(N__45496));
    Span4Mux_v I__9762 (
            .O(N__45503),
            .I(N__45493));
    InMux I__9761 (
            .O(N__45502),
            .I(N__45490));
    CascadeMux I__9760 (
            .O(N__45501),
            .I(N__45487));
    InMux I__9759 (
            .O(N__45500),
            .I(N__45481));
    CascadeMux I__9758 (
            .O(N__45499),
            .I(N__45477));
    InMux I__9757 (
            .O(N__45496),
            .I(N__45473));
    Span4Mux_h I__9756 (
            .O(N__45493),
            .I(N__45468));
    LocalMux I__9755 (
            .O(N__45490),
            .I(N__45468));
    InMux I__9754 (
            .O(N__45487),
            .I(N__45465));
    CascadeMux I__9753 (
            .O(N__45486),
            .I(N__45462));
    CascadeMux I__9752 (
            .O(N__45485),
            .I(N__45458));
    InMux I__9751 (
            .O(N__45484),
            .I(N__45451));
    LocalMux I__9750 (
            .O(N__45481),
            .I(N__45448));
    InMux I__9749 (
            .O(N__45480),
            .I(N__45445));
    InMux I__9748 (
            .O(N__45477),
            .I(N__45440));
    InMux I__9747 (
            .O(N__45476),
            .I(N__45440));
    LocalMux I__9746 (
            .O(N__45473),
            .I(N__45433));
    Span4Mux_v I__9745 (
            .O(N__45468),
            .I(N__45433));
    LocalMux I__9744 (
            .O(N__45465),
            .I(N__45433));
    InMux I__9743 (
            .O(N__45462),
            .I(N__45422));
    InMux I__9742 (
            .O(N__45461),
            .I(N__45422));
    InMux I__9741 (
            .O(N__45458),
            .I(N__45422));
    InMux I__9740 (
            .O(N__45457),
            .I(N__45422));
    InMux I__9739 (
            .O(N__45456),
            .I(N__45422));
    InMux I__9738 (
            .O(N__45455),
            .I(N__45417));
    InMux I__9737 (
            .O(N__45454),
            .I(N__45417));
    LocalMux I__9736 (
            .O(N__45451),
            .I(N__45410));
    Span4Mux_h I__9735 (
            .O(N__45448),
            .I(N__45410));
    LocalMux I__9734 (
            .O(N__45445),
            .I(N__45410));
    LocalMux I__9733 (
            .O(N__45440),
            .I(n1752));
    Odrv4 I__9732 (
            .O(N__45433),
            .I(n1752));
    LocalMux I__9731 (
            .O(N__45422),
            .I(n1752));
    LocalMux I__9730 (
            .O(N__45417),
            .I(n1752));
    Odrv4 I__9729 (
            .O(N__45410),
            .I(n1752));
    InMux I__9728 (
            .O(N__45399),
            .I(N__45396));
    LocalMux I__9727 (
            .O(N__45396),
            .I(N__45393));
    Span4Mux_h I__9726 (
            .O(N__45393),
            .I(N__45390));
    Span4Mux_h I__9725 (
            .O(N__45390),
            .I(N__45386));
    CascadeMux I__9724 (
            .O(N__45389),
            .I(N__45383));
    Span4Mux_v I__9723 (
            .O(N__45386),
            .I(N__45380));
    InMux I__9722 (
            .O(N__45383),
            .I(N__45377));
    Odrv4 I__9721 (
            .O(N__45380),
            .I(n15630));
    LocalMux I__9720 (
            .O(N__45377),
            .I(n15630));
    CascadeMux I__9719 (
            .O(N__45372),
            .I(N__45368));
    InMux I__9718 (
            .O(N__45371),
            .I(N__45365));
    InMux I__9717 (
            .O(N__45368),
            .I(N__45361));
    LocalMux I__9716 (
            .O(N__45365),
            .I(N__45358));
    InMux I__9715 (
            .O(N__45364),
            .I(N__45355));
    LocalMux I__9714 (
            .O(N__45361),
            .I(n1621_adj_601));
    Odrv4 I__9713 (
            .O(N__45358),
            .I(n1621_adj_601));
    LocalMux I__9712 (
            .O(N__45355),
            .I(n1621_adj_601));
    InMux I__9711 (
            .O(N__45348),
            .I(n12590));
    InMux I__9710 (
            .O(N__45345),
            .I(N__45342));
    LocalMux I__9709 (
            .O(N__45342),
            .I(N__45338));
    CascadeMux I__9708 (
            .O(N__45341),
            .I(N__45335));
    Span4Mux_v I__9707 (
            .O(N__45338),
            .I(N__45332));
    InMux I__9706 (
            .O(N__45335),
            .I(N__45329));
    Odrv4 I__9705 (
            .O(N__45332),
            .I(n1719));
    LocalMux I__9704 (
            .O(N__45329),
            .I(n1719));
    InMux I__9703 (
            .O(N__45324),
            .I(N__45321));
    LocalMux I__9702 (
            .O(N__45321),
            .I(n1695));
    CascadeMux I__9701 (
            .O(N__45318),
            .I(N__45315));
    InMux I__9700 (
            .O(N__45315),
            .I(N__45311));
    InMux I__9699 (
            .O(N__45314),
            .I(N__45307));
    LocalMux I__9698 (
            .O(N__45311),
            .I(N__45304));
    InMux I__9697 (
            .O(N__45310),
            .I(N__45301));
    LocalMux I__9696 (
            .O(N__45307),
            .I(n1727));
    Odrv4 I__9695 (
            .O(N__45304),
            .I(n1727));
    LocalMux I__9694 (
            .O(N__45301),
            .I(n1727));
    InMux I__9693 (
            .O(N__45294),
            .I(N__45291));
    LocalMux I__9692 (
            .O(N__45291),
            .I(N__45288));
    Odrv4 I__9691 (
            .O(N__45288),
            .I(n1696));
    CascadeMux I__9690 (
            .O(N__45285),
            .I(n1653_cascade_));
    CascadeMux I__9689 (
            .O(N__45282),
            .I(N__45279));
    InMux I__9688 (
            .O(N__45279),
            .I(N__45274));
    InMux I__9687 (
            .O(N__45278),
            .I(N__45269));
    InMux I__9686 (
            .O(N__45277),
            .I(N__45269));
    LocalMux I__9685 (
            .O(N__45274),
            .I(n1728));
    LocalMux I__9684 (
            .O(N__45269),
            .I(n1728));
    CascadeMux I__9683 (
            .O(N__45264),
            .I(N__45261));
    InMux I__9682 (
            .O(N__45261),
            .I(N__45258));
    LocalMux I__9681 (
            .O(N__45258),
            .I(N__45255));
    Odrv4 I__9680 (
            .O(N__45255),
            .I(n1697));
    InMux I__9679 (
            .O(N__45252),
            .I(N__45249));
    LocalMux I__9678 (
            .O(N__45249),
            .I(n1692));
    CascadeMux I__9677 (
            .O(N__45246),
            .I(N__45242));
    InMux I__9676 (
            .O(N__45245),
            .I(N__45239));
    InMux I__9675 (
            .O(N__45242),
            .I(N__45236));
    LocalMux I__9674 (
            .O(N__45239),
            .I(N__45232));
    LocalMux I__9673 (
            .O(N__45236),
            .I(N__45229));
    InMux I__9672 (
            .O(N__45235),
            .I(N__45226));
    Odrv4 I__9671 (
            .O(N__45232),
            .I(n1724));
    Odrv4 I__9670 (
            .O(N__45229),
            .I(n1724));
    LocalMux I__9669 (
            .O(N__45226),
            .I(n1724));
    CascadeMux I__9668 (
            .O(N__45219),
            .I(N__45216));
    InMux I__9667 (
            .O(N__45216),
            .I(N__45213));
    LocalMux I__9666 (
            .O(N__45213),
            .I(n1693_adj_614));
    CascadeMux I__9665 (
            .O(N__45210),
            .I(N__45206));
    CascadeMux I__9664 (
            .O(N__45209),
            .I(N__45203));
    InMux I__9663 (
            .O(N__45206),
            .I(N__45200));
    InMux I__9662 (
            .O(N__45203),
            .I(N__45197));
    LocalMux I__9661 (
            .O(N__45200),
            .I(N__45193));
    LocalMux I__9660 (
            .O(N__45197),
            .I(N__45190));
    InMux I__9659 (
            .O(N__45196),
            .I(N__45187));
    Odrv4 I__9658 (
            .O(N__45193),
            .I(n1725));
    Odrv4 I__9657 (
            .O(N__45190),
            .I(n1725));
    LocalMux I__9656 (
            .O(N__45187),
            .I(n1725));
    InMux I__9655 (
            .O(N__45180),
            .I(N__45177));
    LocalMux I__9654 (
            .O(N__45177),
            .I(N__45174));
    Span4Mux_h I__9653 (
            .O(N__45174),
            .I(N__45171));
    Span4Mux_v I__9652 (
            .O(N__45171),
            .I(N__45168));
    Span4Mux_v I__9651 (
            .O(N__45168),
            .I(N__45164));
    InMux I__9650 (
            .O(N__45167),
            .I(N__45161));
    Odrv4 I__9649 (
            .O(N__45164),
            .I(n15611));
    LocalMux I__9648 (
            .O(N__45161),
            .I(n15611));
    CascadeMux I__9647 (
            .O(N__45156),
            .I(N__45152));
    InMux I__9646 (
            .O(N__45155),
            .I(N__45149));
    InMux I__9645 (
            .O(N__45152),
            .I(N__45146));
    LocalMux I__9644 (
            .O(N__45149),
            .I(n1625_adj_605));
    LocalMux I__9643 (
            .O(N__45146),
            .I(n1625_adj_605));
    InMux I__9642 (
            .O(N__45141),
            .I(n12581));
    InMux I__9641 (
            .O(N__45138),
            .I(n12582));
    InMux I__9640 (
            .O(N__45135),
            .I(N__45132));
    LocalMux I__9639 (
            .O(N__45132),
            .I(n1694));
    InMux I__9638 (
            .O(N__45129),
            .I(n12583));
    InMux I__9637 (
            .O(N__45126),
            .I(bfn_13_18_0_));
    InMux I__9636 (
            .O(N__45123),
            .I(n12585));
    InMux I__9635 (
            .O(N__45120),
            .I(N__45117));
    LocalMux I__9634 (
            .O(N__45117),
            .I(n1691));
    InMux I__9633 (
            .O(N__45114),
            .I(n12586));
    CascadeMux I__9632 (
            .O(N__45111),
            .I(N__45108));
    InMux I__9631 (
            .O(N__45108),
            .I(N__45105));
    LocalMux I__9630 (
            .O(N__45105),
            .I(n1690));
    InMux I__9629 (
            .O(N__45102),
            .I(n12587));
    CascadeMux I__9628 (
            .O(N__45099),
            .I(N__45096));
    InMux I__9627 (
            .O(N__45096),
            .I(N__45093));
    LocalMux I__9626 (
            .O(N__45093),
            .I(n1689));
    InMux I__9625 (
            .O(N__45090),
            .I(n12588));
    InMux I__9624 (
            .O(N__45087),
            .I(N__45084));
    LocalMux I__9623 (
            .O(N__45084),
            .I(n1688));
    InMux I__9622 (
            .O(N__45081),
            .I(n12589));
    InMux I__9621 (
            .O(N__45078),
            .I(N__45072));
    InMux I__9620 (
            .O(N__45077),
            .I(N__45072));
    LocalMux I__9619 (
            .O(N__45072),
            .I(n33_adj_675));
    CascadeMux I__9618 (
            .O(N__45069),
            .I(N__45066));
    InMux I__9617 (
            .O(N__45066),
            .I(N__45063));
    LocalMux I__9616 (
            .O(N__45063),
            .I(n15104));
    InMux I__9615 (
            .O(N__45060),
            .I(N__45054));
    InMux I__9614 (
            .O(N__45059),
            .I(N__45054));
    LocalMux I__9613 (
            .O(N__45054),
            .I(n31_adj_674));
    CascadeMux I__9612 (
            .O(N__45051),
            .I(N__45046));
    InMux I__9611 (
            .O(N__45050),
            .I(N__45039));
    InMux I__9610 (
            .O(N__45049),
            .I(N__45039));
    InMux I__9609 (
            .O(N__45046),
            .I(N__45039));
    LocalMux I__9608 (
            .O(N__45039),
            .I(n35));
    InMux I__9607 (
            .O(N__45036),
            .I(N__45033));
    LocalMux I__9606 (
            .O(N__45033),
            .I(n15247));
    CascadeMux I__9605 (
            .O(N__45030),
            .I(n15099_cascade_));
    InMux I__9604 (
            .O(N__45027),
            .I(N__45024));
    LocalMux I__9603 (
            .O(N__45024),
            .I(n15220));
    InMux I__9602 (
            .O(N__45021),
            .I(N__45015));
    InMux I__9601 (
            .O(N__45020),
            .I(N__45015));
    LocalMux I__9600 (
            .O(N__45015),
            .I(N__45012));
    Odrv4 I__9599 (
            .O(N__45012),
            .I(pwm_setpoint_18));
    CascadeMux I__9598 (
            .O(N__45009),
            .I(n15257_cascade_));
    InMux I__9597 (
            .O(N__45006),
            .I(N__45000));
    InMux I__9596 (
            .O(N__45005),
            .I(N__45000));
    LocalMux I__9595 (
            .O(N__45000),
            .I(n37));
    InMux I__9594 (
            .O(N__44997),
            .I(N__44994));
    LocalMux I__9593 (
            .O(N__44994),
            .I(N__44991));
    Odrv4 I__9592 (
            .O(N__44991),
            .I(n15258));
    InMux I__9591 (
            .O(N__44988),
            .I(bfn_13_17_0_));
    InMux I__9590 (
            .O(N__44985),
            .I(N__44982));
    LocalMux I__9589 (
            .O(N__44982),
            .I(N__44979));
    Odrv4 I__9588 (
            .O(N__44979),
            .I(n1700));
    InMux I__9587 (
            .O(N__44976),
            .I(n12577));
    InMux I__9586 (
            .O(N__44973),
            .I(N__44970));
    LocalMux I__9585 (
            .O(N__44970),
            .I(N__44967));
    Odrv4 I__9584 (
            .O(N__44967),
            .I(n1699));
    InMux I__9583 (
            .O(N__44964),
            .I(n12578));
    InMux I__9582 (
            .O(N__44961),
            .I(n12579));
    InMux I__9581 (
            .O(N__44958),
            .I(n12580));
    InMux I__9580 (
            .O(N__44955),
            .I(N__44951));
    InMux I__9579 (
            .O(N__44954),
            .I(N__44948));
    LocalMux I__9578 (
            .O(N__44951),
            .I(N__44943));
    LocalMux I__9577 (
            .O(N__44948),
            .I(N__44943));
    Span4Mux_s3_v I__9576 (
            .O(N__44943),
            .I(N__44940));
    Odrv4 I__9575 (
            .O(N__44940),
            .I(duty_12));
    InMux I__9574 (
            .O(N__44937),
            .I(N__44934));
    LocalMux I__9573 (
            .O(N__44934),
            .I(N__44931));
    Span4Mux_h I__9572 (
            .O(N__44931),
            .I(N__44928));
    Odrv4 I__9571 (
            .O(N__44928),
            .I(n13_adj_585));
    CascadeMux I__9570 (
            .O(N__44925),
            .I(n31_adj_674_cascade_));
    InMux I__9569 (
            .O(N__44922),
            .I(N__44919));
    LocalMux I__9568 (
            .O(N__44919),
            .I(n15230));
    InMux I__9567 (
            .O(N__44916),
            .I(N__44913));
    LocalMux I__9566 (
            .O(N__44913),
            .I(n15237));
    CascadeMux I__9565 (
            .O(N__44910),
            .I(n15195_cascade_));
    InMux I__9564 (
            .O(N__44907),
            .I(N__44904));
    LocalMux I__9563 (
            .O(N__44904),
            .I(N__44901));
    Odrv4 I__9562 (
            .O(N__44901),
            .I(n15241));
    InMux I__9561 (
            .O(N__44898),
            .I(N__44895));
    LocalMux I__9560 (
            .O(N__44895),
            .I(n15097));
    InMux I__9559 (
            .O(N__44892),
            .I(N__44889));
    LocalMux I__9558 (
            .O(N__44889),
            .I(n10_adj_659));
    InMux I__9557 (
            .O(N__44886),
            .I(N__44883));
    LocalMux I__9556 (
            .O(N__44883),
            .I(n30_adj_673));
    InMux I__9555 (
            .O(N__44880),
            .I(N__44875));
    InMux I__9554 (
            .O(N__44879),
            .I(N__44870));
    InMux I__9553 (
            .O(N__44878),
            .I(N__44870));
    LocalMux I__9552 (
            .O(N__44875),
            .I(pwm_setpoint_21));
    LocalMux I__9551 (
            .O(N__44870),
            .I(pwm_setpoint_21));
    InMux I__9550 (
            .O(N__44865),
            .I(N__44862));
    LocalMux I__9549 (
            .O(N__44862),
            .I(N__44859));
    Odrv4 I__9548 (
            .O(N__44859),
            .I(pwm_setpoint_23_N_171_12));
    InMux I__9547 (
            .O(N__44856),
            .I(N__44853));
    LocalMux I__9546 (
            .O(N__44853),
            .I(n39_adj_676));
    CascadeMux I__9545 (
            .O(N__44850),
            .I(N__44847));
    InMux I__9544 (
            .O(N__44847),
            .I(N__44844));
    LocalMux I__9543 (
            .O(N__44844),
            .I(N__44841));
    Odrv4 I__9542 (
            .O(N__44841),
            .I(n41_adj_678));
    InMux I__9541 (
            .O(N__44838),
            .I(N__44835));
    LocalMux I__9540 (
            .O(N__44835),
            .I(N__44832));
    Odrv12 I__9539 (
            .O(N__44832),
            .I(n15091));
    InMux I__9538 (
            .O(N__44829),
            .I(N__44826));
    LocalMux I__9537 (
            .O(N__44826),
            .I(N__44823));
    Odrv4 I__9536 (
            .O(N__44823),
            .I(n4_adj_655));
    InMux I__9535 (
            .O(N__44820),
            .I(N__44816));
    InMux I__9534 (
            .O(N__44819),
            .I(N__44813));
    LocalMux I__9533 (
            .O(N__44816),
            .I(pwm_setpoint_12));
    LocalMux I__9532 (
            .O(N__44813),
            .I(pwm_setpoint_12));
    InMux I__9531 (
            .O(N__44808),
            .I(N__44802));
    InMux I__9530 (
            .O(N__44807),
            .I(N__44802));
    LocalMux I__9529 (
            .O(N__44802),
            .I(n25_adj_670));
    InMux I__9528 (
            .O(N__44799),
            .I(N__44796));
    LocalMux I__9527 (
            .O(N__44796),
            .I(N__44793));
    Odrv4 I__9526 (
            .O(N__44793),
            .I(n15110));
    InMux I__9525 (
            .O(N__44790),
            .I(N__44785));
    InMux I__9524 (
            .O(N__44789),
            .I(N__44782));
    InMux I__9523 (
            .O(N__44788),
            .I(N__44779));
    LocalMux I__9522 (
            .O(N__44785),
            .I(N__44774));
    LocalMux I__9521 (
            .O(N__44782),
            .I(N__44774));
    LocalMux I__9520 (
            .O(N__44779),
            .I(n23_adj_668));
    Odrv4 I__9519 (
            .O(N__44774),
            .I(n23_adj_668));
    CascadeMux I__9518 (
            .O(N__44769),
            .I(n25_adj_670_cascade_));
    InMux I__9517 (
            .O(N__44766),
            .I(N__44760));
    InMux I__9516 (
            .O(N__44765),
            .I(N__44760));
    LocalMux I__9515 (
            .O(N__44760),
            .I(n43));
    CascadeMux I__9514 (
            .O(N__44757),
            .I(N__44754));
    InMux I__9513 (
            .O(N__44754),
            .I(N__44751));
    LocalMux I__9512 (
            .O(N__44751),
            .I(n15146));
    InMux I__9511 (
            .O(N__44748),
            .I(N__44744));
    InMux I__9510 (
            .O(N__44747),
            .I(N__44741));
    LocalMux I__9509 (
            .O(N__44744),
            .I(N__44738));
    LocalMux I__9508 (
            .O(N__44741),
            .I(n13_adj_662));
    Odrv4 I__9507 (
            .O(N__44738),
            .I(n13_adj_662));
    InMux I__9506 (
            .O(N__44733),
            .I(N__44729));
    InMux I__9505 (
            .O(N__44732),
            .I(N__44726));
    LocalMux I__9504 (
            .O(N__44729),
            .I(n15_adj_663));
    LocalMux I__9503 (
            .O(N__44726),
            .I(n15_adj_663));
    InMux I__9502 (
            .O(N__44721),
            .I(N__44718));
    LocalMux I__9501 (
            .O(N__44718),
            .I(n15229));
    InMux I__9500 (
            .O(N__44715),
            .I(N__44712));
    LocalMux I__9499 (
            .O(N__44712),
            .I(N__44708));
    InMux I__9498 (
            .O(N__44711),
            .I(N__44705));
    Odrv4 I__9497 (
            .O(N__44708),
            .I(pwm_setpoint_22));
    LocalMux I__9496 (
            .O(N__44705),
            .I(pwm_setpoint_22));
    CascadeMux I__9495 (
            .O(N__44700),
            .I(n45_cascade_));
    InMux I__9494 (
            .O(N__44697),
            .I(N__44691));
    InMux I__9493 (
            .O(N__44696),
            .I(N__44691));
    LocalMux I__9492 (
            .O(N__44691),
            .I(pwm_setpoint_20));
    CascadeMux I__9491 (
            .O(N__44688),
            .I(n41_adj_678_cascade_));
    InMux I__9490 (
            .O(N__44685),
            .I(N__44682));
    LocalMux I__9489 (
            .O(N__44682),
            .I(n40_adj_677));
    InMux I__9488 (
            .O(N__44679),
            .I(N__44674));
    InMux I__9487 (
            .O(N__44678),
            .I(N__44669));
    InMux I__9486 (
            .O(N__44677),
            .I(N__44669));
    LocalMux I__9485 (
            .O(N__44674),
            .I(n45));
    LocalMux I__9484 (
            .O(N__44669),
            .I(n45));
    InMux I__9483 (
            .O(N__44664),
            .I(N__44661));
    LocalMux I__9482 (
            .O(N__44661),
            .I(n15223));
    InMux I__9481 (
            .O(N__44658),
            .I(N__44655));
    LocalMux I__9480 (
            .O(N__44655),
            .I(N__44652));
    Odrv4 I__9479 (
            .O(N__44652),
            .I(n15165));
    InMux I__9478 (
            .O(N__44649),
            .I(N__44646));
    LocalMux I__9477 (
            .O(N__44646),
            .I(n15243));
    InMux I__9476 (
            .O(N__44643),
            .I(N__44640));
    LocalMux I__9475 (
            .O(N__44640),
            .I(N__44636));
    InMux I__9474 (
            .O(N__44639),
            .I(N__44633));
    Span4Mux_h I__9473 (
            .O(N__44636),
            .I(N__44628));
    LocalMux I__9472 (
            .O(N__44633),
            .I(N__44628));
    Odrv4 I__9471 (
            .O(N__44628),
            .I(duty_22));
    InMux I__9470 (
            .O(N__44625),
            .I(N__44622));
    LocalMux I__9469 (
            .O(N__44622),
            .I(n3_adj_575));
    InMux I__9468 (
            .O(N__44619),
            .I(N__44613));
    InMux I__9467 (
            .O(N__44618),
            .I(N__44613));
    LocalMux I__9466 (
            .O(N__44613),
            .I(N__44610));
    Odrv4 I__9465 (
            .O(N__44610),
            .I(pwm_setpoint_19));
    CascadeMux I__9464 (
            .O(N__44607),
            .I(n39_adj_676_cascade_));
    InMux I__9463 (
            .O(N__44604),
            .I(N__44601));
    LocalMux I__9462 (
            .O(N__44601),
            .I(n15254));
    InMux I__9461 (
            .O(N__44598),
            .I(N__44595));
    LocalMux I__9460 (
            .O(N__44595),
            .I(N__44592));
    Span4Mux_s3_v I__9459 (
            .O(N__44592),
            .I(N__44588));
    InMux I__9458 (
            .O(N__44591),
            .I(N__44585));
    Odrv4 I__9457 (
            .O(N__44588),
            .I(duty_17));
    LocalMux I__9456 (
            .O(N__44585),
            .I(duty_17));
    InMux I__9455 (
            .O(N__44580),
            .I(N__44577));
    LocalMux I__9454 (
            .O(N__44577),
            .I(n8_adj_580));
    InMux I__9453 (
            .O(N__44574),
            .I(N__44571));
    LocalMux I__9452 (
            .O(N__44571),
            .I(N__44567));
    InMux I__9451 (
            .O(N__44570),
            .I(N__44564));
    Odrv4 I__9450 (
            .O(N__44567),
            .I(duty_21));
    LocalMux I__9449 (
            .O(N__44564),
            .I(duty_21));
    InMux I__9448 (
            .O(N__44559),
            .I(N__44556));
    LocalMux I__9447 (
            .O(N__44556),
            .I(n4_adj_576));
    InMux I__9446 (
            .O(N__44553),
            .I(N__44550));
    LocalMux I__9445 (
            .O(N__44550),
            .I(N__44547));
    Span4Mux_s2_v I__9444 (
            .O(N__44547),
            .I(N__44544));
    Span4Mux_h I__9443 (
            .O(N__44544),
            .I(N__44540));
    InMux I__9442 (
            .O(N__44543),
            .I(N__44537));
    Odrv4 I__9441 (
            .O(N__44540),
            .I(duty_18));
    LocalMux I__9440 (
            .O(N__44537),
            .I(duty_18));
    InMux I__9439 (
            .O(N__44532),
            .I(N__44529));
    LocalMux I__9438 (
            .O(N__44529),
            .I(n7_adj_579));
    InMux I__9437 (
            .O(N__44526),
            .I(N__44523));
    LocalMux I__9436 (
            .O(N__44523),
            .I(pwm_setpoint_23_N_171_19));
    InMux I__9435 (
            .O(N__44520),
            .I(N__44517));
    LocalMux I__9434 (
            .O(N__44517),
            .I(pwm_setpoint_23_N_171_20));
    InMux I__9433 (
            .O(N__44514),
            .I(N__44511));
    LocalMux I__9432 (
            .O(N__44511),
            .I(N__44508));
    Odrv4 I__9431 (
            .O(N__44508),
            .I(pwm_setpoint_23_N_171_0));
    InMux I__9430 (
            .O(N__44505),
            .I(N__44502));
    LocalMux I__9429 (
            .O(N__44502),
            .I(N__44498));
    InMux I__9428 (
            .O(N__44501),
            .I(N__44495));
    Odrv12 I__9427 (
            .O(N__44498),
            .I(duty_0));
    LocalMux I__9426 (
            .O(N__44495),
            .I(duty_0));
    InMux I__9425 (
            .O(N__44490),
            .I(N__44487));
    LocalMux I__9424 (
            .O(N__44487),
            .I(pwm_setpoint_0));
    InMux I__9423 (
            .O(N__44484),
            .I(N__44478));
    InMux I__9422 (
            .O(N__44483),
            .I(N__44478));
    LocalMux I__9421 (
            .O(N__44478),
            .I(duty_20));
    InMux I__9420 (
            .O(N__44475),
            .I(N__44472));
    LocalMux I__9419 (
            .O(N__44472),
            .I(n5_adj_577));
    InMux I__9418 (
            .O(N__44469),
            .I(N__44466));
    LocalMux I__9417 (
            .O(N__44466),
            .I(N__44463));
    Span4Mux_h I__9416 (
            .O(N__44463),
            .I(N__44460));
    Odrv4 I__9415 (
            .O(N__44460),
            .I(n10_adj_566));
    InMux I__9414 (
            .O(N__44457),
            .I(n12487));
    InMux I__9413 (
            .O(N__44454),
            .I(N__44451));
    LocalMux I__9412 (
            .O(N__44451),
            .I(N__44447));
    InMux I__9411 (
            .O(N__44450),
            .I(N__44444));
    Span4Mux_v I__9410 (
            .O(N__44447),
            .I(N__44439));
    LocalMux I__9409 (
            .O(N__44444),
            .I(N__44439));
    Span4Mux_h I__9408 (
            .O(N__44439),
            .I(N__44436));
    Odrv4 I__9407 (
            .O(N__44436),
            .I(duty_16));
    InMux I__9406 (
            .O(N__44433),
            .I(bfn_12_27_0_));
    InMux I__9405 (
            .O(N__44430),
            .I(N__44427));
    LocalMux I__9404 (
            .O(N__44427),
            .I(N__44424));
    Span4Mux_v I__9403 (
            .O(N__44424),
            .I(N__44421));
    Odrv4 I__9402 (
            .O(N__44421),
            .I(n8_adj_568));
    InMux I__9401 (
            .O(N__44418),
            .I(n12489));
    InMux I__9400 (
            .O(N__44415),
            .I(N__44412));
    LocalMux I__9399 (
            .O(N__44412),
            .I(N__44409));
    Odrv4 I__9398 (
            .O(N__44409),
            .I(n7_adj_569));
    InMux I__9397 (
            .O(N__44406),
            .I(n12490));
    InMux I__9396 (
            .O(N__44403),
            .I(N__44400));
    LocalMux I__9395 (
            .O(N__44400),
            .I(N__44397));
    Odrv4 I__9394 (
            .O(N__44397),
            .I(n6_adj_570));
    InMux I__9393 (
            .O(N__44394),
            .I(n12491));
    InMux I__9392 (
            .O(N__44391),
            .I(N__44388));
    LocalMux I__9391 (
            .O(N__44388),
            .I(N__44385));
    Span4Mux_v I__9390 (
            .O(N__44385),
            .I(N__44382));
    Odrv4 I__9389 (
            .O(N__44382),
            .I(n5_adj_571));
    InMux I__9388 (
            .O(N__44379),
            .I(n12492));
    InMux I__9387 (
            .O(N__44376),
            .I(N__44373));
    LocalMux I__9386 (
            .O(N__44373),
            .I(N__44370));
    Odrv4 I__9385 (
            .O(N__44370),
            .I(n4_adj_572));
    InMux I__9384 (
            .O(N__44367),
            .I(n12493));
    InMux I__9383 (
            .O(N__44364),
            .I(N__44361));
    LocalMux I__9382 (
            .O(N__44361),
            .I(N__44358));
    Odrv4 I__9381 (
            .O(N__44358),
            .I(n3_adj_573));
    InMux I__9380 (
            .O(N__44355),
            .I(n12494));
    InMux I__9379 (
            .O(N__44352),
            .I(N__44349));
    LocalMux I__9378 (
            .O(N__44349),
            .I(N__44346));
    Odrv4 I__9377 (
            .O(N__44346),
            .I(n2_adj_574));
    InMux I__9376 (
            .O(N__44343),
            .I(n12495));
    InMux I__9375 (
            .O(N__44340),
            .I(N__44337));
    LocalMux I__9374 (
            .O(N__44337),
            .I(N__44334));
    Span4Mux_h I__9373 (
            .O(N__44334),
            .I(N__44330));
    InMux I__9372 (
            .O(N__44333),
            .I(N__44327));
    Odrv4 I__9371 (
            .O(N__44330),
            .I(duty_7));
    LocalMux I__9370 (
            .O(N__44327),
            .I(duty_7));
    InMux I__9369 (
            .O(N__44322),
            .I(n12479));
    InMux I__9368 (
            .O(N__44319),
            .I(N__44316));
    LocalMux I__9367 (
            .O(N__44316),
            .I(N__44313));
    Odrv4 I__9366 (
            .O(N__44313),
            .I(n17_adj_559));
    InMux I__9365 (
            .O(N__44310),
            .I(N__44306));
    InMux I__9364 (
            .O(N__44309),
            .I(N__44303));
    LocalMux I__9363 (
            .O(N__44306),
            .I(N__44300));
    LocalMux I__9362 (
            .O(N__44303),
            .I(N__44297));
    Span4Mux_h I__9361 (
            .O(N__44300),
            .I(N__44294));
    Span4Mux_h I__9360 (
            .O(N__44297),
            .I(N__44291));
    Span4Mux_h I__9359 (
            .O(N__44294),
            .I(N__44288));
    Odrv4 I__9358 (
            .O(N__44291),
            .I(duty_8));
    Odrv4 I__9357 (
            .O(N__44288),
            .I(duty_8));
    InMux I__9356 (
            .O(N__44283),
            .I(bfn_12_26_0_));
    InMux I__9355 (
            .O(N__44280),
            .I(N__44277));
    LocalMux I__9354 (
            .O(N__44277),
            .I(N__44274));
    Odrv4 I__9353 (
            .O(N__44274),
            .I(n16_adj_560));
    InMux I__9352 (
            .O(N__44271),
            .I(N__44267));
    InMux I__9351 (
            .O(N__44270),
            .I(N__44264));
    LocalMux I__9350 (
            .O(N__44267),
            .I(N__44261));
    LocalMux I__9349 (
            .O(N__44264),
            .I(N__44258));
    Span4Mux_v I__9348 (
            .O(N__44261),
            .I(N__44255));
    Span12Mux_s6_v I__9347 (
            .O(N__44258),
            .I(N__44252));
    Odrv4 I__9346 (
            .O(N__44255),
            .I(duty_9));
    Odrv12 I__9345 (
            .O(N__44252),
            .I(duty_9));
    InMux I__9344 (
            .O(N__44247),
            .I(n12481));
    InMux I__9343 (
            .O(N__44244),
            .I(N__44241));
    LocalMux I__9342 (
            .O(N__44241),
            .I(N__44238));
    Odrv4 I__9341 (
            .O(N__44238),
            .I(n15_adj_561));
    InMux I__9340 (
            .O(N__44235),
            .I(N__44232));
    LocalMux I__9339 (
            .O(N__44232),
            .I(N__44228));
    InMux I__9338 (
            .O(N__44231),
            .I(N__44225));
    Span4Mux_s3_v I__9337 (
            .O(N__44228),
            .I(N__44222));
    LocalMux I__9336 (
            .O(N__44225),
            .I(N__44219));
    Odrv4 I__9335 (
            .O(N__44222),
            .I(duty_10));
    Odrv4 I__9334 (
            .O(N__44219),
            .I(duty_10));
    InMux I__9333 (
            .O(N__44214),
            .I(n12482));
    InMux I__9332 (
            .O(N__44211),
            .I(N__44208));
    LocalMux I__9331 (
            .O(N__44208),
            .I(N__44205));
    Odrv4 I__9330 (
            .O(N__44205),
            .I(n14_adj_562));
    InMux I__9329 (
            .O(N__44202),
            .I(N__44198));
    InMux I__9328 (
            .O(N__44201),
            .I(N__44195));
    LocalMux I__9327 (
            .O(N__44198),
            .I(N__44192));
    LocalMux I__9326 (
            .O(N__44195),
            .I(N__44189));
    Span4Mux_v I__9325 (
            .O(N__44192),
            .I(N__44186));
    Span4Mux_v I__9324 (
            .O(N__44189),
            .I(N__44181));
    Span4Mux_h I__9323 (
            .O(N__44186),
            .I(N__44181));
    Odrv4 I__9322 (
            .O(N__44181),
            .I(duty_11));
    InMux I__9321 (
            .O(N__44178),
            .I(n12483));
    CascadeMux I__9320 (
            .O(N__44175),
            .I(N__44172));
    InMux I__9319 (
            .O(N__44172),
            .I(N__44169));
    LocalMux I__9318 (
            .O(N__44169),
            .I(N__44166));
    Odrv4 I__9317 (
            .O(N__44166),
            .I(n13_adj_563));
    InMux I__9316 (
            .O(N__44163),
            .I(n12484));
    InMux I__9315 (
            .O(N__44160),
            .I(N__44157));
    LocalMux I__9314 (
            .O(N__44157),
            .I(N__44154));
    Odrv12 I__9313 (
            .O(N__44154),
            .I(n12_adj_564));
    InMux I__9312 (
            .O(N__44151),
            .I(N__44147));
    InMux I__9311 (
            .O(N__44150),
            .I(N__44144));
    LocalMux I__9310 (
            .O(N__44147),
            .I(N__44139));
    LocalMux I__9309 (
            .O(N__44144),
            .I(N__44139));
    Span4Mux_v I__9308 (
            .O(N__44139),
            .I(N__44136));
    Odrv4 I__9307 (
            .O(N__44136),
            .I(duty_13));
    InMux I__9306 (
            .O(N__44133),
            .I(n12485));
    InMux I__9305 (
            .O(N__44130),
            .I(N__44127));
    LocalMux I__9304 (
            .O(N__44127),
            .I(N__44124));
    Odrv12 I__9303 (
            .O(N__44124),
            .I(n11_adj_565));
    InMux I__9302 (
            .O(N__44121),
            .I(N__44117));
    InMux I__9301 (
            .O(N__44120),
            .I(N__44114));
    LocalMux I__9300 (
            .O(N__44117),
            .I(N__44111));
    LocalMux I__9299 (
            .O(N__44114),
            .I(N__44108));
    Span4Mux_h I__9298 (
            .O(N__44111),
            .I(N__44105));
    Span4Mux_v I__9297 (
            .O(N__44108),
            .I(N__44100));
    Span4Mux_h I__9296 (
            .O(N__44105),
            .I(N__44100));
    Odrv4 I__9295 (
            .O(N__44100),
            .I(duty_14));
    InMux I__9294 (
            .O(N__44097),
            .I(n12486));
    InMux I__9293 (
            .O(N__44094),
            .I(N__44086));
    InMux I__9292 (
            .O(N__44093),
            .I(N__44083));
    InMux I__9291 (
            .O(N__44092),
            .I(N__44076));
    InMux I__9290 (
            .O(N__44091),
            .I(N__44076));
    InMux I__9289 (
            .O(N__44090),
            .I(N__44076));
    InMux I__9288 (
            .O(N__44089),
            .I(N__44073));
    LocalMux I__9287 (
            .O(N__44086),
            .I(n861));
    LocalMux I__9286 (
            .O(N__44083),
            .I(n861));
    LocalMux I__9285 (
            .O(N__44076),
            .I(n861));
    LocalMux I__9284 (
            .O(N__44073),
            .I(n861));
    CascadeMux I__9283 (
            .O(N__44064),
            .I(N__44060));
    CascadeMux I__9282 (
            .O(N__44063),
            .I(N__44057));
    InMux I__9281 (
            .O(N__44060),
            .I(N__44054));
    InMux I__9280 (
            .O(N__44057),
            .I(N__44051));
    LocalMux I__9279 (
            .O(N__44054),
            .I(n829));
    LocalMux I__9278 (
            .O(N__44051),
            .I(n829));
    InMux I__9277 (
            .O(N__44046),
            .I(N__44043));
    LocalMux I__9276 (
            .O(N__44043),
            .I(n896));
    InMux I__9275 (
            .O(N__44040),
            .I(bfn_12_25_0_));
    InMux I__9274 (
            .O(N__44037),
            .I(N__44034));
    LocalMux I__9273 (
            .O(N__44034),
            .I(N__44031));
    Odrv4 I__9272 (
            .O(N__44031),
            .I(n24_adj_552));
    InMux I__9271 (
            .O(N__44028),
            .I(n12473));
    InMux I__9270 (
            .O(N__44025),
            .I(N__44022));
    LocalMux I__9269 (
            .O(N__44022),
            .I(n23_adj_553));
    InMux I__9268 (
            .O(N__44019),
            .I(n12474));
    InMux I__9267 (
            .O(N__44016),
            .I(N__44013));
    LocalMux I__9266 (
            .O(N__44013),
            .I(n22_adj_554));
    InMux I__9265 (
            .O(N__44010),
            .I(n12475));
    InMux I__9264 (
            .O(N__44007),
            .I(N__44004));
    LocalMux I__9263 (
            .O(N__44004),
            .I(N__44001));
    Odrv4 I__9262 (
            .O(N__44001),
            .I(n21_adj_555));
    InMux I__9261 (
            .O(N__43998),
            .I(N__43995));
    LocalMux I__9260 (
            .O(N__43995),
            .I(N__43992));
    Span4Mux_v I__9259 (
            .O(N__43992),
            .I(N__43988));
    InMux I__9258 (
            .O(N__43991),
            .I(N__43985));
    Odrv4 I__9257 (
            .O(N__43988),
            .I(duty_4));
    LocalMux I__9256 (
            .O(N__43985),
            .I(duty_4));
    InMux I__9255 (
            .O(N__43980),
            .I(n12476));
    InMux I__9254 (
            .O(N__43977),
            .I(N__43974));
    LocalMux I__9253 (
            .O(N__43974),
            .I(N__43971));
    Odrv4 I__9252 (
            .O(N__43971),
            .I(n20_adj_556));
    InMux I__9251 (
            .O(N__43968),
            .I(N__43965));
    LocalMux I__9250 (
            .O(N__43965),
            .I(N__43962));
    Span4Mux_v I__9249 (
            .O(N__43962),
            .I(N__43959));
    Sp12to4 I__9248 (
            .O(N__43959),
            .I(N__43955));
    InMux I__9247 (
            .O(N__43958),
            .I(N__43952));
    Odrv12 I__9246 (
            .O(N__43955),
            .I(duty_5));
    LocalMux I__9245 (
            .O(N__43952),
            .I(duty_5));
    InMux I__9244 (
            .O(N__43947),
            .I(n12477));
    InMux I__9243 (
            .O(N__43944),
            .I(N__43941));
    LocalMux I__9242 (
            .O(N__43941),
            .I(n19_adj_557));
    InMux I__9241 (
            .O(N__43938),
            .I(n12478));
    InMux I__9240 (
            .O(N__43935),
            .I(N__43932));
    LocalMux I__9239 (
            .O(N__43932),
            .I(N__43929));
    Span4Mux_h I__9238 (
            .O(N__43929),
            .I(N__43926));
    Span4Mux_h I__9237 (
            .O(N__43926),
            .I(N__43923));
    Odrv4 I__9236 (
            .O(N__43923),
            .I(n18_adj_558));
    CascadeMux I__9235 (
            .O(N__43920),
            .I(N__43917));
    InMux I__9234 (
            .O(N__43917),
            .I(N__43913));
    InMux I__9233 (
            .O(N__43916),
            .I(N__43910));
    LocalMux I__9232 (
            .O(N__43913),
            .I(N__43906));
    LocalMux I__9231 (
            .O(N__43910),
            .I(N__43903));
    InMux I__9230 (
            .O(N__43909),
            .I(N__43900));
    Span4Mux_h I__9229 (
            .O(N__43906),
            .I(N__43897));
    Span4Mux_v I__9228 (
            .O(N__43903),
            .I(N__43894));
    LocalMux I__9227 (
            .O(N__43900),
            .I(encoder0_position_25));
    Odrv4 I__9226 (
            .O(N__43897),
            .I(encoder0_position_25));
    Odrv4 I__9225 (
            .O(N__43894),
            .I(encoder0_position_25));
    InMux I__9224 (
            .O(N__43887),
            .I(N__43884));
    LocalMux I__9223 (
            .O(N__43884),
            .I(N__43881));
    Span4Mux_h I__9222 (
            .O(N__43881),
            .I(N__43878));
    Odrv4 I__9221 (
            .O(N__43878),
            .I(n8));
    InMux I__9220 (
            .O(N__43875),
            .I(N__43871));
    InMux I__9219 (
            .O(N__43874),
            .I(N__43868));
    LocalMux I__9218 (
            .O(N__43871),
            .I(n41));
    LocalMux I__9217 (
            .O(N__43868),
            .I(n41));
    InMux I__9216 (
            .O(N__43863),
            .I(N__43860));
    LocalMux I__9215 (
            .O(N__43860),
            .I(n901));
    CascadeMux I__9214 (
            .O(N__43857),
            .I(n41_cascade_));
    CascadeMux I__9213 (
            .O(N__43854),
            .I(n933_cascade_));
    CascadeMux I__9212 (
            .O(N__43851),
            .I(N__43848));
    InMux I__9211 (
            .O(N__43848),
            .I(N__43845));
    LocalMux I__9210 (
            .O(N__43845),
            .I(N__43842));
    Odrv12 I__9209 (
            .O(N__43842),
            .I(n10));
    InMux I__9208 (
            .O(N__43839),
            .I(N__43834));
    InMux I__9207 (
            .O(N__43838),
            .I(N__43831));
    InMux I__9206 (
            .O(N__43837),
            .I(N__43828));
    LocalMux I__9205 (
            .O(N__43834),
            .I(N__43825));
    LocalMux I__9204 (
            .O(N__43831),
            .I(N__43822));
    LocalMux I__9203 (
            .O(N__43828),
            .I(N__43817));
    Span4Mux_v I__9202 (
            .O(N__43825),
            .I(N__43817));
    Span4Mux_h I__9201 (
            .O(N__43822),
            .I(N__43814));
    Odrv4 I__9200 (
            .O(N__43817),
            .I(encoder0_position_23));
    Odrv4 I__9199 (
            .O(N__43814),
            .I(encoder0_position_23));
    CascadeMux I__9198 (
            .O(N__43809),
            .I(N__43805));
    InMux I__9197 (
            .O(N__43808),
            .I(N__43802));
    InMux I__9196 (
            .O(N__43805),
            .I(N__43798));
    LocalMux I__9195 (
            .O(N__43802),
            .I(N__43795));
    InMux I__9194 (
            .O(N__43801),
            .I(N__43792));
    LocalMux I__9193 (
            .O(N__43798),
            .I(N__43787));
    Span4Mux_v I__9192 (
            .O(N__43795),
            .I(N__43787));
    LocalMux I__9191 (
            .O(N__43792),
            .I(N__43784));
    Odrv4 I__9190 (
            .O(N__43787),
            .I(encoder0_position_24));
    Odrv12 I__9189 (
            .O(N__43784),
            .I(encoder0_position_24));
    InMux I__9188 (
            .O(N__43779),
            .I(N__43776));
    LocalMux I__9187 (
            .O(N__43776),
            .I(N__43773));
    Span4Mux_v I__9186 (
            .O(N__43773),
            .I(N__43770));
    Span4Mux_h I__9185 (
            .O(N__43770),
            .I(N__43767));
    Odrv4 I__9184 (
            .O(N__43767),
            .I(n9));
    CascadeMux I__9183 (
            .O(N__43764),
            .I(n295_cascade_));
    CascadeMux I__9182 (
            .O(N__43761),
            .I(n11955_cascade_));
    InMux I__9181 (
            .O(N__43758),
            .I(N__43755));
    LocalMux I__9180 (
            .O(N__43755),
            .I(n14460));
    CascadeMux I__9179 (
            .O(N__43752),
            .I(n960_cascade_));
    CascadeMux I__9178 (
            .O(N__43749),
            .I(N__43745));
    InMux I__9177 (
            .O(N__43748),
            .I(N__43742));
    InMux I__9176 (
            .O(N__43745),
            .I(N__43739));
    LocalMux I__9175 (
            .O(N__43742),
            .I(N__43736));
    LocalMux I__9174 (
            .O(N__43739),
            .I(N__43730));
    Span4Mux_h I__9173 (
            .O(N__43736),
            .I(N__43730));
    InMux I__9172 (
            .O(N__43735),
            .I(N__43727));
    Span4Mux_v I__9171 (
            .O(N__43730),
            .I(N__43724));
    LocalMux I__9170 (
            .O(N__43727),
            .I(n1818));
    Odrv4 I__9169 (
            .O(N__43724),
            .I(n1818));
    CascadeMux I__9168 (
            .O(N__43719),
            .I(N__43716));
    InMux I__9167 (
            .O(N__43716),
            .I(N__43713));
    LocalMux I__9166 (
            .O(N__43713),
            .I(N__43710));
    Span4Mux_v I__9165 (
            .O(N__43710),
            .I(N__43707));
    Odrv4 I__9164 (
            .O(N__43707),
            .I(n10_adj_628));
    InMux I__9163 (
            .O(N__43704),
            .I(N__43701));
    LocalMux I__9162 (
            .O(N__43701),
            .I(N__43698));
    Span4Mux_h I__9161 (
            .O(N__43698),
            .I(N__43695));
    Odrv4 I__9160 (
            .O(N__43695),
            .I(n17));
    InMux I__9159 (
            .O(N__43692),
            .I(N__43689));
    LocalMux I__9158 (
            .O(N__43689),
            .I(N__43684));
    InMux I__9157 (
            .O(N__43688),
            .I(N__43681));
    InMux I__9156 (
            .O(N__43687),
            .I(N__43678));
    Span4Mux_v I__9155 (
            .O(N__43684),
            .I(N__43671));
    LocalMux I__9154 (
            .O(N__43681),
            .I(N__43671));
    LocalMux I__9153 (
            .O(N__43678),
            .I(N__43671));
    Odrv4 I__9152 (
            .O(N__43671),
            .I(n303));
    InMux I__9151 (
            .O(N__43668),
            .I(N__43665));
    LocalMux I__9150 (
            .O(N__43665),
            .I(N__43662));
    Span4Mux_v I__9149 (
            .O(N__43662),
            .I(N__43659));
    Odrv4 I__9148 (
            .O(N__43659),
            .I(n15));
    CascadeMux I__9147 (
            .O(N__43656),
            .I(N__43652));
    InMux I__9146 (
            .O(N__43655),
            .I(N__43649));
    InMux I__9145 (
            .O(N__43652),
            .I(N__43645));
    LocalMux I__9144 (
            .O(N__43649),
            .I(N__43642));
    InMux I__9143 (
            .O(N__43648),
            .I(N__43639));
    LocalMux I__9142 (
            .O(N__43645),
            .I(N__43634));
    Span4Mux_v I__9141 (
            .O(N__43642),
            .I(N__43634));
    LocalMux I__9140 (
            .O(N__43639),
            .I(N__43631));
    Odrv4 I__9139 (
            .O(N__43634),
            .I(encoder0_position_18));
    Odrv12 I__9138 (
            .O(N__43631),
            .I(encoder0_position_18));
    InMux I__9137 (
            .O(N__43626),
            .I(N__43623));
    LocalMux I__9136 (
            .O(N__43623),
            .I(n899));
    CascadeMux I__9135 (
            .O(N__43620),
            .I(N__43616));
    CascadeMux I__9134 (
            .O(N__43619),
            .I(N__43613));
    InMux I__9133 (
            .O(N__43616),
            .I(N__43610));
    InMux I__9132 (
            .O(N__43613),
            .I(N__43607));
    LocalMux I__9131 (
            .O(N__43610),
            .I(N__43604));
    LocalMux I__9130 (
            .O(N__43607),
            .I(n832));
    Odrv4 I__9129 (
            .O(N__43604),
            .I(n832));
    InMux I__9128 (
            .O(N__43599),
            .I(N__43596));
    LocalMux I__9127 (
            .O(N__43596),
            .I(n900));
    CascadeMux I__9126 (
            .O(N__43593),
            .I(N__43589));
    CascadeMux I__9125 (
            .O(N__43592),
            .I(N__43586));
    InMux I__9124 (
            .O(N__43589),
            .I(N__43582));
    InMux I__9123 (
            .O(N__43586),
            .I(N__43579));
    InMux I__9122 (
            .O(N__43585),
            .I(N__43576));
    LocalMux I__9121 (
            .O(N__43582),
            .I(N__43571));
    LocalMux I__9120 (
            .O(N__43579),
            .I(N__43571));
    LocalMux I__9119 (
            .O(N__43576),
            .I(n833));
    Odrv4 I__9118 (
            .O(N__43571),
            .I(n833));
    CascadeMux I__9117 (
            .O(N__43566),
            .I(n932_cascade_));
    InMux I__9116 (
            .O(N__43563),
            .I(n12597));
    CascadeMux I__9115 (
            .O(N__43560),
            .I(N__43557));
    InMux I__9114 (
            .O(N__43557),
            .I(N__43554));
    LocalMux I__9113 (
            .O(N__43554),
            .I(N__43550));
    InMux I__9112 (
            .O(N__43553),
            .I(N__43547));
    Span4Mux_v I__9111 (
            .O(N__43550),
            .I(N__43544));
    LocalMux I__9110 (
            .O(N__43547),
            .I(n1726));
    Odrv4 I__9109 (
            .O(N__43544),
            .I(n1726));
    CascadeMux I__9108 (
            .O(N__43539),
            .I(N__43536));
    InMux I__9107 (
            .O(N__43536),
            .I(N__43533));
    LocalMux I__9106 (
            .O(N__43533),
            .I(N__43530));
    Span4Mux_h I__9105 (
            .O(N__43530),
            .I(N__43527));
    Odrv4 I__9104 (
            .O(N__43527),
            .I(n1793));
    InMux I__9103 (
            .O(N__43524),
            .I(bfn_12_21_0_));
    InMux I__9102 (
            .O(N__43521),
            .I(N__43518));
    LocalMux I__9101 (
            .O(N__43518),
            .I(N__43515));
    Span4Mux_h I__9100 (
            .O(N__43515),
            .I(N__43512));
    Odrv4 I__9099 (
            .O(N__43512),
            .I(n1792));
    InMux I__9098 (
            .O(N__43509),
            .I(n12599));
    InMux I__9097 (
            .O(N__43506),
            .I(N__43503));
    LocalMux I__9096 (
            .O(N__43503),
            .I(N__43500));
    Span4Mux_h I__9095 (
            .O(N__43500),
            .I(N__43497));
    Odrv4 I__9094 (
            .O(N__43497),
            .I(n1791));
    InMux I__9093 (
            .O(N__43494),
            .I(n12600));
    CascadeMux I__9092 (
            .O(N__43491),
            .I(N__43488));
    InMux I__9091 (
            .O(N__43488),
            .I(N__43484));
    InMux I__9090 (
            .O(N__43487),
            .I(N__43480));
    LocalMux I__9089 (
            .O(N__43484),
            .I(N__43477));
    InMux I__9088 (
            .O(N__43483),
            .I(N__43474));
    LocalMux I__9087 (
            .O(N__43480),
            .I(n1723));
    Odrv4 I__9086 (
            .O(N__43477),
            .I(n1723));
    LocalMux I__9085 (
            .O(N__43474),
            .I(n1723));
    InMux I__9084 (
            .O(N__43467),
            .I(N__43464));
    LocalMux I__9083 (
            .O(N__43464),
            .I(N__43461));
    Odrv4 I__9082 (
            .O(N__43461),
            .I(n1790));
    InMux I__9081 (
            .O(N__43458),
            .I(n12601));
    CascadeMux I__9080 (
            .O(N__43455),
            .I(N__43452));
    InMux I__9079 (
            .O(N__43452),
            .I(N__43449));
    LocalMux I__9078 (
            .O(N__43449),
            .I(N__43445));
    InMux I__9077 (
            .O(N__43448),
            .I(N__43442));
    Odrv4 I__9076 (
            .O(N__43445),
            .I(n1722));
    LocalMux I__9075 (
            .O(N__43442),
            .I(n1722));
    InMux I__9074 (
            .O(N__43437),
            .I(N__43434));
    LocalMux I__9073 (
            .O(N__43434),
            .I(N__43431));
    Odrv4 I__9072 (
            .O(N__43431),
            .I(n1789));
    InMux I__9071 (
            .O(N__43428),
            .I(n12602));
    CascadeMux I__9070 (
            .O(N__43425),
            .I(N__43422));
    InMux I__9069 (
            .O(N__43422),
            .I(N__43419));
    LocalMux I__9068 (
            .O(N__43419),
            .I(N__43415));
    InMux I__9067 (
            .O(N__43418),
            .I(N__43412));
    Odrv4 I__9066 (
            .O(N__43415),
            .I(n1721));
    LocalMux I__9065 (
            .O(N__43412),
            .I(n1721));
    InMux I__9064 (
            .O(N__43407),
            .I(N__43404));
    LocalMux I__9063 (
            .O(N__43404),
            .I(N__43401));
    Odrv12 I__9062 (
            .O(N__43401),
            .I(n1788));
    InMux I__9061 (
            .O(N__43398),
            .I(n12603));
    CascadeMux I__9060 (
            .O(N__43395),
            .I(N__43392));
    InMux I__9059 (
            .O(N__43392),
            .I(N__43387));
    InMux I__9058 (
            .O(N__43391),
            .I(N__43384));
    InMux I__9057 (
            .O(N__43390),
            .I(N__43381));
    LocalMux I__9056 (
            .O(N__43387),
            .I(N__43376));
    LocalMux I__9055 (
            .O(N__43384),
            .I(N__43376));
    LocalMux I__9054 (
            .O(N__43381),
            .I(N__43373));
    Odrv4 I__9053 (
            .O(N__43376),
            .I(n1720));
    Odrv4 I__9052 (
            .O(N__43373),
            .I(n1720));
    InMux I__9051 (
            .O(N__43368),
            .I(N__43365));
    LocalMux I__9050 (
            .O(N__43365),
            .I(n1787));
    InMux I__9049 (
            .O(N__43362),
            .I(n12604));
    InMux I__9048 (
            .O(N__43359),
            .I(n12605));
    CascadeMux I__9047 (
            .O(N__43356),
            .I(n1731_cascade_));
    InMux I__9046 (
            .O(N__43353),
            .I(N__43350));
    LocalMux I__9045 (
            .O(N__43350),
            .I(n11991));
    InMux I__9044 (
            .O(N__43347),
            .I(N__43344));
    LocalMux I__9043 (
            .O(N__43344),
            .I(N__43341));
    Span4Mux_h I__9042 (
            .O(N__43341),
            .I(N__43338));
    Odrv4 I__9041 (
            .O(N__43338),
            .I(n1801));
    InMux I__9040 (
            .O(N__43335),
            .I(bfn_12_20_0_));
    InMux I__9039 (
            .O(N__43332),
            .I(N__43329));
    LocalMux I__9038 (
            .O(N__43329),
            .I(N__43326));
    Span4Mux_h I__9037 (
            .O(N__43326),
            .I(N__43323));
    Odrv4 I__9036 (
            .O(N__43323),
            .I(n1800));
    InMux I__9035 (
            .O(N__43320),
            .I(n12591));
    CascadeMux I__9034 (
            .O(N__43317),
            .I(N__43314));
    InMux I__9033 (
            .O(N__43314),
            .I(N__43311));
    LocalMux I__9032 (
            .O(N__43311),
            .I(N__43307));
    CascadeMux I__9031 (
            .O(N__43310),
            .I(N__43304));
    Span4Mux_v I__9030 (
            .O(N__43307),
            .I(N__43300));
    InMux I__9029 (
            .O(N__43304),
            .I(N__43297));
    InMux I__9028 (
            .O(N__43303),
            .I(N__43294));
    Odrv4 I__9027 (
            .O(N__43300),
            .I(n1732));
    LocalMux I__9026 (
            .O(N__43297),
            .I(n1732));
    LocalMux I__9025 (
            .O(N__43294),
            .I(n1732));
    InMux I__9024 (
            .O(N__43287),
            .I(N__43284));
    LocalMux I__9023 (
            .O(N__43284),
            .I(N__43281));
    Span4Mux_h I__9022 (
            .O(N__43281),
            .I(N__43278));
    Odrv4 I__9021 (
            .O(N__43278),
            .I(n1799));
    InMux I__9020 (
            .O(N__43275),
            .I(n12592));
    InMux I__9019 (
            .O(N__43272),
            .I(N__43268));
    CascadeMux I__9018 (
            .O(N__43271),
            .I(N__43265));
    LocalMux I__9017 (
            .O(N__43268),
            .I(N__43262));
    InMux I__9016 (
            .O(N__43265),
            .I(N__43259));
    Odrv4 I__9015 (
            .O(N__43262),
            .I(n1731));
    LocalMux I__9014 (
            .O(N__43259),
            .I(n1731));
    InMux I__9013 (
            .O(N__43254),
            .I(N__43251));
    LocalMux I__9012 (
            .O(N__43251),
            .I(N__43248));
    Odrv4 I__9011 (
            .O(N__43248),
            .I(n1798));
    InMux I__9010 (
            .O(N__43245),
            .I(n12593));
    InMux I__9009 (
            .O(N__43242),
            .I(N__43239));
    LocalMux I__9008 (
            .O(N__43239),
            .I(n1797));
    InMux I__9007 (
            .O(N__43236),
            .I(n12594));
    InMux I__9006 (
            .O(N__43233),
            .I(N__43230));
    LocalMux I__9005 (
            .O(N__43230),
            .I(N__43227));
    Odrv4 I__9004 (
            .O(N__43227),
            .I(n1796));
    InMux I__9003 (
            .O(N__43224),
            .I(n12595));
    CascadeMux I__9002 (
            .O(N__43221),
            .I(N__43218));
    InMux I__9001 (
            .O(N__43218),
            .I(N__43215));
    LocalMux I__9000 (
            .O(N__43215),
            .I(N__43212));
    Odrv4 I__8999 (
            .O(N__43212),
            .I(n1795));
    InMux I__8998 (
            .O(N__43209),
            .I(n12596));
    InMux I__8997 (
            .O(N__43206),
            .I(N__43203));
    LocalMux I__8996 (
            .O(N__43203),
            .I(N__43200));
    Odrv12 I__8995 (
            .O(N__43200),
            .I(n1794));
    CascadeMux I__8994 (
            .O(N__43197),
            .I(n1721_cascade_));
    InMux I__8993 (
            .O(N__43194),
            .I(N__43190));
    CascadeMux I__8992 (
            .O(N__43193),
            .I(N__43187));
    LocalMux I__8991 (
            .O(N__43190),
            .I(N__43183));
    InMux I__8990 (
            .O(N__43187),
            .I(N__43180));
    InMux I__8989 (
            .O(N__43186),
            .I(N__43177));
    Odrv4 I__8988 (
            .O(N__43183),
            .I(n1820));
    LocalMux I__8987 (
            .O(N__43180),
            .I(n1820));
    LocalMux I__8986 (
            .O(N__43177),
            .I(n1820));
    CascadeMux I__8985 (
            .O(N__43170),
            .I(N__43166));
    CascadeMux I__8984 (
            .O(N__43169),
            .I(N__43163));
    InMux I__8983 (
            .O(N__43166),
            .I(N__43159));
    InMux I__8982 (
            .O(N__43163),
            .I(N__43156));
    InMux I__8981 (
            .O(N__43162),
            .I(N__43153));
    LocalMux I__8980 (
            .O(N__43159),
            .I(n1827));
    LocalMux I__8979 (
            .O(N__43156),
            .I(n1827));
    LocalMux I__8978 (
            .O(N__43153),
            .I(n1827));
    CascadeMux I__8977 (
            .O(N__43146),
            .I(n1722_cascade_));
    CascadeMux I__8976 (
            .O(N__43143),
            .I(N__43139));
    CascadeMux I__8975 (
            .O(N__43142),
            .I(N__43136));
    InMux I__8974 (
            .O(N__43139),
            .I(N__43132));
    InMux I__8973 (
            .O(N__43136),
            .I(N__43129));
    InMux I__8972 (
            .O(N__43135),
            .I(N__43126));
    LocalMux I__8971 (
            .O(N__43132),
            .I(n1821));
    LocalMux I__8970 (
            .O(N__43129),
            .I(n1821));
    LocalMux I__8969 (
            .O(N__43126),
            .I(n1821));
    CascadeMux I__8968 (
            .O(N__43119),
            .I(N__43116));
    InMux I__8967 (
            .O(N__43116),
            .I(N__43113));
    LocalMux I__8966 (
            .O(N__43113),
            .I(N__43108));
    InMux I__8965 (
            .O(N__43112),
            .I(N__43105));
    CascadeMux I__8964 (
            .O(N__43111),
            .I(N__43102));
    Span4Mux_h I__8963 (
            .O(N__43108),
            .I(N__43099));
    LocalMux I__8962 (
            .O(N__43105),
            .I(N__43096));
    InMux I__8961 (
            .O(N__43102),
            .I(N__43093));
    Odrv4 I__8960 (
            .O(N__43099),
            .I(n1830));
    Odrv4 I__8959 (
            .O(N__43096),
            .I(n1830));
    LocalMux I__8958 (
            .O(N__43093),
            .I(n1830));
    CascadeMux I__8957 (
            .O(N__43086),
            .I(n1752_cascade_));
    InMux I__8956 (
            .O(N__43083),
            .I(N__43079));
    CascadeMux I__8955 (
            .O(N__43082),
            .I(N__43076));
    LocalMux I__8954 (
            .O(N__43079),
            .I(N__43072));
    InMux I__8953 (
            .O(N__43076),
            .I(N__43069));
    InMux I__8952 (
            .O(N__43075),
            .I(N__43066));
    Odrv4 I__8951 (
            .O(N__43072),
            .I(n1826));
    LocalMux I__8950 (
            .O(N__43069),
            .I(n1826));
    LocalMux I__8949 (
            .O(N__43066),
            .I(n1826));
    CascadeMux I__8948 (
            .O(N__43059),
            .I(N__43054));
    CascadeMux I__8947 (
            .O(N__43058),
            .I(N__43051));
    InMux I__8946 (
            .O(N__43057),
            .I(N__43046));
    InMux I__8945 (
            .O(N__43054),
            .I(N__43046));
    InMux I__8944 (
            .O(N__43051),
            .I(N__43043));
    LocalMux I__8943 (
            .O(N__43046),
            .I(N__43040));
    LocalMux I__8942 (
            .O(N__43043),
            .I(n1824));
    Odrv4 I__8941 (
            .O(N__43040),
            .I(n1824));
    CascadeMux I__8940 (
            .O(N__43035),
            .I(N__43032));
    InMux I__8939 (
            .O(N__43032),
            .I(N__43028));
    CascadeMux I__8938 (
            .O(N__43031),
            .I(N__43024));
    LocalMux I__8937 (
            .O(N__43028),
            .I(N__43021));
    InMux I__8936 (
            .O(N__43027),
            .I(N__43018));
    InMux I__8935 (
            .O(N__43024),
            .I(N__43015));
    Span4Mux_h I__8934 (
            .O(N__43021),
            .I(N__43010));
    LocalMux I__8933 (
            .O(N__43018),
            .I(N__43010));
    LocalMux I__8932 (
            .O(N__43015),
            .I(n1823));
    Odrv4 I__8931 (
            .O(N__43010),
            .I(n1823));
    CascadeMux I__8930 (
            .O(N__43005),
            .I(n1726_cascade_));
    CascadeMux I__8929 (
            .O(N__43002),
            .I(n14244_cascade_));
    CascadeMux I__8928 (
            .O(N__42999),
            .I(n14250_cascade_));
    InMux I__8927 (
            .O(N__42996),
            .I(N__42993));
    LocalMux I__8926 (
            .O(N__42993),
            .I(n14254));
    InMux I__8925 (
            .O(N__42990),
            .I(N__42987));
    LocalMux I__8924 (
            .O(N__42987),
            .I(N__42984));
    Odrv12 I__8923 (
            .O(N__42984),
            .I(pwm_setpoint_23_N_171_17));
    InMux I__8922 (
            .O(N__42981),
            .I(N__42972));
    InMux I__8921 (
            .O(N__42980),
            .I(N__42972));
    InMux I__8920 (
            .O(N__42979),
            .I(N__42972));
    LocalMux I__8919 (
            .O(N__42972),
            .I(pwm_setpoint_16));
    CascadeMux I__8918 (
            .O(N__42969),
            .I(N__42966));
    InMux I__8917 (
            .O(N__42966),
            .I(N__42961));
    InMux I__8916 (
            .O(N__42965),
            .I(N__42958));
    InMux I__8915 (
            .O(N__42964),
            .I(N__42955));
    LocalMux I__8914 (
            .O(N__42961),
            .I(N__42952));
    LocalMux I__8913 (
            .O(N__42958),
            .I(N__42947));
    LocalMux I__8912 (
            .O(N__42955),
            .I(N__42947));
    Span4Mux_s3_v I__8911 (
            .O(N__42952),
            .I(N__42942));
    Span4Mux_s3_v I__8910 (
            .O(N__42947),
            .I(N__42942));
    Odrv4 I__8909 (
            .O(N__42942),
            .I(pwm_setpoint_7));
    InMux I__8908 (
            .O(N__42939),
            .I(N__42936));
    LocalMux I__8907 (
            .O(N__42936),
            .I(N__42933));
    Odrv12 I__8906 (
            .O(N__42933),
            .I(pwm_setpoint_23_N_171_10));
    InMux I__8905 (
            .O(N__42930),
            .I(N__42926));
    InMux I__8904 (
            .O(N__42929),
            .I(N__42923));
    LocalMux I__8903 (
            .O(N__42926),
            .I(N__42920));
    LocalMux I__8902 (
            .O(N__42923),
            .I(N__42917));
    Span4Mux_s2_v I__8901 (
            .O(N__42920),
            .I(N__42914));
    Span4Mux_h I__8900 (
            .O(N__42917),
            .I(N__42911));
    Odrv4 I__8899 (
            .O(N__42914),
            .I(pwm_setpoint_11));
    Odrv4 I__8898 (
            .O(N__42911),
            .I(pwm_setpoint_11));
    InMux I__8897 (
            .O(N__42906),
            .I(N__42903));
    LocalMux I__8896 (
            .O(N__42903),
            .I(N__42900));
    Odrv4 I__8895 (
            .O(N__42900),
            .I(n15204));
    InMux I__8894 (
            .O(N__42897),
            .I(N__42891));
    InMux I__8893 (
            .O(N__42896),
            .I(N__42891));
    LocalMux I__8892 (
            .O(N__42891),
            .I(pwm_setpoint_17));
    CascadeMux I__8891 (
            .O(N__42888),
            .I(n35_cascade_));
    InMux I__8890 (
            .O(N__42885),
            .I(N__42882));
    LocalMux I__8889 (
            .O(N__42882),
            .I(n12_adj_661));
    InMux I__8888 (
            .O(N__42879),
            .I(N__42875));
    CascadeMux I__8887 (
            .O(N__42878),
            .I(N__42872));
    LocalMux I__8886 (
            .O(N__42875),
            .I(N__42869));
    InMux I__8885 (
            .O(N__42872),
            .I(N__42866));
    Odrv4 I__8884 (
            .O(N__42869),
            .I(n1825));
    LocalMux I__8883 (
            .O(N__42866),
            .I(n1825));
    CascadeMux I__8882 (
            .O(N__42861),
            .I(n1825_cascade_));
    InMux I__8881 (
            .O(N__42858),
            .I(N__42855));
    LocalMux I__8880 (
            .O(N__42855),
            .I(N__42852));
    Odrv4 I__8879 (
            .O(N__42852),
            .I(n14520));
    InMux I__8878 (
            .O(N__42849),
            .I(N__42845));
    CascadeMux I__8877 (
            .O(N__42848),
            .I(N__42842));
    LocalMux I__8876 (
            .O(N__42845),
            .I(N__42838));
    InMux I__8875 (
            .O(N__42842),
            .I(N__42835));
    InMux I__8874 (
            .O(N__42841),
            .I(N__42832));
    Odrv4 I__8873 (
            .O(N__42838),
            .I(n1828));
    LocalMux I__8872 (
            .O(N__42835),
            .I(n1828));
    LocalMux I__8871 (
            .O(N__42832),
            .I(n1828));
    InMux I__8870 (
            .O(N__42825),
            .I(N__42822));
    LocalMux I__8869 (
            .O(N__42822),
            .I(N__42819));
    Odrv12 I__8868 (
            .O(N__42819),
            .I(pwm_setpoint_23_N_171_22));
    InMux I__8867 (
            .O(N__42816),
            .I(N__42810));
    InMux I__8866 (
            .O(N__42815),
            .I(N__42810));
    LocalMux I__8865 (
            .O(N__42810),
            .I(N__42807));
    Odrv4 I__8864 (
            .O(N__42807),
            .I(n9_adj_658));
    InMux I__8863 (
            .O(N__42804),
            .I(N__42800));
    InMux I__8862 (
            .O(N__42803),
            .I(N__42797));
    LocalMux I__8861 (
            .O(N__42800),
            .I(N__42794));
    LocalMux I__8860 (
            .O(N__42797),
            .I(pwm_setpoint_8));
    Odrv4 I__8859 (
            .O(N__42794),
            .I(pwm_setpoint_8));
    CascadeMux I__8858 (
            .O(N__42789),
            .I(N__42786));
    InMux I__8857 (
            .O(N__42786),
            .I(N__42783));
    LocalMux I__8856 (
            .O(N__42783),
            .I(n17_adj_665));
    InMux I__8855 (
            .O(N__42780),
            .I(N__42774));
    InMux I__8854 (
            .O(N__42779),
            .I(N__42774));
    LocalMux I__8853 (
            .O(N__42774),
            .I(n19_adj_666));
    InMux I__8852 (
            .O(N__42771),
            .I(N__42768));
    LocalMux I__8851 (
            .O(N__42768),
            .I(n15178));
    CascadeMux I__8850 (
            .O(N__42765),
            .I(n17_adj_665_cascade_));
    InMux I__8849 (
            .O(N__42762),
            .I(N__42759));
    LocalMux I__8848 (
            .O(N__42759),
            .I(N__42756));
    Odrv12 I__8847 (
            .O(N__42756),
            .I(pwm_setpoint_23_N_171_16));
    InMux I__8846 (
            .O(N__42753),
            .I(N__42750));
    LocalMux I__8845 (
            .O(N__42750),
            .I(n15174));
    CascadeMux I__8844 (
            .O(N__42747),
            .I(n16_adj_664_cascade_));
    CascadeMux I__8843 (
            .O(N__42744),
            .I(n24_adj_669_cascade_));
    InMux I__8842 (
            .O(N__42741),
            .I(N__42738));
    LocalMux I__8841 (
            .O(N__42738),
            .I(N__42735));
    Span4Mux_v I__8840 (
            .O(N__42735),
            .I(N__42732));
    Odrv4 I__8839 (
            .O(N__42732),
            .I(n8_adj_657));
    InMux I__8838 (
            .O(N__42729),
            .I(N__42726));
    LocalMux I__8837 (
            .O(N__42726),
            .I(n15144));
    InMux I__8836 (
            .O(N__42723),
            .I(N__42720));
    LocalMux I__8835 (
            .O(N__42720),
            .I(pwm_setpoint_23_N_171_21));
    CascadeMux I__8834 (
            .O(N__42717),
            .I(N__42714));
    InMux I__8833 (
            .O(N__42714),
            .I(N__42711));
    LocalMux I__8832 (
            .O(N__42711),
            .I(N__42708));
    Odrv4 I__8831 (
            .O(N__42708),
            .I(pwm_setpoint_23_N_171_9));
    InMux I__8830 (
            .O(N__42705),
            .I(N__42696));
    InMux I__8829 (
            .O(N__42704),
            .I(N__42696));
    InMux I__8828 (
            .O(N__42703),
            .I(N__42696));
    LocalMux I__8827 (
            .O(N__42696),
            .I(pwm_setpoint_9));
    InMux I__8826 (
            .O(N__42693),
            .I(N__42690));
    LocalMux I__8825 (
            .O(N__42690),
            .I(N__42687));
    Odrv4 I__8824 (
            .O(N__42687),
            .I(pwm_setpoint_23_N_171_14));
    InMux I__8823 (
            .O(N__42684),
            .I(N__42681));
    LocalMux I__8822 (
            .O(N__42681),
            .I(N__42678));
    Odrv4 I__8821 (
            .O(N__42678),
            .I(n9_adj_581));
    InMux I__8820 (
            .O(N__42675),
            .I(bfn_11_28_0_));
    InMux I__8819 (
            .O(N__42672),
            .I(n12442));
    InMux I__8818 (
            .O(N__42669),
            .I(N__42666));
    LocalMux I__8817 (
            .O(N__42666),
            .I(N__42663));
    Span4Mux_v I__8816 (
            .O(N__42663),
            .I(N__42660));
    Odrv4 I__8815 (
            .O(N__42660),
            .I(pwm_setpoint_23_N_171_18));
    InMux I__8814 (
            .O(N__42657),
            .I(n12443));
    InMux I__8813 (
            .O(N__42654),
            .I(n12444));
    InMux I__8812 (
            .O(N__42651),
            .I(n12445));
    InMux I__8811 (
            .O(N__42648),
            .I(n12446));
    InMux I__8810 (
            .O(N__42645),
            .I(n12447));
    InMux I__8809 (
            .O(N__42642),
            .I(n12448));
    InMux I__8808 (
            .O(N__42639),
            .I(N__42636));
    LocalMux I__8807 (
            .O(N__42636),
            .I(N__42633));
    Span4Mux_h I__8806 (
            .O(N__42633),
            .I(N__42630));
    Odrv4 I__8805 (
            .O(N__42630),
            .I(n17_adj_589));
    InMux I__8804 (
            .O(N__42627),
            .I(N__42624));
    LocalMux I__8803 (
            .O(N__42624),
            .I(pwm_setpoint_23_N_171_8));
    InMux I__8802 (
            .O(N__42621),
            .I(bfn_11_27_0_));
    InMux I__8801 (
            .O(N__42618),
            .I(N__42615));
    LocalMux I__8800 (
            .O(N__42615),
            .I(N__42612));
    Span4Mux_h I__8799 (
            .O(N__42612),
            .I(N__42609));
    Odrv4 I__8798 (
            .O(N__42609),
            .I(n16_adj_588));
    InMux I__8797 (
            .O(N__42606),
            .I(n12434));
    InMux I__8796 (
            .O(N__42603),
            .I(N__42600));
    LocalMux I__8795 (
            .O(N__42600),
            .I(N__42597));
    Span4Mux_h I__8794 (
            .O(N__42597),
            .I(N__42594));
    Odrv4 I__8793 (
            .O(N__42594),
            .I(n15_adj_587));
    InMux I__8792 (
            .O(N__42591),
            .I(n12435));
    InMux I__8791 (
            .O(N__42588),
            .I(N__42585));
    LocalMux I__8790 (
            .O(N__42585),
            .I(N__42582));
    Span4Mux_h I__8789 (
            .O(N__42582),
            .I(N__42579));
    Odrv4 I__8788 (
            .O(N__42579),
            .I(n14_adj_586));
    InMux I__8787 (
            .O(N__42576),
            .I(N__42573));
    LocalMux I__8786 (
            .O(N__42573),
            .I(pwm_setpoint_23_N_171_11));
    InMux I__8785 (
            .O(N__42570),
            .I(n12436));
    InMux I__8784 (
            .O(N__42567),
            .I(n12437));
    InMux I__8783 (
            .O(N__42564),
            .I(N__42561));
    LocalMux I__8782 (
            .O(N__42561),
            .I(n12_adj_584));
    InMux I__8781 (
            .O(N__42558),
            .I(N__42555));
    LocalMux I__8780 (
            .O(N__42555),
            .I(pwm_setpoint_23_N_171_13));
    InMux I__8779 (
            .O(N__42552),
            .I(n12438));
    InMux I__8778 (
            .O(N__42549),
            .I(N__42546));
    LocalMux I__8777 (
            .O(N__42546),
            .I(N__42543));
    Span4Mux_v I__8776 (
            .O(N__42543),
            .I(N__42540));
    Odrv4 I__8775 (
            .O(N__42540),
            .I(n11_adj_583));
    InMux I__8774 (
            .O(N__42537),
            .I(n12439));
    InMux I__8773 (
            .O(N__42534),
            .I(N__42531));
    LocalMux I__8772 (
            .O(N__42531),
            .I(N__42528));
    Span4Mux_h I__8771 (
            .O(N__42528),
            .I(N__42525));
    Span4Mux_h I__8770 (
            .O(N__42525),
            .I(N__42522));
    Span4Mux_h I__8769 (
            .O(N__42522),
            .I(N__42519));
    Odrv4 I__8768 (
            .O(N__42519),
            .I(n10_adj_582));
    InMux I__8767 (
            .O(N__42516),
            .I(n12440));
    InMux I__8766 (
            .O(N__42513),
            .I(N__42510));
    LocalMux I__8765 (
            .O(N__42510),
            .I(N__42507));
    Odrv12 I__8764 (
            .O(N__42507),
            .I(encoder0_position_scaled_2));
    InMux I__8763 (
            .O(N__42504),
            .I(N__42501));
    LocalMux I__8762 (
            .O(N__42501),
            .I(n25_adj_597));
    InMux I__8761 (
            .O(N__42498),
            .I(bfn_11_26_0_));
    InMux I__8760 (
            .O(N__42495),
            .I(n12426));
    InMux I__8759 (
            .O(N__42492),
            .I(n12427));
    InMux I__8758 (
            .O(N__42489),
            .I(N__42486));
    LocalMux I__8757 (
            .O(N__42486),
            .I(n22_adj_594));
    InMux I__8756 (
            .O(N__42483),
            .I(n12428));
    InMux I__8755 (
            .O(N__42480),
            .I(N__42477));
    LocalMux I__8754 (
            .O(N__42477),
            .I(n21_adj_593));
    InMux I__8753 (
            .O(N__42474),
            .I(N__42471));
    LocalMux I__8752 (
            .O(N__42471),
            .I(pwm_setpoint_23_N_171_4));
    InMux I__8751 (
            .O(N__42468),
            .I(n12429));
    InMux I__8750 (
            .O(N__42465),
            .I(N__42462));
    LocalMux I__8749 (
            .O(N__42462),
            .I(n20_adj_592));
    InMux I__8748 (
            .O(N__42459),
            .I(N__42456));
    LocalMux I__8747 (
            .O(N__42456),
            .I(pwm_setpoint_23_N_171_5));
    InMux I__8746 (
            .O(N__42453),
            .I(n12430));
    InMux I__8745 (
            .O(N__42450),
            .I(n12431));
    InMux I__8744 (
            .O(N__42447),
            .I(N__42444));
    LocalMux I__8743 (
            .O(N__42444),
            .I(n18_adj_590));
    InMux I__8742 (
            .O(N__42441),
            .I(N__42438));
    LocalMux I__8741 (
            .O(N__42438),
            .I(pwm_setpoint_23_N_171_7));
    InMux I__8740 (
            .O(N__42435),
            .I(n12432));
    InMux I__8739 (
            .O(N__42432),
            .I(n12506));
    InMux I__8738 (
            .O(N__42429),
            .I(N__42424));
    InMux I__8737 (
            .O(N__42428),
            .I(N__42421));
    InMux I__8736 (
            .O(N__42427),
            .I(N__42418));
    LocalMux I__8735 (
            .O(N__42424),
            .I(N__42415));
    LocalMux I__8734 (
            .O(N__42421),
            .I(N__42410));
    LocalMux I__8733 (
            .O(N__42418),
            .I(N__42410));
    Span4Mux_h I__8732 (
            .O(N__42415),
            .I(N__42407));
    Span4Mux_h I__8731 (
            .O(N__42410),
            .I(N__42404));
    Odrv4 I__8730 (
            .O(N__42407),
            .I(n2));
    Odrv4 I__8729 (
            .O(N__42404),
            .I(n2));
    CascadeMux I__8728 (
            .O(N__42399),
            .I(N__42396));
    InMux I__8727 (
            .O(N__42396),
            .I(N__42393));
    LocalMux I__8726 (
            .O(N__42393),
            .I(n14568));
    InMux I__8725 (
            .O(N__42390),
            .I(N__42387));
    LocalMux I__8724 (
            .O(N__42387),
            .I(N__42384));
    Odrv4 I__8723 (
            .O(N__42384),
            .I(n2561));
    CascadeMux I__8722 (
            .O(N__42381),
            .I(N__42378));
    InMux I__8721 (
            .O(N__42378),
            .I(N__42374));
    InMux I__8720 (
            .O(N__42377),
            .I(N__42371));
    LocalMux I__8719 (
            .O(N__42374),
            .I(n828));
    LocalMux I__8718 (
            .O(N__42371),
            .I(n828));
    InMux I__8717 (
            .O(N__42366),
            .I(N__42363));
    LocalMux I__8716 (
            .O(N__42363),
            .I(N__42360));
    Odrv12 I__8715 (
            .O(N__42360),
            .I(encoder0_position_scaled_3));
    InMux I__8714 (
            .O(N__42357),
            .I(N__42354));
    LocalMux I__8713 (
            .O(N__42354),
            .I(N__42351));
    Odrv12 I__8712 (
            .O(N__42351),
            .I(encoder0_position_scaled_6));
    InMux I__8711 (
            .O(N__42348),
            .I(N__42344));
    InMux I__8710 (
            .O(N__42347),
            .I(N__42341));
    LocalMux I__8709 (
            .O(N__42344),
            .I(N__42337));
    LocalMux I__8708 (
            .O(N__42341),
            .I(N__42334));
    InMux I__8707 (
            .O(N__42340),
            .I(N__42331));
    Span4Mux_v I__8706 (
            .O(N__42337),
            .I(N__42326));
    Span4Mux_v I__8705 (
            .O(N__42334),
            .I(N__42326));
    LocalMux I__8704 (
            .O(N__42331),
            .I(N__42323));
    Odrv4 I__8703 (
            .O(N__42326),
            .I(n6));
    Odrv4 I__8702 (
            .O(N__42323),
            .I(n6));
    CascadeMux I__8701 (
            .O(N__42318),
            .I(N__42313));
    InMux I__8700 (
            .O(N__42317),
            .I(N__42310));
    InMux I__8699 (
            .O(N__42316),
            .I(N__42307));
    InMux I__8698 (
            .O(N__42313),
            .I(N__42304));
    LocalMux I__8697 (
            .O(N__42310),
            .I(N__42301));
    LocalMux I__8696 (
            .O(N__42307),
            .I(N__42298));
    LocalMux I__8695 (
            .O(N__42304),
            .I(N__42295));
    Span4Mux_h I__8694 (
            .O(N__42301),
            .I(N__42292));
    Span4Mux_h I__8693 (
            .O(N__42298),
            .I(N__42289));
    Odrv4 I__8692 (
            .O(N__42295),
            .I(n4));
    Odrv4 I__8691 (
            .O(N__42292),
            .I(n4));
    Odrv4 I__8690 (
            .O(N__42289),
            .I(n4));
    CascadeMux I__8689 (
            .O(N__42282),
            .I(N__42278));
    CascadeMux I__8688 (
            .O(N__42281),
            .I(N__42275));
    InMux I__8687 (
            .O(N__42278),
            .I(N__42272));
    InMux I__8686 (
            .O(N__42275),
            .I(N__42269));
    LocalMux I__8685 (
            .O(N__42272),
            .I(n40));
    LocalMux I__8684 (
            .O(N__42269),
            .I(n40));
    InMux I__8683 (
            .O(N__42264),
            .I(N__42260));
    InMux I__8682 (
            .O(N__42263),
            .I(N__42257));
    LocalMux I__8681 (
            .O(N__42260),
            .I(N__42253));
    LocalMux I__8680 (
            .O(N__42257),
            .I(N__42250));
    InMux I__8679 (
            .O(N__42256),
            .I(N__42247));
    Span4Mux_v I__8678 (
            .O(N__42253),
            .I(N__42244));
    Span4Mux_h I__8677 (
            .O(N__42250),
            .I(N__42241));
    LocalMux I__8676 (
            .O(N__42247),
            .I(N__42238));
    Odrv4 I__8675 (
            .O(N__42244),
            .I(n5));
    Odrv4 I__8674 (
            .O(N__42241),
            .I(n5));
    Odrv4 I__8673 (
            .O(N__42238),
            .I(n5));
    InMux I__8672 (
            .O(N__42231),
            .I(N__42228));
    LocalMux I__8671 (
            .O(N__42228),
            .I(n5_adj_682));
    CascadeMux I__8670 (
            .O(N__42225),
            .I(N__42222));
    InMux I__8669 (
            .O(N__42222),
            .I(N__42212));
    InMux I__8668 (
            .O(N__42221),
            .I(N__42212));
    InMux I__8667 (
            .O(N__42220),
            .I(N__42212));
    InMux I__8666 (
            .O(N__42219),
            .I(N__42209));
    LocalMux I__8665 (
            .O(N__42212),
            .I(N__42204));
    LocalMux I__8664 (
            .O(N__42209),
            .I(N__42204));
    Span4Mux_h I__8663 (
            .O(N__42204),
            .I(N__42201));
    Odrv4 I__8662 (
            .O(N__42201),
            .I(n3));
    CascadeMux I__8661 (
            .O(N__42198),
            .I(n5_adj_682_cascade_));
    CascadeMux I__8660 (
            .O(N__42195),
            .I(N__42190));
    InMux I__8659 (
            .O(N__42194),
            .I(N__42185));
    InMux I__8658 (
            .O(N__42193),
            .I(N__42182));
    InMux I__8657 (
            .O(N__42190),
            .I(N__42175));
    InMux I__8656 (
            .O(N__42189),
            .I(N__42175));
    InMux I__8655 (
            .O(N__42188),
            .I(N__42175));
    LocalMux I__8654 (
            .O(N__42185),
            .I(n13653));
    LocalMux I__8653 (
            .O(N__42182),
            .I(n13653));
    LocalMux I__8652 (
            .O(N__42175),
            .I(n13653));
    InMux I__8651 (
            .O(N__42168),
            .I(bfn_11_24_0_));
    InMux I__8650 (
            .O(N__42165),
            .I(n12501));
    InMux I__8649 (
            .O(N__42162),
            .I(n12502));
    CascadeMux I__8648 (
            .O(N__42159),
            .I(N__42156));
    InMux I__8647 (
            .O(N__42156),
            .I(N__42152));
    InMux I__8646 (
            .O(N__42155),
            .I(N__42148));
    LocalMux I__8645 (
            .O(N__42152),
            .I(N__42145));
    InMux I__8644 (
            .O(N__42151),
            .I(N__42142));
    LocalMux I__8643 (
            .O(N__42148),
            .I(n831));
    Odrv4 I__8642 (
            .O(N__42145),
            .I(n831));
    LocalMux I__8641 (
            .O(N__42142),
            .I(n831));
    InMux I__8640 (
            .O(N__42135),
            .I(N__42132));
    LocalMux I__8639 (
            .O(N__42132),
            .I(n898));
    InMux I__8638 (
            .O(N__42129),
            .I(n12503));
    CascadeMux I__8637 (
            .O(N__42126),
            .I(N__42122));
    CascadeMux I__8636 (
            .O(N__42125),
            .I(N__42119));
    InMux I__8635 (
            .O(N__42122),
            .I(N__42115));
    InMux I__8634 (
            .O(N__42119),
            .I(N__42112));
    InMux I__8633 (
            .O(N__42118),
            .I(N__42109));
    LocalMux I__8632 (
            .O(N__42115),
            .I(N__42106));
    LocalMux I__8631 (
            .O(N__42112),
            .I(n830));
    LocalMux I__8630 (
            .O(N__42109),
            .I(n830));
    Odrv4 I__8629 (
            .O(N__42106),
            .I(n830));
    InMux I__8628 (
            .O(N__42099),
            .I(N__42096));
    LocalMux I__8627 (
            .O(N__42096),
            .I(n897));
    InMux I__8626 (
            .O(N__42093),
            .I(n12504));
    InMux I__8625 (
            .O(N__42090),
            .I(n12505));
    CascadeMux I__8624 (
            .O(N__42087),
            .I(n832_cascade_));
    InMux I__8623 (
            .O(N__42084),
            .I(N__42081));
    LocalMux I__8622 (
            .O(N__42081),
            .I(n2564));
    CascadeMux I__8621 (
            .O(N__42078),
            .I(n13658_cascade_));
    CascadeMux I__8620 (
            .O(N__42075),
            .I(N__42070));
    CascadeMux I__8619 (
            .O(N__42074),
            .I(N__42067));
    CascadeMux I__8618 (
            .O(N__42073),
            .I(N__42064));
    InMux I__8617 (
            .O(N__42070),
            .I(N__42060));
    InMux I__8616 (
            .O(N__42067),
            .I(N__42057));
    InMux I__8615 (
            .O(N__42064),
            .I(N__42054));
    InMux I__8614 (
            .O(N__42063),
            .I(N__42051));
    LocalMux I__8613 (
            .O(N__42060),
            .I(N__42048));
    LocalMux I__8612 (
            .O(N__42057),
            .I(N__42045));
    LocalMux I__8611 (
            .O(N__42054),
            .I(encoder0_position_28));
    LocalMux I__8610 (
            .O(N__42051),
            .I(encoder0_position_28));
    Odrv4 I__8609 (
            .O(N__42048),
            .I(encoder0_position_28));
    Odrv12 I__8608 (
            .O(N__42045),
            .I(encoder0_position_28));
    InMux I__8607 (
            .O(N__42036),
            .I(N__42033));
    LocalMux I__8606 (
            .O(N__42033),
            .I(N__42030));
    Span4Mux_v I__8605 (
            .O(N__42030),
            .I(N__42027));
    Odrv4 I__8604 (
            .O(N__42027),
            .I(encoder0_position_scaled_4));
    CascadeMux I__8603 (
            .O(N__42024),
            .I(n929_cascade_));
    CascadeMux I__8602 (
            .O(N__42021),
            .I(N__42016));
    CascadeMux I__8601 (
            .O(N__42020),
            .I(N__42013));
    CascadeMux I__8600 (
            .O(N__42019),
            .I(N__42010));
    InMux I__8599 (
            .O(N__42016),
            .I(N__42007));
    InMux I__8598 (
            .O(N__42013),
            .I(N__42004));
    InMux I__8597 (
            .O(N__42010),
            .I(N__42000));
    LocalMux I__8596 (
            .O(N__42007),
            .I(N__41995));
    LocalMux I__8595 (
            .O(N__42004),
            .I(N__41995));
    InMux I__8594 (
            .O(N__42003),
            .I(N__41992));
    LocalMux I__8593 (
            .O(N__42000),
            .I(encoder0_position_30));
    Odrv4 I__8592 (
            .O(N__41995),
            .I(encoder0_position_30));
    LocalMux I__8591 (
            .O(N__41992),
            .I(encoder0_position_30));
    InMux I__8590 (
            .O(N__41985),
            .I(N__41982));
    LocalMux I__8589 (
            .O(N__41982),
            .I(n13654));
    CascadeMux I__8588 (
            .O(N__41979),
            .I(n829_cascade_));
    InMux I__8587 (
            .O(N__41976),
            .I(N__41973));
    LocalMux I__8586 (
            .O(N__41973),
            .I(n12027));
    CascadeMux I__8585 (
            .O(N__41970),
            .I(n861_cascade_));
    InMux I__8584 (
            .O(N__41967),
            .I(N__41964));
    LocalMux I__8583 (
            .O(N__41964),
            .I(N__41961));
    Span4Mux_h I__8582 (
            .O(N__41961),
            .I(N__41958));
    Odrv4 I__8581 (
            .O(N__41958),
            .I(n16));
    CascadeMux I__8580 (
            .O(N__41955),
            .I(N__41951));
    InMux I__8579 (
            .O(N__41954),
            .I(N__41946));
    InMux I__8578 (
            .O(N__41951),
            .I(N__41943));
    InMux I__8577 (
            .O(N__41950),
            .I(N__41940));
    InMux I__8576 (
            .O(N__41949),
            .I(N__41937));
    LocalMux I__8575 (
            .O(N__41946),
            .I(encoder0_position_29));
    LocalMux I__8574 (
            .O(N__41943),
            .I(encoder0_position_29));
    LocalMux I__8573 (
            .O(N__41940),
            .I(encoder0_position_29));
    LocalMux I__8572 (
            .O(N__41937),
            .I(encoder0_position_29));
    CascadeMux I__8571 (
            .O(N__41928),
            .I(N__41925));
    InMux I__8570 (
            .O(N__41925),
            .I(N__41922));
    LocalMux I__8569 (
            .O(N__41922),
            .I(n404));
    InMux I__8568 (
            .O(N__41919),
            .I(N__41914));
    InMux I__8567 (
            .O(N__41918),
            .I(N__41909));
    InMux I__8566 (
            .O(N__41917),
            .I(N__41909));
    LocalMux I__8565 (
            .O(N__41914),
            .I(encoder0_position_17));
    LocalMux I__8564 (
            .O(N__41909),
            .I(encoder0_position_17));
    CascadeMux I__8563 (
            .O(N__41904),
            .I(N__41901));
    InMux I__8562 (
            .O(N__41901),
            .I(N__41898));
    LocalMux I__8561 (
            .O(N__41898),
            .I(N__41895));
    Span4Mux_h I__8560 (
            .O(N__41895),
            .I(N__41892));
    Odrv4 I__8559 (
            .O(N__41892),
            .I(n16_adj_634));
    CascadeMux I__8558 (
            .O(N__41889),
            .I(N__41886));
    InMux I__8557 (
            .O(N__41886),
            .I(N__41883));
    LocalMux I__8556 (
            .O(N__41883),
            .I(N__41880));
    Span4Mux_v I__8555 (
            .O(N__41880),
            .I(N__41877));
    Odrv4 I__8554 (
            .O(N__41877),
            .I(n7_adj_625));
    CascadeMux I__8553 (
            .O(N__41874),
            .I(N__41871));
    InMux I__8552 (
            .O(N__41871),
            .I(N__41868));
    LocalMux I__8551 (
            .O(N__41868),
            .I(N__41865));
    Span4Mux_v I__8550 (
            .O(N__41865),
            .I(N__41862));
    Odrv4 I__8549 (
            .O(N__41862),
            .I(n3_adj_621));
    InMux I__8548 (
            .O(N__41859),
            .I(N__41856));
    LocalMux I__8547 (
            .O(N__41856),
            .I(n2566));
    CascadeMux I__8546 (
            .O(N__41853),
            .I(N__41850));
    InMux I__8545 (
            .O(N__41850),
            .I(N__41847));
    LocalMux I__8544 (
            .O(N__41847),
            .I(N__41843));
    InMux I__8543 (
            .O(N__41846),
            .I(N__41840));
    Span4Mux_h I__8542 (
            .O(N__41843),
            .I(N__41835));
    LocalMux I__8541 (
            .O(N__41840),
            .I(N__41835));
    Odrv4 I__8540 (
            .O(N__41835),
            .I(n7));
    CascadeMux I__8539 (
            .O(N__41832),
            .I(n13662_cascade_));
    CascadeMux I__8538 (
            .O(N__41829),
            .I(N__41825));
    CascadeMux I__8537 (
            .O(N__41828),
            .I(N__41822));
    InMux I__8536 (
            .O(N__41825),
            .I(N__41818));
    InMux I__8535 (
            .O(N__41822),
            .I(N__41814));
    InMux I__8534 (
            .O(N__41821),
            .I(N__41811));
    LocalMux I__8533 (
            .O(N__41818),
            .I(N__41808));
    InMux I__8532 (
            .O(N__41817),
            .I(N__41805));
    LocalMux I__8531 (
            .O(N__41814),
            .I(encoder0_position_26));
    LocalMux I__8530 (
            .O(N__41811),
            .I(encoder0_position_26));
    Odrv4 I__8529 (
            .O(N__41808),
            .I(encoder0_position_26));
    LocalMux I__8528 (
            .O(N__41805),
            .I(encoder0_position_26));
    CascadeMux I__8527 (
            .O(N__41796),
            .I(N__41793));
    InMux I__8526 (
            .O(N__41793),
            .I(N__41790));
    LocalMux I__8525 (
            .O(N__41790),
            .I(n2565));
    InMux I__8524 (
            .O(N__41787),
            .I(N__41781));
    InMux I__8523 (
            .O(N__41786),
            .I(N__41778));
    InMux I__8522 (
            .O(N__41785),
            .I(N__41775));
    InMux I__8521 (
            .O(N__41784),
            .I(N__41772));
    LocalMux I__8520 (
            .O(N__41781),
            .I(N__41767));
    LocalMux I__8519 (
            .O(N__41778),
            .I(N__41767));
    LocalMux I__8518 (
            .O(N__41775),
            .I(encoder0_position_27));
    LocalMux I__8517 (
            .O(N__41772),
            .I(encoder0_position_27));
    Odrv4 I__8516 (
            .O(N__41767),
            .I(encoder0_position_27));
    CascadeMux I__8515 (
            .O(N__41760),
            .I(n13660_cascade_));
    CascadeMux I__8514 (
            .O(N__41757),
            .I(N__41754));
    InMux I__8513 (
            .O(N__41754),
            .I(N__41751));
    LocalMux I__8512 (
            .O(N__41751),
            .I(N__41748));
    Odrv4 I__8511 (
            .O(N__41748),
            .I(n1895));
    CascadeMux I__8510 (
            .O(N__41745),
            .I(N__41741));
    CascadeMux I__8509 (
            .O(N__41744),
            .I(N__41738));
    InMux I__8508 (
            .O(N__41741),
            .I(N__41735));
    InMux I__8507 (
            .O(N__41738),
            .I(N__41732));
    LocalMux I__8506 (
            .O(N__41735),
            .I(N__41729));
    LocalMux I__8505 (
            .O(N__41732),
            .I(N__41726));
    Span4Mux_h I__8504 (
            .O(N__41729),
            .I(N__41720));
    Span4Mux_v I__8503 (
            .O(N__41726),
            .I(N__41720));
    InMux I__8502 (
            .O(N__41725),
            .I(N__41717));
    Odrv4 I__8501 (
            .O(N__41720),
            .I(n1927));
    LocalMux I__8500 (
            .O(N__41717),
            .I(n1927));
    InMux I__8499 (
            .O(N__41712),
            .I(N__41709));
    LocalMux I__8498 (
            .O(N__41709),
            .I(N__41706));
    Odrv4 I__8497 (
            .O(N__41706),
            .I(n1894));
    CascadeMux I__8496 (
            .O(N__41703),
            .I(N__41699));
    CascadeMux I__8495 (
            .O(N__41702),
            .I(N__41696));
    InMux I__8494 (
            .O(N__41699),
            .I(N__41693));
    InMux I__8493 (
            .O(N__41696),
            .I(N__41690));
    LocalMux I__8492 (
            .O(N__41693),
            .I(N__41687));
    LocalMux I__8491 (
            .O(N__41690),
            .I(N__41684));
    Span4Mux_h I__8490 (
            .O(N__41687),
            .I(N__41680));
    Span4Mux_h I__8489 (
            .O(N__41684),
            .I(N__41677));
    InMux I__8488 (
            .O(N__41683),
            .I(N__41674));
    Odrv4 I__8487 (
            .O(N__41680),
            .I(n1926));
    Odrv4 I__8486 (
            .O(N__41677),
            .I(n1926));
    LocalMux I__8485 (
            .O(N__41674),
            .I(n1926));
    CascadeMux I__8484 (
            .O(N__41667),
            .I(N__41662));
    InMux I__8483 (
            .O(N__41666),
            .I(N__41657));
    InMux I__8482 (
            .O(N__41665),
            .I(N__41657));
    InMux I__8481 (
            .O(N__41662),
            .I(N__41654));
    LocalMux I__8480 (
            .O(N__41657),
            .I(N__41649));
    LocalMux I__8479 (
            .O(N__41654),
            .I(N__41649));
    Odrv4 I__8478 (
            .O(N__41649),
            .I(n1829));
    CascadeMux I__8477 (
            .O(N__41646),
            .I(N__41643));
    InMux I__8476 (
            .O(N__41643),
            .I(N__41640));
    LocalMux I__8475 (
            .O(N__41640),
            .I(n1885));
    InMux I__8474 (
            .O(N__41637),
            .I(N__41633));
    InMux I__8473 (
            .O(N__41636),
            .I(N__41630));
    LocalMux I__8472 (
            .O(N__41633),
            .I(N__41627));
    LocalMux I__8471 (
            .O(N__41630),
            .I(N__41624));
    Span4Mux_v I__8470 (
            .O(N__41627),
            .I(N__41621));
    Span4Mux_v I__8469 (
            .O(N__41624),
            .I(N__41618));
    Odrv4 I__8468 (
            .O(N__41621),
            .I(n1917));
    Odrv4 I__8467 (
            .O(N__41618),
            .I(n1917));
    InMux I__8466 (
            .O(N__41613),
            .I(N__41610));
    LocalMux I__8465 (
            .O(N__41610),
            .I(N__41607));
    Span4Mux_v I__8464 (
            .O(N__41607),
            .I(N__41604));
    Odrv4 I__8463 (
            .O(N__41604),
            .I(n30));
    CascadeMux I__8462 (
            .O(N__41601),
            .I(N__41597));
    CascadeMux I__8461 (
            .O(N__41600),
            .I(N__41593));
    InMux I__8460 (
            .O(N__41597),
            .I(N__41590));
    InMux I__8459 (
            .O(N__41596),
            .I(N__41587));
    InMux I__8458 (
            .O(N__41593),
            .I(N__41584));
    LocalMux I__8457 (
            .O(N__41590),
            .I(N__41581));
    LocalMux I__8456 (
            .O(N__41587),
            .I(N__41578));
    LocalMux I__8455 (
            .O(N__41584),
            .I(encoder0_position_3));
    Odrv4 I__8454 (
            .O(N__41581),
            .I(encoder0_position_3));
    Odrv4 I__8453 (
            .O(N__41578),
            .I(encoder0_position_3));
    InMux I__8452 (
            .O(N__41571),
            .I(N__41567));
    InMux I__8451 (
            .O(N__41570),
            .I(N__41564));
    LocalMux I__8450 (
            .O(N__41567),
            .I(N__41560));
    LocalMux I__8449 (
            .O(N__41564),
            .I(N__41557));
    InMux I__8448 (
            .O(N__41563),
            .I(N__41554));
    Span4Mux_v I__8447 (
            .O(N__41560),
            .I(N__41551));
    Span4Mux_s3_h I__8446 (
            .O(N__41557),
            .I(N__41546));
    LocalMux I__8445 (
            .O(N__41554),
            .I(N__41546));
    Span4Mux_h I__8444 (
            .O(N__41551),
            .I(N__41541));
    Span4Mux_h I__8443 (
            .O(N__41546),
            .I(N__41541));
    Span4Mux_v I__8442 (
            .O(N__41541),
            .I(N__41538));
    Span4Mux_v I__8441 (
            .O(N__41538),
            .I(N__41535));
    Odrv4 I__8440 (
            .O(N__41535),
            .I(n316));
    InMux I__8439 (
            .O(N__41532),
            .I(N__41529));
    LocalMux I__8438 (
            .O(N__41529),
            .I(N__41526));
    Odrv4 I__8437 (
            .O(N__41526),
            .I(n1888));
    InMux I__8436 (
            .O(N__41523),
            .I(N__41520));
    LocalMux I__8435 (
            .O(N__41520),
            .I(N__41516));
    InMux I__8434 (
            .O(N__41519),
            .I(N__41509));
    Span4Mux_v I__8433 (
            .O(N__41516),
            .I(N__41506));
    InMux I__8432 (
            .O(N__41515),
            .I(N__41498));
    CascadeMux I__8431 (
            .O(N__41514),
            .I(N__41491));
    CascadeMux I__8430 (
            .O(N__41513),
            .I(N__41486));
    CascadeMux I__8429 (
            .O(N__41512),
            .I(N__41483));
    LocalMux I__8428 (
            .O(N__41509),
            .I(N__41477));
    Span4Mux_v I__8427 (
            .O(N__41506),
            .I(N__41477));
    InMux I__8426 (
            .O(N__41505),
            .I(N__41472));
    InMux I__8425 (
            .O(N__41504),
            .I(N__41472));
    InMux I__8424 (
            .O(N__41503),
            .I(N__41465));
    InMux I__8423 (
            .O(N__41502),
            .I(N__41465));
    InMux I__8422 (
            .O(N__41501),
            .I(N__41465));
    LocalMux I__8421 (
            .O(N__41498),
            .I(N__41462));
    InMux I__8420 (
            .O(N__41497),
            .I(N__41455));
    InMux I__8419 (
            .O(N__41496),
            .I(N__41455));
    InMux I__8418 (
            .O(N__41495),
            .I(N__41455));
    InMux I__8417 (
            .O(N__41494),
            .I(N__41446));
    InMux I__8416 (
            .O(N__41491),
            .I(N__41446));
    InMux I__8415 (
            .O(N__41490),
            .I(N__41446));
    InMux I__8414 (
            .O(N__41489),
            .I(N__41446));
    InMux I__8413 (
            .O(N__41486),
            .I(N__41439));
    InMux I__8412 (
            .O(N__41483),
            .I(N__41439));
    InMux I__8411 (
            .O(N__41482),
            .I(N__41439));
    Span4Mux_h I__8410 (
            .O(N__41477),
            .I(N__41432));
    LocalMux I__8409 (
            .O(N__41472),
            .I(N__41432));
    LocalMux I__8408 (
            .O(N__41465),
            .I(N__41432));
    Odrv4 I__8407 (
            .O(N__41462),
            .I(n1851));
    LocalMux I__8406 (
            .O(N__41455),
            .I(n1851));
    LocalMux I__8405 (
            .O(N__41446),
            .I(n1851));
    LocalMux I__8404 (
            .O(N__41439),
            .I(n1851));
    Odrv4 I__8403 (
            .O(N__41432),
            .I(n1851));
    InMux I__8402 (
            .O(N__41421),
            .I(N__41417));
    InMux I__8401 (
            .O(N__41420),
            .I(N__41414));
    LocalMux I__8400 (
            .O(N__41417),
            .I(N__41411));
    LocalMux I__8399 (
            .O(N__41414),
            .I(N__41408));
    Span4Mux_h I__8398 (
            .O(N__41411),
            .I(N__41405));
    Span4Mux_h I__8397 (
            .O(N__41408),
            .I(N__41402));
    Odrv4 I__8396 (
            .O(N__41405),
            .I(n1920));
    Odrv4 I__8395 (
            .O(N__41402),
            .I(n1920));
    InMux I__8394 (
            .O(N__41397),
            .I(N__41394));
    LocalMux I__8393 (
            .O(N__41394),
            .I(N__41391));
    Span4Mux_h I__8392 (
            .O(N__41391),
            .I(N__41388));
    Odrv4 I__8391 (
            .O(N__41388),
            .I(n1987));
    CascadeMux I__8390 (
            .O(N__41385),
            .I(n1920_cascade_));
    InMux I__8389 (
            .O(N__41382),
            .I(N__41379));
    LocalMux I__8388 (
            .O(N__41379),
            .I(N__41375));
    InMux I__8387 (
            .O(N__41378),
            .I(N__41371));
    Span4Mux_v I__8386 (
            .O(N__41375),
            .I(N__41363));
    InMux I__8385 (
            .O(N__41374),
            .I(N__41360));
    LocalMux I__8384 (
            .O(N__41371),
            .I(N__41353));
    InMux I__8383 (
            .O(N__41370),
            .I(N__41350));
    CascadeMux I__8382 (
            .O(N__41369),
            .I(N__41347));
    CascadeMux I__8381 (
            .O(N__41368),
            .I(N__41344));
    CascadeMux I__8380 (
            .O(N__41367),
            .I(N__41337));
    CascadeMux I__8379 (
            .O(N__41366),
            .I(N__41334));
    Span4Mux_v I__8378 (
            .O(N__41363),
            .I(N__41327));
    LocalMux I__8377 (
            .O(N__41360),
            .I(N__41327));
    InMux I__8376 (
            .O(N__41359),
            .I(N__41324));
    InMux I__8375 (
            .O(N__41358),
            .I(N__41317));
    InMux I__8374 (
            .O(N__41357),
            .I(N__41317));
    InMux I__8373 (
            .O(N__41356),
            .I(N__41317));
    Span4Mux_h I__8372 (
            .O(N__41353),
            .I(N__41314));
    LocalMux I__8371 (
            .O(N__41350),
            .I(N__41311));
    InMux I__8370 (
            .O(N__41347),
            .I(N__41298));
    InMux I__8369 (
            .O(N__41344),
            .I(N__41298));
    InMux I__8368 (
            .O(N__41343),
            .I(N__41298));
    InMux I__8367 (
            .O(N__41342),
            .I(N__41298));
    InMux I__8366 (
            .O(N__41341),
            .I(N__41298));
    InMux I__8365 (
            .O(N__41340),
            .I(N__41298));
    InMux I__8364 (
            .O(N__41337),
            .I(N__41289));
    InMux I__8363 (
            .O(N__41334),
            .I(N__41289));
    InMux I__8362 (
            .O(N__41333),
            .I(N__41289));
    InMux I__8361 (
            .O(N__41332),
            .I(N__41289));
    Odrv4 I__8360 (
            .O(N__41327),
            .I(n1950));
    LocalMux I__8359 (
            .O(N__41324),
            .I(n1950));
    LocalMux I__8358 (
            .O(N__41317),
            .I(n1950));
    Odrv4 I__8357 (
            .O(N__41314),
            .I(n1950));
    Odrv4 I__8356 (
            .O(N__41311),
            .I(n1950));
    LocalMux I__8355 (
            .O(N__41298),
            .I(n1950));
    LocalMux I__8354 (
            .O(N__41289),
            .I(n1950));
    CascadeMux I__8353 (
            .O(N__41274),
            .I(N__41269));
    CascadeMux I__8352 (
            .O(N__41273),
            .I(N__41266));
    CascadeMux I__8351 (
            .O(N__41272),
            .I(N__41263));
    InMux I__8350 (
            .O(N__41269),
            .I(N__41260));
    InMux I__8349 (
            .O(N__41266),
            .I(N__41257));
    InMux I__8348 (
            .O(N__41263),
            .I(N__41254));
    LocalMux I__8347 (
            .O(N__41260),
            .I(N__41251));
    LocalMux I__8346 (
            .O(N__41257),
            .I(N__41248));
    LocalMux I__8345 (
            .O(N__41254),
            .I(N__41245));
    Span4Mux_v I__8344 (
            .O(N__41251),
            .I(N__41240));
    Span4Mux_h I__8343 (
            .O(N__41248),
            .I(N__41240));
    Span4Mux_h I__8342 (
            .O(N__41245),
            .I(N__41237));
    Span4Mux_h I__8341 (
            .O(N__41240),
            .I(N__41234));
    Odrv4 I__8340 (
            .O(N__41237),
            .I(n2019));
    Odrv4 I__8339 (
            .O(N__41234),
            .I(n2019));
    InMux I__8338 (
            .O(N__41229),
            .I(N__41224));
    CascadeMux I__8337 (
            .O(N__41228),
            .I(N__41221));
    InMux I__8336 (
            .O(N__41227),
            .I(N__41218));
    LocalMux I__8335 (
            .O(N__41224),
            .I(N__41215));
    InMux I__8334 (
            .O(N__41221),
            .I(N__41212));
    LocalMux I__8333 (
            .O(N__41218),
            .I(N__41209));
    Span4Mux_h I__8332 (
            .O(N__41215),
            .I(N__41206));
    LocalMux I__8331 (
            .O(N__41212),
            .I(N__41203));
    Span4Mux_h I__8330 (
            .O(N__41209),
            .I(N__41200));
    Odrv4 I__8329 (
            .O(N__41206),
            .I(n1819));
    Odrv4 I__8328 (
            .O(N__41203),
            .I(n1819));
    Odrv4 I__8327 (
            .O(N__41200),
            .I(n1819));
    CascadeMux I__8326 (
            .O(N__41193),
            .I(N__41190));
    InMux I__8325 (
            .O(N__41190),
            .I(N__41187));
    LocalMux I__8324 (
            .O(N__41187),
            .I(N__41184));
    Odrv4 I__8323 (
            .O(N__41184),
            .I(n1889));
    InMux I__8322 (
            .O(N__41181),
            .I(n12617));
    InMux I__8321 (
            .O(N__41178),
            .I(n12618));
    CascadeMux I__8320 (
            .O(N__41175),
            .I(N__41172));
    InMux I__8319 (
            .O(N__41172),
            .I(N__41169));
    LocalMux I__8318 (
            .O(N__41169),
            .I(N__41166));
    Odrv4 I__8317 (
            .O(N__41166),
            .I(n1887));
    InMux I__8316 (
            .O(N__41163),
            .I(n12619));
    CascadeMux I__8315 (
            .O(N__41160),
            .I(N__41157));
    InMux I__8314 (
            .O(N__41157),
            .I(N__41154));
    LocalMux I__8313 (
            .O(N__41154),
            .I(N__41151));
    Odrv4 I__8312 (
            .O(N__41151),
            .I(n1886));
    InMux I__8311 (
            .O(N__41148),
            .I(n12620));
    InMux I__8310 (
            .O(N__41145),
            .I(bfn_11_19_0_));
    CascadeMux I__8309 (
            .O(N__41142),
            .I(N__41139));
    InMux I__8308 (
            .O(N__41139),
            .I(N__41136));
    LocalMux I__8307 (
            .O(N__41136),
            .I(n1892));
    CascadeMux I__8306 (
            .O(N__41133),
            .I(N__41129));
    CascadeMux I__8305 (
            .O(N__41132),
            .I(N__41126));
    InMux I__8304 (
            .O(N__41129),
            .I(N__41123));
    InMux I__8303 (
            .O(N__41126),
            .I(N__41120));
    LocalMux I__8302 (
            .O(N__41123),
            .I(N__41117));
    LocalMux I__8301 (
            .O(N__41120),
            .I(N__41114));
    Span4Mux_h I__8300 (
            .O(N__41117),
            .I(N__41111));
    Odrv12 I__8299 (
            .O(N__41114),
            .I(n1924));
    Odrv4 I__8298 (
            .O(N__41111),
            .I(n1924));
    CascadeMux I__8297 (
            .O(N__41106),
            .I(n1924_cascade_));
    InMux I__8296 (
            .O(N__41103),
            .I(N__41100));
    LocalMux I__8295 (
            .O(N__41100),
            .I(N__41097));
    Span4Mux_h I__8294 (
            .O(N__41097),
            .I(N__41094));
    Odrv4 I__8293 (
            .O(N__41094),
            .I(n14438));
    InMux I__8292 (
            .O(N__41091),
            .I(N__41088));
    LocalMux I__8291 (
            .O(N__41088),
            .I(N__41084));
    CascadeMux I__8290 (
            .O(N__41087),
            .I(N__41081));
    Span4Mux_h I__8289 (
            .O(N__41084),
            .I(N__41078));
    InMux I__8288 (
            .O(N__41081),
            .I(N__41075));
    Odrv4 I__8287 (
            .O(N__41078),
            .I(n1822));
    LocalMux I__8286 (
            .O(N__41075),
            .I(n1822));
    CascadeMux I__8285 (
            .O(N__41070),
            .I(n1822_cascade_));
    InMux I__8284 (
            .O(N__41067),
            .I(N__41064));
    LocalMux I__8283 (
            .O(N__41064),
            .I(N__41061));
    Odrv4 I__8282 (
            .O(N__41061),
            .I(n14534));
    InMux I__8281 (
            .O(N__41058),
            .I(n12608));
    InMux I__8280 (
            .O(N__41055),
            .I(N__41052));
    LocalMux I__8279 (
            .O(N__41052),
            .I(n1897));
    InMux I__8278 (
            .O(N__41049),
            .I(n12609));
    InMux I__8277 (
            .O(N__41046),
            .I(N__41043));
    LocalMux I__8276 (
            .O(N__41043),
            .I(n1896));
    InMux I__8275 (
            .O(N__41040),
            .I(n12610));
    InMux I__8274 (
            .O(N__41037),
            .I(n12611));
    InMux I__8273 (
            .O(N__41034),
            .I(n12612));
    InMux I__8272 (
            .O(N__41031),
            .I(N__41028));
    LocalMux I__8271 (
            .O(N__41028),
            .I(n1893));
    InMux I__8270 (
            .O(N__41025),
            .I(bfn_11_18_0_));
    InMux I__8269 (
            .O(N__41022),
            .I(n12614));
    CascadeMux I__8268 (
            .O(N__41019),
            .I(N__41016));
    InMux I__8267 (
            .O(N__41016),
            .I(N__41013));
    LocalMux I__8266 (
            .O(N__41013),
            .I(n1891));
    InMux I__8265 (
            .O(N__41010),
            .I(n12615));
    InMux I__8264 (
            .O(N__41007),
            .I(N__41004));
    LocalMux I__8263 (
            .O(N__41004),
            .I(N__41001));
    Span4Mux_v I__8262 (
            .O(N__41001),
            .I(N__40998));
    Odrv4 I__8261 (
            .O(N__40998),
            .I(n1890));
    InMux I__8260 (
            .O(N__40995),
            .I(n12616));
    InMux I__8259 (
            .O(N__40992),
            .I(N__40985));
    InMux I__8258 (
            .O(N__40991),
            .I(N__40985));
    InMux I__8257 (
            .O(N__40990),
            .I(N__40982));
    LocalMux I__8256 (
            .O(N__40985),
            .I(blink_counter_24));
    LocalMux I__8255 (
            .O(N__40982),
            .I(blink_counter_24));
    InMux I__8254 (
            .O(N__40977),
            .I(bfn_10_32_0_));
    InMux I__8253 (
            .O(N__40974),
            .I(n13094));
    InMux I__8252 (
            .O(N__40971),
            .I(N__40967));
    InMux I__8251 (
            .O(N__40970),
            .I(N__40964));
    LocalMux I__8250 (
            .O(N__40967),
            .I(blink_counter_25));
    LocalMux I__8249 (
            .O(N__40964),
            .I(blink_counter_25));
    CascadeMux I__8248 (
            .O(N__40959),
            .I(n1833_cascade_));
    InMux I__8247 (
            .O(N__40956),
            .I(N__40953));
    LocalMux I__8246 (
            .O(N__40953),
            .I(n11989));
    InMux I__8245 (
            .O(N__40950),
            .I(N__40945));
    InMux I__8244 (
            .O(N__40949),
            .I(N__40942));
    InMux I__8243 (
            .O(N__40948),
            .I(N__40939));
    LocalMux I__8242 (
            .O(N__40945),
            .I(N__40934));
    LocalMux I__8241 (
            .O(N__40942),
            .I(N__40934));
    LocalMux I__8240 (
            .O(N__40939),
            .I(N__40931));
    Span4Mux_h I__8239 (
            .O(N__40934),
            .I(N__40928));
    Span4Mux_h I__8238 (
            .O(N__40931),
            .I(N__40925));
    Odrv4 I__8237 (
            .O(N__40928),
            .I(n304));
    Odrv4 I__8236 (
            .O(N__40925),
            .I(n304));
    InMux I__8235 (
            .O(N__40920),
            .I(N__40917));
    LocalMux I__8234 (
            .O(N__40917),
            .I(n1901));
    InMux I__8233 (
            .O(N__40914),
            .I(bfn_11_17_0_));
    InMux I__8232 (
            .O(N__40911),
            .I(N__40907));
    CascadeMux I__8231 (
            .O(N__40910),
            .I(N__40904));
    LocalMux I__8230 (
            .O(N__40907),
            .I(N__40901));
    InMux I__8229 (
            .O(N__40904),
            .I(N__40898));
    Odrv4 I__8228 (
            .O(N__40901),
            .I(n1833));
    LocalMux I__8227 (
            .O(N__40898),
            .I(n1833));
    InMux I__8226 (
            .O(N__40893),
            .I(N__40890));
    LocalMux I__8225 (
            .O(N__40890),
            .I(n1900));
    InMux I__8224 (
            .O(N__40887),
            .I(n12606));
    CascadeMux I__8223 (
            .O(N__40884),
            .I(N__40880));
    InMux I__8222 (
            .O(N__40883),
            .I(N__40876));
    InMux I__8221 (
            .O(N__40880),
            .I(N__40873));
    InMux I__8220 (
            .O(N__40879),
            .I(N__40870));
    LocalMux I__8219 (
            .O(N__40876),
            .I(n1832));
    LocalMux I__8218 (
            .O(N__40873),
            .I(n1832));
    LocalMux I__8217 (
            .O(N__40870),
            .I(n1832));
    CascadeMux I__8216 (
            .O(N__40863),
            .I(N__40860));
    InMux I__8215 (
            .O(N__40860),
            .I(N__40857));
    LocalMux I__8214 (
            .O(N__40857),
            .I(n1899));
    InMux I__8213 (
            .O(N__40854),
            .I(n12607));
    CascadeMux I__8212 (
            .O(N__40851),
            .I(N__40848));
    InMux I__8211 (
            .O(N__40848),
            .I(N__40844));
    InMux I__8210 (
            .O(N__40847),
            .I(N__40841));
    LocalMux I__8209 (
            .O(N__40844),
            .I(n1831));
    LocalMux I__8208 (
            .O(N__40841),
            .I(n1831));
    InMux I__8207 (
            .O(N__40836),
            .I(N__40833));
    LocalMux I__8206 (
            .O(N__40833),
            .I(n1898));
    InMux I__8205 (
            .O(N__40830),
            .I(N__40827));
    LocalMux I__8204 (
            .O(N__40827),
            .I(n10_adj_687));
    InMux I__8203 (
            .O(N__40824),
            .I(bfn_10_31_0_));
    InMux I__8202 (
            .O(N__40821),
            .I(N__40818));
    LocalMux I__8201 (
            .O(N__40818),
            .I(n9_adj_686));
    InMux I__8200 (
            .O(N__40815),
            .I(n13086));
    InMux I__8199 (
            .O(N__40812),
            .I(N__40809));
    LocalMux I__8198 (
            .O(N__40809),
            .I(n8_adj_685));
    InMux I__8197 (
            .O(N__40806),
            .I(n13087));
    InMux I__8196 (
            .O(N__40803),
            .I(N__40800));
    LocalMux I__8195 (
            .O(N__40800),
            .I(n7_adj_684));
    InMux I__8194 (
            .O(N__40797),
            .I(n13088));
    InMux I__8193 (
            .O(N__40794),
            .I(N__40791));
    LocalMux I__8192 (
            .O(N__40791),
            .I(n6_adj_683));
    InMux I__8191 (
            .O(N__40788),
            .I(n13089));
    CascadeMux I__8190 (
            .O(N__40785),
            .I(N__40781));
    InMux I__8189 (
            .O(N__40784),
            .I(N__40775));
    InMux I__8188 (
            .O(N__40781),
            .I(N__40775));
    InMux I__8187 (
            .O(N__40780),
            .I(N__40772));
    LocalMux I__8186 (
            .O(N__40775),
            .I(blink_counter_21));
    LocalMux I__8185 (
            .O(N__40772),
            .I(blink_counter_21));
    InMux I__8184 (
            .O(N__40767),
            .I(n13090));
    InMux I__8183 (
            .O(N__40764),
            .I(N__40757));
    InMux I__8182 (
            .O(N__40763),
            .I(N__40757));
    InMux I__8181 (
            .O(N__40762),
            .I(N__40754));
    LocalMux I__8180 (
            .O(N__40757),
            .I(blink_counter_22));
    LocalMux I__8179 (
            .O(N__40754),
            .I(blink_counter_22));
    InMux I__8178 (
            .O(N__40749),
            .I(n13091));
    CascadeMux I__8177 (
            .O(N__40746),
            .I(N__40743));
    InMux I__8176 (
            .O(N__40743),
            .I(N__40736));
    InMux I__8175 (
            .O(N__40742),
            .I(N__40736));
    InMux I__8174 (
            .O(N__40741),
            .I(N__40733));
    LocalMux I__8173 (
            .O(N__40736),
            .I(blink_counter_23));
    LocalMux I__8172 (
            .O(N__40733),
            .I(blink_counter_23));
    InMux I__8171 (
            .O(N__40728),
            .I(n13092));
    InMux I__8170 (
            .O(N__40725),
            .I(N__40722));
    LocalMux I__8169 (
            .O(N__40722),
            .I(n19_adj_696));
    InMux I__8168 (
            .O(N__40719),
            .I(n13076));
    InMux I__8167 (
            .O(N__40716),
            .I(N__40713));
    LocalMux I__8166 (
            .O(N__40713),
            .I(n18_adj_695));
    InMux I__8165 (
            .O(N__40710),
            .I(bfn_10_30_0_));
    InMux I__8164 (
            .O(N__40707),
            .I(N__40704));
    LocalMux I__8163 (
            .O(N__40704),
            .I(n17_adj_694));
    InMux I__8162 (
            .O(N__40701),
            .I(n13078));
    InMux I__8161 (
            .O(N__40698),
            .I(N__40695));
    LocalMux I__8160 (
            .O(N__40695),
            .I(n16_adj_693));
    InMux I__8159 (
            .O(N__40692),
            .I(n13079));
    InMux I__8158 (
            .O(N__40689),
            .I(N__40686));
    LocalMux I__8157 (
            .O(N__40686),
            .I(n15_adj_692));
    InMux I__8156 (
            .O(N__40683),
            .I(n13080));
    InMux I__8155 (
            .O(N__40680),
            .I(N__40677));
    LocalMux I__8154 (
            .O(N__40677),
            .I(n14_adj_691));
    InMux I__8153 (
            .O(N__40674),
            .I(n13081));
    InMux I__8152 (
            .O(N__40671),
            .I(N__40668));
    LocalMux I__8151 (
            .O(N__40668),
            .I(n13_adj_690));
    InMux I__8150 (
            .O(N__40665),
            .I(n13082));
    InMux I__8149 (
            .O(N__40662),
            .I(N__40659));
    LocalMux I__8148 (
            .O(N__40659),
            .I(n12_adj_689));
    InMux I__8147 (
            .O(N__40656),
            .I(n13083));
    InMux I__8146 (
            .O(N__40653),
            .I(N__40650));
    LocalMux I__8145 (
            .O(N__40650),
            .I(n11_adj_688));
    InMux I__8144 (
            .O(N__40647),
            .I(n13084));
    InMux I__8143 (
            .O(N__40644),
            .I(N__40641));
    LocalMux I__8142 (
            .O(N__40641),
            .I(n26_adj_703));
    InMux I__8141 (
            .O(N__40638),
            .I(bfn_10_29_0_));
    InMux I__8140 (
            .O(N__40635),
            .I(N__40632));
    LocalMux I__8139 (
            .O(N__40632),
            .I(n25_adj_702));
    InMux I__8138 (
            .O(N__40629),
            .I(n13070));
    InMux I__8137 (
            .O(N__40626),
            .I(N__40623));
    LocalMux I__8136 (
            .O(N__40623),
            .I(n24_adj_701));
    InMux I__8135 (
            .O(N__40620),
            .I(n13071));
    InMux I__8134 (
            .O(N__40617),
            .I(N__40614));
    LocalMux I__8133 (
            .O(N__40614),
            .I(n23_adj_700));
    InMux I__8132 (
            .O(N__40611),
            .I(n13072));
    InMux I__8131 (
            .O(N__40608),
            .I(N__40605));
    LocalMux I__8130 (
            .O(N__40605),
            .I(n22_adj_699));
    InMux I__8129 (
            .O(N__40602),
            .I(n13073));
    InMux I__8128 (
            .O(N__40599),
            .I(N__40596));
    LocalMux I__8127 (
            .O(N__40596),
            .I(n21_adj_698));
    InMux I__8126 (
            .O(N__40593),
            .I(n13074));
    InMux I__8125 (
            .O(N__40590),
            .I(N__40587));
    LocalMux I__8124 (
            .O(N__40587),
            .I(n20_adj_697));
    InMux I__8123 (
            .O(N__40584),
            .I(n13075));
    InMux I__8122 (
            .O(N__40581),
            .I(N__40578));
    LocalMux I__8121 (
            .O(N__40578),
            .I(N__40575));
    Odrv12 I__8120 (
            .O(N__40575),
            .I(encoder0_position_scaled_21));
    InMux I__8119 (
            .O(N__40572),
            .I(N__40569));
    LocalMux I__8118 (
            .O(N__40569),
            .I(N__40566));
    Odrv4 I__8117 (
            .O(N__40566),
            .I(encoder0_position_scaled_19));
    InMux I__8116 (
            .O(N__40563),
            .I(N__40559));
    InMux I__8115 (
            .O(N__40562),
            .I(N__40556));
    LocalMux I__8114 (
            .O(N__40559),
            .I(pwm_setpoint_4));
    LocalMux I__8113 (
            .O(N__40556),
            .I(pwm_setpoint_4));
    InMux I__8112 (
            .O(N__40551),
            .I(N__40548));
    LocalMux I__8111 (
            .O(N__40548),
            .I(N__40545));
    Odrv12 I__8110 (
            .O(N__40545),
            .I(encoder0_position_scaled_22));
    InMux I__8109 (
            .O(N__40542),
            .I(N__40538));
    InMux I__8108 (
            .O(N__40541),
            .I(N__40535));
    LocalMux I__8107 (
            .O(N__40538),
            .I(N__40532));
    LocalMux I__8106 (
            .O(N__40535),
            .I(\quad_counter0.a_prev ));
    Odrv4 I__8105 (
            .O(N__40532),
            .I(\quad_counter0.a_prev ));
    CascadeMux I__8104 (
            .O(N__40527),
            .I(N__40509));
    CascadeMux I__8103 (
            .O(N__40526),
            .I(N__40505));
    CascadeMux I__8102 (
            .O(N__40525),
            .I(N__40501));
    CascadeMux I__8101 (
            .O(N__40524),
            .I(N__40497));
    CascadeMux I__8100 (
            .O(N__40523),
            .I(N__40493));
    CascadeMux I__8099 (
            .O(N__40522),
            .I(N__40489));
    CascadeMux I__8098 (
            .O(N__40521),
            .I(N__40485));
    CascadeMux I__8097 (
            .O(N__40520),
            .I(N__40481));
    CascadeMux I__8096 (
            .O(N__40519),
            .I(N__40477));
    CascadeMux I__8095 (
            .O(N__40518),
            .I(N__40473));
    CascadeMux I__8094 (
            .O(N__40517),
            .I(N__40469));
    CascadeMux I__8093 (
            .O(N__40516),
            .I(N__40464));
    CascadeMux I__8092 (
            .O(N__40515),
            .I(N__40460));
    CascadeMux I__8091 (
            .O(N__40514),
            .I(N__40456));
    InMux I__8090 (
            .O(N__40513),
            .I(N__40438));
    InMux I__8089 (
            .O(N__40512),
            .I(N__40438));
    InMux I__8088 (
            .O(N__40509),
            .I(N__40438));
    InMux I__8087 (
            .O(N__40508),
            .I(N__40438));
    InMux I__8086 (
            .O(N__40505),
            .I(N__40438));
    InMux I__8085 (
            .O(N__40504),
            .I(N__40438));
    InMux I__8084 (
            .O(N__40501),
            .I(N__40438));
    InMux I__8083 (
            .O(N__40500),
            .I(N__40438));
    InMux I__8082 (
            .O(N__40497),
            .I(N__40421));
    InMux I__8081 (
            .O(N__40496),
            .I(N__40421));
    InMux I__8080 (
            .O(N__40493),
            .I(N__40421));
    InMux I__8079 (
            .O(N__40492),
            .I(N__40421));
    InMux I__8078 (
            .O(N__40489),
            .I(N__40421));
    InMux I__8077 (
            .O(N__40488),
            .I(N__40421));
    InMux I__8076 (
            .O(N__40485),
            .I(N__40421));
    InMux I__8075 (
            .O(N__40484),
            .I(N__40421));
    InMux I__8074 (
            .O(N__40481),
            .I(N__40404));
    InMux I__8073 (
            .O(N__40480),
            .I(N__40404));
    InMux I__8072 (
            .O(N__40477),
            .I(N__40404));
    InMux I__8071 (
            .O(N__40476),
            .I(N__40404));
    InMux I__8070 (
            .O(N__40473),
            .I(N__40404));
    InMux I__8069 (
            .O(N__40472),
            .I(N__40404));
    InMux I__8068 (
            .O(N__40469),
            .I(N__40404));
    InMux I__8067 (
            .O(N__40468),
            .I(N__40404));
    InMux I__8066 (
            .O(N__40467),
            .I(N__40389));
    InMux I__8065 (
            .O(N__40464),
            .I(N__40389));
    InMux I__8064 (
            .O(N__40463),
            .I(N__40389));
    InMux I__8063 (
            .O(N__40460),
            .I(N__40389));
    InMux I__8062 (
            .O(N__40459),
            .I(N__40389));
    InMux I__8061 (
            .O(N__40456),
            .I(N__40389));
    InMux I__8060 (
            .O(N__40455),
            .I(N__40389));
    LocalMux I__8059 (
            .O(N__40438),
            .I(N__40386));
    LocalMux I__8058 (
            .O(N__40421),
            .I(N__40379));
    LocalMux I__8057 (
            .O(N__40404),
            .I(N__40379));
    LocalMux I__8056 (
            .O(N__40389),
            .I(N__40379));
    Sp12to4 I__8055 (
            .O(N__40386),
            .I(N__40374));
    Span12Mux_v I__8054 (
            .O(N__40379),
            .I(N__40374));
    Odrv12 I__8053 (
            .O(N__40374),
            .I(\quad_counter0.direction_N_536 ));
    InMux I__8052 (
            .O(N__40371),
            .I(N__40368));
    LocalMux I__8051 (
            .O(N__40368),
            .I(N__40365));
    Odrv4 I__8050 (
            .O(N__40365),
            .I(encoder0_position_scaled_1));
    InMux I__8049 (
            .O(N__40362),
            .I(N__40359));
    LocalMux I__8048 (
            .O(N__40359),
            .I(\quad_counter0.direction_N_540 ));
    InMux I__8047 (
            .O(N__40356),
            .I(N__40353));
    LocalMux I__8046 (
            .O(N__40353),
            .I(N__40350));
    Odrv4 I__8045 (
            .O(N__40350),
            .I(encoder0_position_scaled_9));
    InMux I__8044 (
            .O(N__40347),
            .I(N__40344));
    LocalMux I__8043 (
            .O(N__40344),
            .I(N__40341));
    Span4Mux_h I__8042 (
            .O(N__40341),
            .I(N__40338));
    Odrv4 I__8041 (
            .O(N__40338),
            .I(encoder0_position_scaled_20));
    InMux I__8040 (
            .O(N__40335),
            .I(N__40332));
    LocalMux I__8039 (
            .O(N__40332),
            .I(N__40329));
    Odrv12 I__8038 (
            .O(N__40329),
            .I(encoder0_position_scaled_11));
    CascadeMux I__8037 (
            .O(N__40326),
            .I(N__40323));
    InMux I__8036 (
            .O(N__40323),
            .I(N__40320));
    LocalMux I__8035 (
            .O(N__40320),
            .I(n15_adj_633));
    CascadeMux I__8034 (
            .O(N__40317),
            .I(N__40314));
    InMux I__8033 (
            .O(N__40314),
            .I(N__40311));
    LocalMux I__8032 (
            .O(N__40311),
            .I(n6_adj_624));
    CEMux I__8031 (
            .O(N__40308),
            .I(N__40305));
    LocalMux I__8030 (
            .O(N__40305),
            .I(N__40299));
    CEMux I__8029 (
            .O(N__40304),
            .I(N__40296));
    CEMux I__8028 (
            .O(N__40303),
            .I(N__40293));
    CEMux I__8027 (
            .O(N__40302),
            .I(N__40290));
    Span4Mux_v I__8026 (
            .O(N__40299),
            .I(N__40287));
    LocalMux I__8025 (
            .O(N__40296),
            .I(N__40284));
    LocalMux I__8024 (
            .O(N__40293),
            .I(N__40281));
    LocalMux I__8023 (
            .O(N__40290),
            .I(N__40278));
    Span4Mux_v I__8022 (
            .O(N__40287),
            .I(N__40275));
    Span12Mux_v I__8021 (
            .O(N__40284),
            .I(N__40272));
    Span4Mux_v I__8020 (
            .O(N__40281),
            .I(N__40267));
    Span4Mux_h I__8019 (
            .O(N__40278),
            .I(N__40267));
    Odrv4 I__8018 (
            .O(N__40275),
            .I(direction_N_537));
    Odrv12 I__8017 (
            .O(N__40272),
            .I(direction_N_537));
    Odrv4 I__8016 (
            .O(N__40267),
            .I(direction_N_537));
    CascadeMux I__8015 (
            .O(N__40260),
            .I(direction_N_537_cascade_));
    InMux I__8014 (
            .O(N__40257),
            .I(N__40254));
    LocalMux I__8013 (
            .O(N__40254),
            .I(n1302));
    CascadeMux I__8012 (
            .O(N__40251),
            .I(N__40248));
    InMux I__8011 (
            .O(N__40248),
            .I(N__40245));
    LocalMux I__8010 (
            .O(N__40245),
            .I(n8_adj_626));
    CascadeMux I__8009 (
            .O(N__40242),
            .I(N__40239));
    InMux I__8008 (
            .O(N__40239),
            .I(N__40236));
    LocalMux I__8007 (
            .O(N__40236),
            .I(n5_adj_623));
    CascadeMux I__8006 (
            .O(N__40233),
            .I(N__40217));
    CascadeMux I__8005 (
            .O(N__40232),
            .I(N__40214));
    CascadeMux I__8004 (
            .O(N__40231),
            .I(N__40211));
    CascadeMux I__8003 (
            .O(N__40230),
            .I(N__40207));
    CascadeMux I__8002 (
            .O(N__40229),
            .I(N__40203));
    CascadeMux I__8001 (
            .O(N__40228),
            .I(N__40200));
    CascadeMux I__8000 (
            .O(N__40227),
            .I(N__40197));
    CascadeMux I__7999 (
            .O(N__40226),
            .I(N__40194));
    CascadeMux I__7998 (
            .O(N__40225),
            .I(N__40191));
    CascadeMux I__7997 (
            .O(N__40224),
            .I(N__40188));
    CascadeMux I__7996 (
            .O(N__40223),
            .I(N__40185));
    CascadeMux I__7995 (
            .O(N__40222),
            .I(N__40182));
    CascadeMux I__7994 (
            .O(N__40221),
            .I(N__40179));
    CascadeMux I__7993 (
            .O(N__40220),
            .I(N__40176));
    InMux I__7992 (
            .O(N__40217),
            .I(N__40164));
    InMux I__7991 (
            .O(N__40214),
            .I(N__40164));
    InMux I__7990 (
            .O(N__40211),
            .I(N__40151));
    InMux I__7989 (
            .O(N__40210),
            .I(N__40151));
    InMux I__7988 (
            .O(N__40207),
            .I(N__40151));
    InMux I__7987 (
            .O(N__40206),
            .I(N__40151));
    InMux I__7986 (
            .O(N__40203),
            .I(N__40151));
    InMux I__7985 (
            .O(N__40200),
            .I(N__40151));
    InMux I__7984 (
            .O(N__40197),
            .I(N__40142));
    InMux I__7983 (
            .O(N__40194),
            .I(N__40142));
    InMux I__7982 (
            .O(N__40191),
            .I(N__40142));
    InMux I__7981 (
            .O(N__40188),
            .I(N__40142));
    InMux I__7980 (
            .O(N__40185),
            .I(N__40133));
    InMux I__7979 (
            .O(N__40182),
            .I(N__40133));
    InMux I__7978 (
            .O(N__40179),
            .I(N__40133));
    InMux I__7977 (
            .O(N__40176),
            .I(N__40133));
    CascadeMux I__7976 (
            .O(N__40175),
            .I(N__40130));
    CascadeMux I__7975 (
            .O(N__40174),
            .I(N__40127));
    CascadeMux I__7974 (
            .O(N__40173),
            .I(N__40124));
    CascadeMux I__7973 (
            .O(N__40172),
            .I(N__40121));
    CascadeMux I__7972 (
            .O(N__40171),
            .I(N__40118));
    CascadeMux I__7971 (
            .O(N__40170),
            .I(N__40115));
    CascadeMux I__7970 (
            .O(N__40169),
            .I(N__40112));
    LocalMux I__7969 (
            .O(N__40164),
            .I(N__40102));
    LocalMux I__7968 (
            .O(N__40151),
            .I(N__40102));
    LocalMux I__7967 (
            .O(N__40142),
            .I(N__40102));
    LocalMux I__7966 (
            .O(N__40133),
            .I(N__40102));
    InMux I__7965 (
            .O(N__40130),
            .I(N__40095));
    InMux I__7964 (
            .O(N__40127),
            .I(N__40095));
    InMux I__7963 (
            .O(N__40124),
            .I(N__40095));
    InMux I__7962 (
            .O(N__40121),
            .I(N__40084));
    InMux I__7961 (
            .O(N__40118),
            .I(N__40084));
    InMux I__7960 (
            .O(N__40115),
            .I(N__40084));
    InMux I__7959 (
            .O(N__40112),
            .I(N__40084));
    InMux I__7958 (
            .O(N__40111),
            .I(N__40084));
    Span4Mux_v I__7957 (
            .O(N__40102),
            .I(N__40080));
    LocalMux I__7956 (
            .O(N__40095),
            .I(N__40075));
    LocalMux I__7955 (
            .O(N__40084),
            .I(N__40075));
    InMux I__7954 (
            .O(N__40083),
            .I(N__40072));
    Odrv4 I__7953 (
            .O(N__40080),
            .I(n2_adj_620));
    Odrv12 I__7952 (
            .O(N__40075),
            .I(n2_adj_620));
    LocalMux I__7951 (
            .O(N__40072),
            .I(n2_adj_620));
    CascadeMux I__7950 (
            .O(N__40065),
            .I(N__40062));
    InMux I__7949 (
            .O(N__40062),
            .I(N__40059));
    LocalMux I__7948 (
            .O(N__40059),
            .I(n9_adj_627));
    InMux I__7947 (
            .O(N__40056),
            .I(N__40053));
    LocalMux I__7946 (
            .O(N__40053),
            .I(N__40050));
    Odrv4 I__7945 (
            .O(N__40050),
            .I(encoder0_position_scaled_5));
    CascadeMux I__7944 (
            .O(N__40047),
            .I(N__40044));
    InMux I__7943 (
            .O(N__40044),
            .I(N__40041));
    LocalMux I__7942 (
            .O(N__40041),
            .I(n38));
    CascadeMux I__7941 (
            .O(N__40038),
            .I(N__40035));
    InMux I__7940 (
            .O(N__40035),
            .I(N__40032));
    LocalMux I__7939 (
            .O(N__40032),
            .I(n402));
    CascadeMux I__7938 (
            .O(N__40029),
            .I(N__40026));
    InMux I__7937 (
            .O(N__40026),
            .I(N__40023));
    LocalMux I__7936 (
            .O(N__40023),
            .I(n39));
    InMux I__7935 (
            .O(N__40020),
            .I(N__40017));
    LocalMux I__7934 (
            .O(N__40017),
            .I(n2562));
    CEMux I__7933 (
            .O(N__40014),
            .I(N__40011));
    LocalMux I__7932 (
            .O(N__40011),
            .I(N__40008));
    Span4Mux_h I__7931 (
            .O(N__40008),
            .I(N__40005));
    Odrv4 I__7930 (
            .O(N__40005),
            .I(n5187));
    InMux I__7929 (
            .O(N__40002),
            .I(N__39997));
    InMux I__7928 (
            .O(N__40001),
            .I(N__39994));
    InMux I__7927 (
            .O(N__40000),
            .I(N__39991));
    LocalMux I__7926 (
            .O(N__39997),
            .I(N__39988));
    LocalMux I__7925 (
            .O(N__39994),
            .I(encoder0_position_11));
    LocalMux I__7924 (
            .O(N__39991),
            .I(encoder0_position_11));
    Odrv12 I__7923 (
            .O(N__39988),
            .I(encoder0_position_11));
    CascadeMux I__7922 (
            .O(N__39981),
            .I(N__39978));
    InMux I__7921 (
            .O(N__39978),
            .I(N__39975));
    LocalMux I__7920 (
            .O(N__39975),
            .I(n22_adj_640));
    InMux I__7919 (
            .O(N__39972),
            .I(N__39967));
    InMux I__7918 (
            .O(N__39971),
            .I(N__39964));
    CascadeMux I__7917 (
            .O(N__39970),
            .I(N__39961));
    LocalMux I__7916 (
            .O(N__39967),
            .I(N__39958));
    LocalMux I__7915 (
            .O(N__39964),
            .I(N__39955));
    InMux I__7914 (
            .O(N__39961),
            .I(N__39952));
    Span4Mux_h I__7913 (
            .O(N__39958),
            .I(N__39949));
    Span4Mux_v I__7912 (
            .O(N__39955),
            .I(N__39946));
    LocalMux I__7911 (
            .O(N__39952),
            .I(encoder0_position_12));
    Odrv4 I__7910 (
            .O(N__39949),
            .I(encoder0_position_12));
    Odrv4 I__7909 (
            .O(N__39946),
            .I(encoder0_position_12));
    CascadeMux I__7908 (
            .O(N__39939),
            .I(N__39936));
    InMux I__7907 (
            .O(N__39936),
            .I(N__39933));
    LocalMux I__7906 (
            .O(N__39933),
            .I(n21_adj_639));
    InMux I__7905 (
            .O(N__39930),
            .I(N__39925));
    InMux I__7904 (
            .O(N__39929),
            .I(N__39922));
    InMux I__7903 (
            .O(N__39928),
            .I(N__39919));
    LocalMux I__7902 (
            .O(N__39925),
            .I(N__39916));
    LocalMux I__7901 (
            .O(N__39922),
            .I(encoder0_position_13));
    LocalMux I__7900 (
            .O(N__39919),
            .I(encoder0_position_13));
    Odrv12 I__7899 (
            .O(N__39916),
            .I(encoder0_position_13));
    CascadeMux I__7898 (
            .O(N__39909),
            .I(N__39906));
    InMux I__7897 (
            .O(N__39906),
            .I(N__39903));
    LocalMux I__7896 (
            .O(N__39903),
            .I(n20_adj_638));
    InMux I__7895 (
            .O(N__39900),
            .I(n12496));
    InMux I__7894 (
            .O(N__39897),
            .I(n12497));
    InMux I__7893 (
            .O(N__39894),
            .I(n12498));
    InMux I__7892 (
            .O(N__39891),
            .I(n12499));
    InMux I__7891 (
            .O(N__39888),
            .I(n12500));
    InMux I__7890 (
            .O(N__39885),
            .I(N__39882));
    LocalMux I__7889 (
            .O(N__39882),
            .I(n2563));
    InMux I__7888 (
            .O(N__39879),
            .I(N__39876));
    LocalMux I__7887 (
            .O(N__39876),
            .I(n13656));
    CascadeMux I__7886 (
            .O(N__39873),
            .I(N__39870));
    InMux I__7885 (
            .O(N__39870),
            .I(N__39867));
    LocalMux I__7884 (
            .O(N__39867),
            .I(n403));
    CascadeMux I__7883 (
            .O(N__39864),
            .I(N__39861));
    InMux I__7882 (
            .O(N__39861),
            .I(N__39858));
    LocalMux I__7881 (
            .O(N__39858),
            .I(n13_adj_631));
    InMux I__7880 (
            .O(N__39855),
            .I(bfn_10_21_0_));
    InMux I__7879 (
            .O(N__39852),
            .I(\quad_counter0.n13119 ));
    InMux I__7878 (
            .O(N__39849),
            .I(\quad_counter0.n13120 ));
    InMux I__7877 (
            .O(N__39846),
            .I(\quad_counter0.n13121 ));
    InMux I__7876 (
            .O(N__39843),
            .I(\quad_counter0.n13122 ));
    InMux I__7875 (
            .O(N__39840),
            .I(\quad_counter0.n13123 ));
    InMux I__7874 (
            .O(N__39837),
            .I(\quad_counter0.n13124 ));
    InMux I__7873 (
            .O(N__39834),
            .I(\quad_counter0.n13125 ));
    InMux I__7872 (
            .O(N__39831),
            .I(bfn_10_22_0_));
    InMux I__7871 (
            .O(N__39828),
            .I(N__39823));
    InMux I__7870 (
            .O(N__39827),
            .I(N__39818));
    InMux I__7869 (
            .O(N__39826),
            .I(N__39818));
    LocalMux I__7868 (
            .O(N__39823),
            .I(encoder0_position_15));
    LocalMux I__7867 (
            .O(N__39818),
            .I(encoder0_position_15));
    InMux I__7866 (
            .O(N__39813),
            .I(\quad_counter0.n13109 ));
    InMux I__7865 (
            .O(N__39810),
            .I(bfn_10_20_0_));
    InMux I__7864 (
            .O(N__39807),
            .I(\quad_counter0.n13111 ));
    InMux I__7863 (
            .O(N__39804),
            .I(\quad_counter0.n13112 ));
    CascadeMux I__7862 (
            .O(N__39801),
            .I(N__39796));
    InMux I__7861 (
            .O(N__39800),
            .I(N__39793));
    InMux I__7860 (
            .O(N__39799),
            .I(N__39790));
    InMux I__7859 (
            .O(N__39796),
            .I(N__39787));
    LocalMux I__7858 (
            .O(N__39793),
            .I(encoder0_position_19));
    LocalMux I__7857 (
            .O(N__39790),
            .I(encoder0_position_19));
    LocalMux I__7856 (
            .O(N__39787),
            .I(encoder0_position_19));
    InMux I__7855 (
            .O(N__39780),
            .I(\quad_counter0.n13113 ));
    InMux I__7854 (
            .O(N__39777),
            .I(\quad_counter0.n13114 ));
    InMux I__7853 (
            .O(N__39774),
            .I(\quad_counter0.n13115 ));
    InMux I__7852 (
            .O(N__39771),
            .I(\quad_counter0.n13116 ));
    InMux I__7851 (
            .O(N__39768),
            .I(\quad_counter0.n13117 ));
    InMux I__7850 (
            .O(N__39765),
            .I(N__39761));
    CascadeMux I__7849 (
            .O(N__39764),
            .I(N__39757));
    LocalMux I__7848 (
            .O(N__39761),
            .I(N__39754));
    InMux I__7847 (
            .O(N__39760),
            .I(N__39751));
    InMux I__7846 (
            .O(N__39757),
            .I(N__39748));
    Span4Mux_h I__7845 (
            .O(N__39754),
            .I(N__39743));
    LocalMux I__7844 (
            .O(N__39751),
            .I(N__39743));
    LocalMux I__7843 (
            .O(N__39748),
            .I(encoder0_position_7));
    Odrv4 I__7842 (
            .O(N__39743),
            .I(encoder0_position_7));
    InMux I__7841 (
            .O(N__39738),
            .I(\quad_counter0.n13101 ));
    InMux I__7840 (
            .O(N__39735),
            .I(N__39732));
    LocalMux I__7839 (
            .O(N__39732),
            .I(N__39728));
    CascadeMux I__7838 (
            .O(N__39731),
            .I(N__39724));
    Span4Mux_h I__7837 (
            .O(N__39728),
            .I(N__39721));
    CascadeMux I__7836 (
            .O(N__39727),
            .I(N__39718));
    InMux I__7835 (
            .O(N__39724),
            .I(N__39715));
    Span4Mux_v I__7834 (
            .O(N__39721),
            .I(N__39712));
    InMux I__7833 (
            .O(N__39718),
            .I(N__39709));
    LocalMux I__7832 (
            .O(N__39715),
            .I(encoder0_position_8));
    Odrv4 I__7831 (
            .O(N__39712),
            .I(encoder0_position_8));
    LocalMux I__7830 (
            .O(N__39709),
            .I(encoder0_position_8));
    InMux I__7829 (
            .O(N__39702),
            .I(bfn_10_19_0_));
    InMux I__7828 (
            .O(N__39699),
            .I(N__39696));
    LocalMux I__7827 (
            .O(N__39696),
            .I(N__39692));
    InMux I__7826 (
            .O(N__39695),
            .I(N__39688));
    Span4Mux_h I__7825 (
            .O(N__39692),
            .I(N__39685));
    InMux I__7824 (
            .O(N__39691),
            .I(N__39682));
    LocalMux I__7823 (
            .O(N__39688),
            .I(encoder0_position_9));
    Odrv4 I__7822 (
            .O(N__39685),
            .I(encoder0_position_9));
    LocalMux I__7821 (
            .O(N__39682),
            .I(encoder0_position_9));
    InMux I__7820 (
            .O(N__39675),
            .I(\quad_counter0.n13103 ));
    CascadeMux I__7819 (
            .O(N__39672),
            .I(N__39668));
    InMux I__7818 (
            .O(N__39671),
            .I(N__39665));
    InMux I__7817 (
            .O(N__39668),
            .I(N__39661));
    LocalMux I__7816 (
            .O(N__39665),
            .I(N__39658));
    InMux I__7815 (
            .O(N__39664),
            .I(N__39655));
    LocalMux I__7814 (
            .O(N__39661),
            .I(encoder0_position_10));
    Odrv4 I__7813 (
            .O(N__39658),
            .I(encoder0_position_10));
    LocalMux I__7812 (
            .O(N__39655),
            .I(encoder0_position_10));
    InMux I__7811 (
            .O(N__39648),
            .I(\quad_counter0.n13104 ));
    InMux I__7810 (
            .O(N__39645),
            .I(\quad_counter0.n13105 ));
    InMux I__7809 (
            .O(N__39642),
            .I(\quad_counter0.n13106 ));
    InMux I__7808 (
            .O(N__39639),
            .I(\quad_counter0.n13107 ));
    CascadeMux I__7807 (
            .O(N__39636),
            .I(N__39633));
    InMux I__7806 (
            .O(N__39633),
            .I(N__39628));
    InMux I__7805 (
            .O(N__39632),
            .I(N__39625));
    InMux I__7804 (
            .O(N__39631),
            .I(N__39622));
    LocalMux I__7803 (
            .O(N__39628),
            .I(encoder0_position_14));
    LocalMux I__7802 (
            .O(N__39625),
            .I(encoder0_position_14));
    LocalMux I__7801 (
            .O(N__39622),
            .I(encoder0_position_14));
    InMux I__7800 (
            .O(N__39615),
            .I(\quad_counter0.n13108 ));
    InMux I__7799 (
            .O(N__39612),
            .I(N__39609));
    LocalMux I__7798 (
            .O(N__39609),
            .I(N__39605));
    CascadeMux I__7797 (
            .O(N__39608),
            .I(N__39602));
    Span4Mux_h I__7796 (
            .O(N__39605),
            .I(N__39598));
    InMux I__7795 (
            .O(N__39602),
            .I(N__39595));
    InMux I__7794 (
            .O(N__39601),
            .I(N__39592));
    Odrv4 I__7793 (
            .O(N__39598),
            .I(n1925));
    LocalMux I__7792 (
            .O(N__39595),
            .I(n1925));
    LocalMux I__7791 (
            .O(N__39592),
            .I(n1925));
    CascadeMux I__7790 (
            .O(N__39585),
            .I(n1928_cascade_));
    InMux I__7789 (
            .O(N__39582),
            .I(N__39579));
    LocalMux I__7788 (
            .O(N__39579),
            .I(N__39575));
    CascadeMux I__7787 (
            .O(N__39578),
            .I(N__39572));
    Span4Mux_h I__7786 (
            .O(N__39575),
            .I(N__39568));
    InMux I__7785 (
            .O(N__39572),
            .I(N__39565));
    InMux I__7784 (
            .O(N__39571),
            .I(N__39562));
    Odrv4 I__7783 (
            .O(N__39568),
            .I(n1923));
    LocalMux I__7782 (
            .O(N__39565),
            .I(n1923));
    LocalMux I__7781 (
            .O(N__39562),
            .I(n1923));
    CascadeMux I__7780 (
            .O(N__39555),
            .I(N__39552));
    InMux I__7779 (
            .O(N__39552),
            .I(N__39549));
    LocalMux I__7778 (
            .O(N__39549),
            .I(N__39546));
    Span4Mux_h I__7777 (
            .O(N__39546),
            .I(N__39543));
    Odrv4 I__7776 (
            .O(N__39543),
            .I(n14440));
    InMux I__7775 (
            .O(N__39540),
            .I(N__39537));
    LocalMux I__7774 (
            .O(N__39537),
            .I(N__39532));
    InMux I__7773 (
            .O(N__39536),
            .I(N__39529));
    CascadeMux I__7772 (
            .O(N__39535),
            .I(N__39526));
    Span4Mux_v I__7771 (
            .O(N__39532),
            .I(N__39521));
    LocalMux I__7770 (
            .O(N__39529),
            .I(N__39521));
    InMux I__7769 (
            .O(N__39526),
            .I(N__39518));
    Odrv4 I__7768 (
            .O(N__39521),
            .I(n1932));
    LocalMux I__7767 (
            .O(N__39518),
            .I(n1932));
    InMux I__7766 (
            .O(N__39513),
            .I(N__39510));
    LocalMux I__7765 (
            .O(N__39510),
            .I(N__39507));
    Span4Mux_h I__7764 (
            .O(N__39507),
            .I(N__39502));
    CascadeMux I__7763 (
            .O(N__39506),
            .I(N__39499));
    InMux I__7762 (
            .O(N__39505),
            .I(N__39496));
    Span4Mux_v I__7761 (
            .O(N__39502),
            .I(N__39493));
    InMux I__7760 (
            .O(N__39499),
            .I(N__39490));
    LocalMux I__7759 (
            .O(N__39496),
            .I(encoder0_position_0));
    Odrv4 I__7758 (
            .O(N__39493),
            .I(encoder0_position_0));
    LocalMux I__7757 (
            .O(N__39490),
            .I(encoder0_position_0));
    InMux I__7756 (
            .O(N__39483),
            .I(bfn_10_18_0_));
    InMux I__7755 (
            .O(N__39480),
            .I(\quad_counter0.n13095 ));
    InMux I__7754 (
            .O(N__39477),
            .I(N__39474));
    LocalMux I__7753 (
            .O(N__39474),
            .I(N__39470));
    InMux I__7752 (
            .O(N__39473),
            .I(N__39466));
    Span4Mux_v I__7751 (
            .O(N__39470),
            .I(N__39463));
    InMux I__7750 (
            .O(N__39469),
            .I(N__39460));
    LocalMux I__7749 (
            .O(N__39466),
            .I(encoder0_position_2));
    Odrv4 I__7748 (
            .O(N__39463),
            .I(encoder0_position_2));
    LocalMux I__7747 (
            .O(N__39460),
            .I(encoder0_position_2));
    InMux I__7746 (
            .O(N__39453),
            .I(\quad_counter0.n13096 ));
    InMux I__7745 (
            .O(N__39450),
            .I(\quad_counter0.n13097 ));
    InMux I__7744 (
            .O(N__39447),
            .I(N__39444));
    LocalMux I__7743 (
            .O(N__39444),
            .I(N__39441));
    Span4Mux_h I__7742 (
            .O(N__39441),
            .I(N__39436));
    InMux I__7741 (
            .O(N__39440),
            .I(N__39433));
    InMux I__7740 (
            .O(N__39439),
            .I(N__39430));
    Span4Mux_v I__7739 (
            .O(N__39436),
            .I(N__39427));
    LocalMux I__7738 (
            .O(N__39433),
            .I(N__39424));
    LocalMux I__7737 (
            .O(N__39430),
            .I(encoder0_position_4));
    Odrv4 I__7736 (
            .O(N__39427),
            .I(encoder0_position_4));
    Odrv4 I__7735 (
            .O(N__39424),
            .I(encoder0_position_4));
    InMux I__7734 (
            .O(N__39417),
            .I(\quad_counter0.n13098 ));
    InMux I__7733 (
            .O(N__39414),
            .I(N__39410));
    CascadeMux I__7732 (
            .O(N__39413),
            .I(N__39407));
    LocalMux I__7731 (
            .O(N__39410),
            .I(N__39404));
    InMux I__7730 (
            .O(N__39407),
            .I(N__39400));
    Span4Mux_v I__7729 (
            .O(N__39404),
            .I(N__39397));
    InMux I__7728 (
            .O(N__39403),
            .I(N__39394));
    LocalMux I__7727 (
            .O(N__39400),
            .I(encoder0_position_5));
    Odrv4 I__7726 (
            .O(N__39397),
            .I(encoder0_position_5));
    LocalMux I__7725 (
            .O(N__39394),
            .I(encoder0_position_5));
    InMux I__7724 (
            .O(N__39387),
            .I(\quad_counter0.n13099 ));
    InMux I__7723 (
            .O(N__39384),
            .I(N__39381));
    LocalMux I__7722 (
            .O(N__39381),
            .I(N__39376));
    InMux I__7721 (
            .O(N__39380),
            .I(N__39373));
    InMux I__7720 (
            .O(N__39379),
            .I(N__39370));
    Span4Mux_v I__7719 (
            .O(N__39376),
            .I(N__39367));
    LocalMux I__7718 (
            .O(N__39373),
            .I(N__39364));
    LocalMux I__7717 (
            .O(N__39370),
            .I(encoder0_position_6));
    Odrv4 I__7716 (
            .O(N__39367),
            .I(encoder0_position_6));
    Odrv4 I__7715 (
            .O(N__39364),
            .I(encoder0_position_6));
    InMux I__7714 (
            .O(N__39357),
            .I(\quad_counter0.n13100 ));
    CascadeMux I__7713 (
            .O(N__39354),
            .I(N__39350));
    InMux I__7712 (
            .O(N__39353),
            .I(N__39346));
    InMux I__7711 (
            .O(N__39350),
            .I(N__39343));
    CascadeMux I__7710 (
            .O(N__39349),
            .I(N__39340));
    LocalMux I__7709 (
            .O(N__39346),
            .I(N__39337));
    LocalMux I__7708 (
            .O(N__39343),
            .I(N__39334));
    InMux I__7707 (
            .O(N__39340),
            .I(N__39331));
    Span4Mux_v I__7706 (
            .O(N__39337),
            .I(N__39328));
    Odrv4 I__7705 (
            .O(N__39334),
            .I(n1931));
    LocalMux I__7704 (
            .O(N__39331),
            .I(n1931));
    Odrv4 I__7703 (
            .O(N__39328),
            .I(n1931));
    CascadeMux I__7702 (
            .O(N__39321),
            .I(N__39317));
    InMux I__7701 (
            .O(N__39320),
            .I(N__39314));
    InMux I__7700 (
            .O(N__39317),
            .I(N__39310));
    LocalMux I__7699 (
            .O(N__39314),
            .I(N__39307));
    CascadeMux I__7698 (
            .O(N__39313),
            .I(N__39304));
    LocalMux I__7697 (
            .O(N__39310),
            .I(N__39301));
    Span4Mux_h I__7696 (
            .O(N__39307),
            .I(N__39298));
    InMux I__7695 (
            .O(N__39304),
            .I(N__39295));
    Span4Mux_h I__7694 (
            .O(N__39301),
            .I(N__39292));
    Odrv4 I__7693 (
            .O(N__39298),
            .I(n1933));
    LocalMux I__7692 (
            .O(N__39295),
            .I(n1933));
    Odrv4 I__7691 (
            .O(N__39292),
            .I(n1933));
    InMux I__7690 (
            .O(N__39285),
            .I(N__39282));
    LocalMux I__7689 (
            .O(N__39282),
            .I(N__39277));
    CascadeMux I__7688 (
            .O(N__39281),
            .I(N__39274));
    InMux I__7687 (
            .O(N__39280),
            .I(N__39271));
    Span4Mux_h I__7686 (
            .O(N__39277),
            .I(N__39268));
    InMux I__7685 (
            .O(N__39274),
            .I(N__39265));
    LocalMux I__7684 (
            .O(N__39271),
            .I(N__39262));
    Odrv4 I__7683 (
            .O(N__39268),
            .I(n1929));
    LocalMux I__7682 (
            .O(N__39265),
            .I(n1929));
    Odrv4 I__7681 (
            .O(N__39262),
            .I(n1929));
    CascadeMux I__7680 (
            .O(N__39255),
            .I(n14524_cascade_));
    CascadeMux I__7679 (
            .O(N__39252),
            .I(n14526_cascade_));
    CascadeMux I__7678 (
            .O(N__39249),
            .I(n1851_cascade_));
    InMux I__7677 (
            .O(N__39246),
            .I(N__39243));
    LocalMux I__7676 (
            .O(N__39243),
            .I(N__39239));
    CascadeMux I__7675 (
            .O(N__39242),
            .I(N__39236));
    Span4Mux_v I__7674 (
            .O(N__39239),
            .I(N__39233));
    InMux I__7673 (
            .O(N__39236),
            .I(N__39230));
    Odrv4 I__7672 (
            .O(N__39233),
            .I(n1928));
    LocalMux I__7671 (
            .O(N__39230),
            .I(n1928));
    CascadeMux I__7670 (
            .O(N__39225),
            .I(N__39221));
    CascadeMux I__7669 (
            .O(N__39224),
            .I(N__39218));
    InMux I__7668 (
            .O(N__39221),
            .I(N__39215));
    InMux I__7667 (
            .O(N__39218),
            .I(N__39211));
    LocalMux I__7666 (
            .O(N__39215),
            .I(N__39208));
    InMux I__7665 (
            .O(N__39214),
            .I(N__39205));
    LocalMux I__7664 (
            .O(N__39211),
            .I(dti_counter_1));
    Odrv4 I__7663 (
            .O(N__39208),
            .I(dti_counter_1));
    LocalMux I__7662 (
            .O(N__39205),
            .I(dti_counter_1));
    InMux I__7661 (
            .O(N__39198),
            .I(N__39195));
    LocalMux I__7660 (
            .O(N__39195),
            .I(N__39192));
    Odrv4 I__7659 (
            .O(N__39192),
            .I(n15076));
    InMux I__7658 (
            .O(N__39189),
            .I(N__39176));
    InMux I__7657 (
            .O(N__39188),
            .I(N__39176));
    InMux I__7656 (
            .O(N__39187),
            .I(N__39165));
    InMux I__7655 (
            .O(N__39186),
            .I(N__39165));
    InMux I__7654 (
            .O(N__39185),
            .I(N__39165));
    InMux I__7653 (
            .O(N__39184),
            .I(N__39165));
    InMux I__7652 (
            .O(N__39183),
            .I(N__39165));
    InMux I__7651 (
            .O(N__39182),
            .I(N__39160));
    InMux I__7650 (
            .O(N__39181),
            .I(N__39160));
    LocalMux I__7649 (
            .O(N__39176),
            .I(N__39157));
    LocalMux I__7648 (
            .O(N__39165),
            .I(commutation_state_prev_0));
    LocalMux I__7647 (
            .O(N__39160),
            .I(commutation_state_prev_0));
    Odrv12 I__7646 (
            .O(N__39157),
            .I(commutation_state_prev_0));
    InMux I__7645 (
            .O(N__39150),
            .I(N__39147));
    LocalMux I__7644 (
            .O(N__39147),
            .I(n14929));
    InMux I__7643 (
            .O(N__39144),
            .I(N__39141));
    LocalMux I__7642 (
            .O(N__39141),
            .I(n14928));
    IoInMux I__7641 (
            .O(N__39138),
            .I(N__39135));
    LocalMux I__7640 (
            .O(N__39135),
            .I(N__39132));
    IoSpan4Mux I__7639 (
            .O(N__39132),
            .I(N__39129));
    Odrv4 I__7638 (
            .O(N__39129),
            .I(LED_c));
    CascadeMux I__7637 (
            .O(N__39126),
            .I(n1831_cascade_));
    InMux I__7636 (
            .O(N__39123),
            .I(N__39119));
    CascadeMux I__7635 (
            .O(N__39122),
            .I(N__39115));
    LocalMux I__7634 (
            .O(N__39119),
            .I(N__39112));
    CascadeMux I__7633 (
            .O(N__39118),
            .I(N__39109));
    InMux I__7632 (
            .O(N__39115),
            .I(N__39106));
    Span4Mux_h I__7631 (
            .O(N__39112),
            .I(N__39103));
    InMux I__7630 (
            .O(N__39109),
            .I(N__39100));
    LocalMux I__7629 (
            .O(N__39106),
            .I(N__39097));
    Odrv4 I__7628 (
            .O(N__39103),
            .I(n1930));
    LocalMux I__7627 (
            .O(N__39100),
            .I(n1930));
    Odrv4 I__7626 (
            .O(N__39097),
            .I(n1930));
    InMux I__7625 (
            .O(N__39090),
            .I(N__39087));
    LocalMux I__7624 (
            .O(N__39087),
            .I(n15075));
    InMux I__7623 (
            .O(N__39084),
            .I(N__39081));
    LocalMux I__7622 (
            .O(N__39081),
            .I(n15071));
    CascadeMux I__7621 (
            .O(N__39078),
            .I(N__39074));
    CascadeMux I__7620 (
            .O(N__39077),
            .I(N__39071));
    InMux I__7619 (
            .O(N__39074),
            .I(N__39067));
    InMux I__7618 (
            .O(N__39071),
            .I(N__39064));
    InMux I__7617 (
            .O(N__39070),
            .I(N__39061));
    LocalMux I__7616 (
            .O(N__39067),
            .I(dti_counter_5));
    LocalMux I__7615 (
            .O(N__39064),
            .I(dti_counter_5));
    LocalMux I__7614 (
            .O(N__39061),
            .I(dti_counter_5));
    CascadeMux I__7613 (
            .O(N__39054),
            .I(N__39049));
    CascadeMux I__7612 (
            .O(N__39053),
            .I(N__39046));
    InMux I__7611 (
            .O(N__39052),
            .I(N__39043));
    InMux I__7610 (
            .O(N__39049),
            .I(N__39040));
    InMux I__7609 (
            .O(N__39046),
            .I(N__39037));
    LocalMux I__7608 (
            .O(N__39043),
            .I(dti_counter_6));
    LocalMux I__7607 (
            .O(N__39040),
            .I(dti_counter_6));
    LocalMux I__7606 (
            .O(N__39037),
            .I(dti_counter_6));
    CascadeMux I__7605 (
            .O(N__39030),
            .I(n14_adj_705_cascade_));
    InMux I__7604 (
            .O(N__39027),
            .I(N__39022));
    InMux I__7603 (
            .O(N__39026),
            .I(N__39017));
    InMux I__7602 (
            .O(N__39025),
            .I(N__39017));
    LocalMux I__7601 (
            .O(N__39022),
            .I(dti_counter_2));
    LocalMux I__7600 (
            .O(N__39017),
            .I(dti_counter_2));
    InMux I__7599 (
            .O(N__39012),
            .I(N__39009));
    LocalMux I__7598 (
            .O(N__39009),
            .I(n10_adj_706));
    CascadeMux I__7597 (
            .O(N__39006),
            .I(N__39003));
    InMux I__7596 (
            .O(N__39003),
            .I(N__38998));
    InMux I__7595 (
            .O(N__39002),
            .I(N__38995));
    InMux I__7594 (
            .O(N__39001),
            .I(N__38992));
    LocalMux I__7593 (
            .O(N__38998),
            .I(dti_counter_0));
    LocalMux I__7592 (
            .O(N__38995),
            .I(dti_counter_0));
    LocalMux I__7591 (
            .O(N__38992),
            .I(dti_counter_0));
    InMux I__7590 (
            .O(N__38985),
            .I(N__38982));
    LocalMux I__7589 (
            .O(N__38982),
            .I(n15081));
    CascadeMux I__7588 (
            .O(N__38979),
            .I(N__38976));
    InMux I__7587 (
            .O(N__38976),
            .I(N__38971));
    InMux I__7586 (
            .O(N__38975),
            .I(N__38966));
    InMux I__7585 (
            .O(N__38974),
            .I(N__38966));
    LocalMux I__7584 (
            .O(N__38971),
            .I(dti_counter_3));
    LocalMux I__7583 (
            .O(N__38966),
            .I(dti_counter_3));
    InMux I__7582 (
            .O(N__38961),
            .I(N__38958));
    LocalMux I__7581 (
            .O(N__38958),
            .I(n15074));
    CascadeMux I__7580 (
            .O(N__38955),
            .I(N__38951));
    InMux I__7579 (
            .O(N__38954),
            .I(N__38947));
    InMux I__7578 (
            .O(N__38951),
            .I(N__38942));
    InMux I__7577 (
            .O(N__38950),
            .I(N__38942));
    LocalMux I__7576 (
            .O(N__38947),
            .I(dti_counter_4));
    LocalMux I__7575 (
            .O(N__38942),
            .I(dti_counter_4));
    InMux I__7574 (
            .O(N__38937),
            .I(N__38934));
    LocalMux I__7573 (
            .O(N__38934),
            .I(n15073));
    CascadeMux I__7572 (
            .O(N__38931),
            .I(N__38928));
    InMux I__7571 (
            .O(N__38928),
            .I(N__38924));
    InMux I__7570 (
            .O(N__38927),
            .I(N__38920));
    LocalMux I__7569 (
            .O(N__38924),
            .I(N__38917));
    InMux I__7568 (
            .O(N__38923),
            .I(N__38914));
    LocalMux I__7567 (
            .O(N__38920),
            .I(dti_counter_7));
    Odrv4 I__7566 (
            .O(N__38917),
            .I(dti_counter_7));
    LocalMux I__7565 (
            .O(N__38914),
            .I(dti_counter_7));
    CascadeMux I__7564 (
            .O(N__38907),
            .I(N__38904));
    InMux I__7563 (
            .O(N__38904),
            .I(N__38901));
    LocalMux I__7562 (
            .O(N__38901),
            .I(N__38898));
    Odrv4 I__7561 (
            .O(N__38898),
            .I(n15070));
    InMux I__7560 (
            .O(N__38895),
            .I(N__38892));
    LocalMux I__7559 (
            .O(N__38892),
            .I(N__38889));
    Span4Mux_v I__7558 (
            .O(N__38889),
            .I(N__38886));
    Sp12to4 I__7557 (
            .O(N__38886),
            .I(N__38882));
    InMux I__7556 (
            .O(N__38885),
            .I(N__38879));
    Odrv12 I__7555 (
            .O(N__38882),
            .I(reg_B_1));
    LocalMux I__7554 (
            .O(N__38879),
            .I(reg_B_1));
    InMux I__7553 (
            .O(N__38874),
            .I(N__38871));
    LocalMux I__7552 (
            .O(N__38871),
            .I(N__38867));
    InMux I__7551 (
            .O(N__38870),
            .I(N__38864));
    Span4Mux_h I__7550 (
            .O(N__38867),
            .I(N__38861));
    LocalMux I__7549 (
            .O(N__38864),
            .I(N__38858));
    Span4Mux_h I__7548 (
            .O(N__38861),
            .I(N__38854));
    Span4Mux_v I__7547 (
            .O(N__38858),
            .I(N__38851));
    InMux I__7546 (
            .O(N__38857),
            .I(N__38848));
    Odrv4 I__7545 (
            .O(N__38854),
            .I(n14129));
    Odrv4 I__7544 (
            .O(N__38851),
            .I(n14129));
    LocalMux I__7543 (
            .O(N__38848),
            .I(n14129));
    CascadeMux I__7542 (
            .O(N__38841),
            .I(N__38838));
    InMux I__7541 (
            .O(N__38838),
            .I(N__38835));
    LocalMux I__7540 (
            .O(N__38835),
            .I(N__38832));
    Odrv4 I__7539 (
            .O(N__38832),
            .I(n1377));
    InMux I__7538 (
            .O(N__38829),
            .I(bfn_9_29_0_));
    InMux I__7537 (
            .O(N__38826),
            .I(n13006));
    InMux I__7536 (
            .O(N__38823),
            .I(n13007));
    InMux I__7535 (
            .O(N__38820),
            .I(n13008));
    InMux I__7534 (
            .O(N__38817),
            .I(n13009));
    InMux I__7533 (
            .O(N__38814),
            .I(N__38811));
    LocalMux I__7532 (
            .O(N__38811),
            .I(n15072));
    InMux I__7531 (
            .O(N__38808),
            .I(n13010));
    InMux I__7530 (
            .O(N__38805),
            .I(n13011));
    CascadeMux I__7529 (
            .O(N__38802),
            .I(N__38796));
    CascadeMux I__7528 (
            .O(N__38801),
            .I(N__38792));
    CascadeMux I__7527 (
            .O(N__38800),
            .I(N__38788));
    InMux I__7526 (
            .O(N__38799),
            .I(N__38772));
    InMux I__7525 (
            .O(N__38796),
            .I(N__38772));
    InMux I__7524 (
            .O(N__38795),
            .I(N__38772));
    InMux I__7523 (
            .O(N__38792),
            .I(N__38772));
    InMux I__7522 (
            .O(N__38791),
            .I(N__38772));
    InMux I__7521 (
            .O(N__38788),
            .I(N__38772));
    InMux I__7520 (
            .O(N__38787),
            .I(N__38772));
    LocalMux I__7519 (
            .O(N__38772),
            .I(N__38769));
    Odrv4 I__7518 (
            .O(N__38769),
            .I(n11526));
    InMux I__7517 (
            .O(N__38766),
            .I(n13012));
    InMux I__7516 (
            .O(N__38763),
            .I(N__38760));
    LocalMux I__7515 (
            .O(N__38760),
            .I(N__38757));
    Odrv4 I__7514 (
            .O(N__38757),
            .I(encoder0_position_scaled_18));
    InMux I__7513 (
            .O(N__38754),
            .I(N__38751));
    LocalMux I__7512 (
            .O(N__38751),
            .I(N__38748));
    Odrv4 I__7511 (
            .O(N__38748),
            .I(encoder0_position_scaled_23));
    InMux I__7510 (
            .O(N__38745),
            .I(N__38742));
    LocalMux I__7509 (
            .O(N__38742),
            .I(N__38739));
    Odrv4 I__7508 (
            .O(N__38739),
            .I(encoder0_position_scaled_17));
    CascadeMux I__7507 (
            .O(N__38736),
            .I(dti_N_333_cascade_));
    InMux I__7506 (
            .O(N__38733),
            .I(n13004));
    InMux I__7505 (
            .O(N__38730),
            .I(n13005));
    InMux I__7504 (
            .O(N__38727),
            .I(N__38724));
    LocalMux I__7503 (
            .O(N__38724),
            .I(N__38721));
    Odrv4 I__7502 (
            .O(N__38721),
            .I(encoder0_position_scaled_8));
    InMux I__7501 (
            .O(N__38718),
            .I(N__38715));
    LocalMux I__7500 (
            .O(N__38715),
            .I(N__38712));
    Odrv4 I__7499 (
            .O(N__38712),
            .I(encoder0_position_scaled_14));
    InMux I__7498 (
            .O(N__38709),
            .I(N__38706));
    LocalMux I__7497 (
            .O(N__38706),
            .I(N__38703));
    Odrv4 I__7496 (
            .O(N__38703),
            .I(encoder0_position_scaled_10));
    InMux I__7495 (
            .O(N__38700),
            .I(N__38697));
    LocalMux I__7494 (
            .O(N__38697),
            .I(N__38694));
    Odrv4 I__7493 (
            .O(N__38694),
            .I(encoder0_position_scaled_12));
    InMux I__7492 (
            .O(N__38691),
            .I(N__38688));
    LocalMux I__7491 (
            .O(N__38688),
            .I(N__38685));
    Odrv4 I__7490 (
            .O(N__38685),
            .I(encoder0_position_scaled_13));
    InMux I__7489 (
            .O(N__38682),
            .I(N__38679));
    LocalMux I__7488 (
            .O(N__38679),
            .I(N__38676));
    Odrv4 I__7487 (
            .O(N__38676),
            .I(encoder0_position_scaled_15));
    InMux I__7486 (
            .O(N__38673),
            .I(N__38670));
    LocalMux I__7485 (
            .O(N__38670),
            .I(N__38667));
    Odrv4 I__7484 (
            .O(N__38667),
            .I(n15508));
    InMux I__7483 (
            .O(N__38664),
            .I(n12995));
    InMux I__7482 (
            .O(N__38661),
            .I(n12996));
    InMux I__7481 (
            .O(N__38658),
            .I(n12997));
    InMux I__7480 (
            .O(N__38655),
            .I(bfn_9_25_0_));
    InMux I__7479 (
            .O(N__38652),
            .I(n12999));
    InMux I__7478 (
            .O(N__38649),
            .I(n13000));
    InMux I__7477 (
            .O(N__38646),
            .I(n13001));
    InMux I__7476 (
            .O(N__38643),
            .I(n13002));
    InMux I__7475 (
            .O(N__38640),
            .I(N__38637));
    LocalMux I__7474 (
            .O(N__38637),
            .I(N__38634));
    Span4Mux_v I__7473 (
            .O(N__38634),
            .I(N__38631));
    Odrv4 I__7472 (
            .O(N__38631),
            .I(n4_adj_622));
    InMux I__7471 (
            .O(N__38628),
            .I(n13003));
    InMux I__7470 (
            .O(N__38625),
            .I(N__38622));
    LocalMux I__7469 (
            .O(N__38622),
            .I(N__38619));
    Span4Mux_h I__7468 (
            .O(N__38619),
            .I(N__38616));
    Odrv4 I__7467 (
            .O(N__38616),
            .I(n20));
    InMux I__7466 (
            .O(N__38613),
            .I(n12987));
    CascadeMux I__7465 (
            .O(N__38610),
            .I(N__38607));
    InMux I__7464 (
            .O(N__38607),
            .I(N__38604));
    LocalMux I__7463 (
            .O(N__38604),
            .I(N__38601));
    Odrv4 I__7462 (
            .O(N__38601),
            .I(n19_adj_637));
    InMux I__7461 (
            .O(N__38598),
            .I(N__38595));
    LocalMux I__7460 (
            .O(N__38595),
            .I(N__38592));
    Odrv12 I__7459 (
            .O(N__38592),
            .I(n19));
    InMux I__7458 (
            .O(N__38589),
            .I(n12988));
    CascadeMux I__7457 (
            .O(N__38586),
            .I(N__38583));
    InMux I__7456 (
            .O(N__38583),
            .I(N__38580));
    LocalMux I__7455 (
            .O(N__38580),
            .I(N__38577));
    Odrv4 I__7454 (
            .O(N__38577),
            .I(n18_adj_636));
    InMux I__7453 (
            .O(N__38574),
            .I(N__38571));
    LocalMux I__7452 (
            .O(N__38571),
            .I(N__38568));
    Span4Mux_h I__7451 (
            .O(N__38568),
            .I(N__38565));
    Odrv4 I__7450 (
            .O(N__38565),
            .I(n18));
    InMux I__7449 (
            .O(N__38562),
            .I(n12989));
    InMux I__7448 (
            .O(N__38559),
            .I(bfn_9_24_0_));
    InMux I__7447 (
            .O(N__38556),
            .I(n12991));
    InMux I__7446 (
            .O(N__38553),
            .I(n12992));
    CascadeMux I__7445 (
            .O(N__38550),
            .I(N__38547));
    InMux I__7444 (
            .O(N__38547),
            .I(N__38544));
    LocalMux I__7443 (
            .O(N__38544),
            .I(N__38541));
    Odrv12 I__7442 (
            .O(N__38541),
            .I(n14_adj_632));
    InMux I__7441 (
            .O(N__38538),
            .I(N__38535));
    LocalMux I__7440 (
            .O(N__38535),
            .I(N__38532));
    Odrv12 I__7439 (
            .O(N__38532),
            .I(n14));
    InMux I__7438 (
            .O(N__38529),
            .I(n12993));
    InMux I__7437 (
            .O(N__38526),
            .I(n12994));
    CascadeMux I__7436 (
            .O(N__38523),
            .I(N__38520));
    InMux I__7435 (
            .O(N__38520),
            .I(N__38517));
    LocalMux I__7434 (
            .O(N__38517),
            .I(N__38514));
    Odrv12 I__7433 (
            .O(N__38514),
            .I(n28_adj_646));
    InMux I__7432 (
            .O(N__38511),
            .I(N__38508));
    LocalMux I__7431 (
            .O(N__38508),
            .I(N__38505));
    Odrv4 I__7430 (
            .O(N__38505),
            .I(n28));
    InMux I__7429 (
            .O(N__38502),
            .I(n12979));
    CascadeMux I__7428 (
            .O(N__38499),
            .I(N__38496));
    InMux I__7427 (
            .O(N__38496),
            .I(N__38493));
    LocalMux I__7426 (
            .O(N__38493),
            .I(n27_adj_645));
    InMux I__7425 (
            .O(N__38490),
            .I(N__38487));
    LocalMux I__7424 (
            .O(N__38487),
            .I(N__38484));
    Odrv4 I__7423 (
            .O(N__38484),
            .I(n27));
    InMux I__7422 (
            .O(N__38481),
            .I(n12980));
    CascadeMux I__7421 (
            .O(N__38478),
            .I(N__38475));
    InMux I__7420 (
            .O(N__38475),
            .I(N__38472));
    LocalMux I__7419 (
            .O(N__38472),
            .I(n26_adj_644));
    InMux I__7418 (
            .O(N__38469),
            .I(N__38466));
    LocalMux I__7417 (
            .O(N__38466),
            .I(N__38463));
    Span4Mux_h I__7416 (
            .O(N__38463),
            .I(N__38460));
    Odrv4 I__7415 (
            .O(N__38460),
            .I(n26));
    InMux I__7414 (
            .O(N__38457),
            .I(n12981));
    CascadeMux I__7413 (
            .O(N__38454),
            .I(N__38451));
    InMux I__7412 (
            .O(N__38451),
            .I(N__38448));
    LocalMux I__7411 (
            .O(N__38448),
            .I(N__38445));
    Odrv4 I__7410 (
            .O(N__38445),
            .I(n25_adj_643));
    InMux I__7409 (
            .O(N__38442),
            .I(N__38439));
    LocalMux I__7408 (
            .O(N__38439),
            .I(N__38436));
    Span4Mux_h I__7407 (
            .O(N__38436),
            .I(N__38433));
    Odrv4 I__7406 (
            .O(N__38433),
            .I(n25));
    InMux I__7405 (
            .O(N__38430),
            .I(bfn_9_23_0_));
    CascadeMux I__7404 (
            .O(N__38427),
            .I(N__38424));
    InMux I__7403 (
            .O(N__38424),
            .I(N__38421));
    LocalMux I__7402 (
            .O(N__38421),
            .I(N__38418));
    Odrv4 I__7401 (
            .O(N__38418),
            .I(n24_adj_642));
    InMux I__7400 (
            .O(N__38415),
            .I(N__38412));
    LocalMux I__7399 (
            .O(N__38412),
            .I(N__38409));
    Span4Mux_v I__7398 (
            .O(N__38409),
            .I(N__38406));
    Odrv4 I__7397 (
            .O(N__38406),
            .I(n24));
    InMux I__7396 (
            .O(N__38403),
            .I(n12983));
    CascadeMux I__7395 (
            .O(N__38400),
            .I(N__38397));
    InMux I__7394 (
            .O(N__38397),
            .I(N__38394));
    LocalMux I__7393 (
            .O(N__38394),
            .I(N__38391));
    Odrv4 I__7392 (
            .O(N__38391),
            .I(n23_adj_641));
    InMux I__7391 (
            .O(N__38388),
            .I(N__38385));
    LocalMux I__7390 (
            .O(N__38385),
            .I(N__38382));
    Odrv4 I__7389 (
            .O(N__38382),
            .I(n23));
    InMux I__7388 (
            .O(N__38379),
            .I(n12984));
    InMux I__7387 (
            .O(N__38376),
            .I(N__38373));
    LocalMux I__7386 (
            .O(N__38373),
            .I(N__38370));
    Odrv4 I__7385 (
            .O(N__38370),
            .I(n22));
    InMux I__7384 (
            .O(N__38367),
            .I(n12985));
    InMux I__7383 (
            .O(N__38364),
            .I(N__38361));
    LocalMux I__7382 (
            .O(N__38361),
            .I(N__38358));
    Span4Mux_h I__7381 (
            .O(N__38358),
            .I(N__38355));
    Odrv4 I__7380 (
            .O(N__38355),
            .I(n21));
    InMux I__7379 (
            .O(N__38352),
            .I(n12986));
    InMux I__7378 (
            .O(N__38349),
            .I(N__38346));
    LocalMux I__7377 (
            .O(N__38346),
            .I(N__38341));
    InMux I__7376 (
            .O(N__38345),
            .I(N__38338));
    InMux I__7375 (
            .O(N__38344),
            .I(N__38335));
    Span4Mux_v I__7374 (
            .O(N__38341),
            .I(N__38330));
    LocalMux I__7373 (
            .O(N__38338),
            .I(N__38330));
    LocalMux I__7372 (
            .O(N__38335),
            .I(N__38327));
    Span4Mux_h I__7371 (
            .O(N__38330),
            .I(N__38324));
    Span4Mux_h I__7370 (
            .O(N__38327),
            .I(N__38321));
    Span4Mux_h I__7369 (
            .O(N__38324),
            .I(N__38318));
    Odrv4 I__7368 (
            .O(N__38321),
            .I(n309));
    Odrv4 I__7367 (
            .O(N__38318),
            .I(n309));
    CascadeMux I__7366 (
            .O(N__38313),
            .I(N__38310));
    InMux I__7365 (
            .O(N__38310),
            .I(N__38307));
    LocalMux I__7364 (
            .O(N__38307),
            .I(N__38304));
    Odrv4 I__7363 (
            .O(N__38304),
            .I(n33_adj_651));
    InMux I__7362 (
            .O(N__38301),
            .I(N__38298));
    LocalMux I__7361 (
            .O(N__38298),
            .I(N__38295));
    Span4Mux_h I__7360 (
            .O(N__38295),
            .I(N__38292));
    Odrv4 I__7359 (
            .O(N__38292),
            .I(n33));
    InMux I__7358 (
            .O(N__38289),
            .I(bfn_9_22_0_));
    InMux I__7357 (
            .O(N__38286),
            .I(N__38283));
    LocalMux I__7356 (
            .O(N__38283),
            .I(N__38280));
    Odrv12 I__7355 (
            .O(N__38280),
            .I(n32));
    InMux I__7354 (
            .O(N__38277),
            .I(n12975));
    CascadeMux I__7353 (
            .O(N__38274),
            .I(N__38271));
    InMux I__7352 (
            .O(N__38271),
            .I(N__38268));
    LocalMux I__7351 (
            .O(N__38268),
            .I(N__38265));
    Odrv12 I__7350 (
            .O(N__38265),
            .I(n31_adj_649));
    InMux I__7349 (
            .O(N__38262),
            .I(N__38259));
    LocalMux I__7348 (
            .O(N__38259),
            .I(N__38256));
    Span4Mux_h I__7347 (
            .O(N__38256),
            .I(N__38253));
    Odrv4 I__7346 (
            .O(N__38253),
            .I(n31));
    InMux I__7345 (
            .O(N__38250),
            .I(n12976));
    CascadeMux I__7344 (
            .O(N__38247),
            .I(N__38244));
    InMux I__7343 (
            .O(N__38244),
            .I(N__38241));
    LocalMux I__7342 (
            .O(N__38241),
            .I(n30_adj_648));
    InMux I__7341 (
            .O(N__38238),
            .I(n12977));
    CascadeMux I__7340 (
            .O(N__38235),
            .I(N__38232));
    InMux I__7339 (
            .O(N__38232),
            .I(N__38229));
    LocalMux I__7338 (
            .O(N__38229),
            .I(n29_adj_647));
    InMux I__7337 (
            .O(N__38226),
            .I(N__38223));
    LocalMux I__7336 (
            .O(N__38223),
            .I(N__38220));
    Span4Mux_h I__7335 (
            .O(N__38220),
            .I(N__38217));
    Odrv4 I__7334 (
            .O(N__38217),
            .I(n29));
    InMux I__7333 (
            .O(N__38214),
            .I(n12978));
    InMux I__7332 (
            .O(N__38211),
            .I(N__38207));
    InMux I__7331 (
            .O(N__38210),
            .I(N__38203));
    LocalMux I__7330 (
            .O(N__38207),
            .I(N__38200));
    InMux I__7329 (
            .O(N__38206),
            .I(N__38197));
    LocalMux I__7328 (
            .O(N__38203),
            .I(N__38194));
    Span4Mux_h I__7327 (
            .O(N__38200),
            .I(N__38191));
    LocalMux I__7326 (
            .O(N__38197),
            .I(N__38188));
    Span4Mux_h I__7325 (
            .O(N__38194),
            .I(N__38185));
    Span4Mux_h I__7324 (
            .O(N__38191),
            .I(N__38182));
    Span12Mux_s8_h I__7323 (
            .O(N__38188),
            .I(N__38179));
    Span4Mux_v I__7322 (
            .O(N__38185),
            .I(N__38176));
    Odrv4 I__7321 (
            .O(N__38182),
            .I(n308));
    Odrv12 I__7320 (
            .O(N__38179),
            .I(n308));
    Odrv4 I__7319 (
            .O(N__38176),
            .I(n308));
    InMux I__7318 (
            .O(N__38169),
            .I(N__38166));
    LocalMux I__7317 (
            .O(N__38166),
            .I(N__38163));
    Odrv4 I__7316 (
            .O(N__38163),
            .I(n14530));
    InMux I__7315 (
            .O(N__38160),
            .I(N__38153));
    InMux I__7314 (
            .O(N__38159),
            .I(N__38153));
    InMux I__7313 (
            .O(N__38158),
            .I(N__38150));
    LocalMux I__7312 (
            .O(N__38153),
            .I(N__38147));
    LocalMux I__7311 (
            .O(N__38150),
            .I(n1918));
    Odrv4 I__7310 (
            .O(N__38147),
            .I(n1918));
    InMux I__7309 (
            .O(N__38142),
            .I(N__38139));
    LocalMux I__7308 (
            .O(N__38139),
            .I(N__38134));
    InMux I__7307 (
            .O(N__38138),
            .I(N__38131));
    InMux I__7306 (
            .O(N__38137),
            .I(N__38128));
    Span4Mux_v I__7305 (
            .O(N__38134),
            .I(N__38123));
    LocalMux I__7304 (
            .O(N__38131),
            .I(N__38123));
    LocalMux I__7303 (
            .O(N__38128),
            .I(n1919));
    Odrv4 I__7302 (
            .O(N__38123),
            .I(n1919));
    InMux I__7301 (
            .O(N__38118),
            .I(N__38114));
    InMux I__7300 (
            .O(N__38117),
            .I(N__38111));
    LocalMux I__7299 (
            .O(N__38114),
            .I(N__38108));
    LocalMux I__7298 (
            .O(N__38111),
            .I(N__38102));
    Span4Mux_v I__7297 (
            .O(N__38108),
            .I(N__38102));
    InMux I__7296 (
            .O(N__38107),
            .I(N__38099));
    Span4Mux_h I__7295 (
            .O(N__38102),
            .I(N__38096));
    LocalMux I__7294 (
            .O(N__38099),
            .I(N__38093));
    Odrv4 I__7293 (
            .O(N__38096),
            .I(n305));
    Odrv4 I__7292 (
            .O(N__38093),
            .I(n305));
    InMux I__7291 (
            .O(N__38088),
            .I(N__38084));
    InMux I__7290 (
            .O(N__38087),
            .I(N__38081));
    LocalMux I__7289 (
            .O(N__38084),
            .I(N__38075));
    LocalMux I__7288 (
            .O(N__38081),
            .I(N__38075));
    InMux I__7287 (
            .O(N__38080),
            .I(N__38072));
    Span4Mux_v I__7286 (
            .O(N__38075),
            .I(N__38067));
    LocalMux I__7285 (
            .O(N__38072),
            .I(N__38067));
    Odrv4 I__7284 (
            .O(N__38067),
            .I(n306));
    InMux I__7283 (
            .O(N__38064),
            .I(N__38061));
    LocalMux I__7282 (
            .O(N__38061),
            .I(N__38058));
    Span4Mux_v I__7281 (
            .O(N__38058),
            .I(N__38055));
    Odrv4 I__7280 (
            .O(N__38055),
            .I(n1991));
    InMux I__7279 (
            .O(N__38052),
            .I(n12631));
    InMux I__7278 (
            .O(N__38049),
            .I(N__38046));
    LocalMux I__7277 (
            .O(N__38046),
            .I(N__38043));
    Span4Mux_v I__7276 (
            .O(N__38043),
            .I(N__38040));
    Odrv4 I__7275 (
            .O(N__38040),
            .I(n1990));
    InMux I__7274 (
            .O(N__38037),
            .I(n12632));
    CascadeMux I__7273 (
            .O(N__38034),
            .I(N__38031));
    InMux I__7272 (
            .O(N__38031),
            .I(N__38028));
    LocalMux I__7271 (
            .O(N__38028),
            .I(N__38024));
    InMux I__7270 (
            .O(N__38027),
            .I(N__38021));
    Odrv4 I__7269 (
            .O(N__38024),
            .I(n1922));
    LocalMux I__7268 (
            .O(N__38021),
            .I(n1922));
    InMux I__7267 (
            .O(N__38016),
            .I(N__38013));
    LocalMux I__7266 (
            .O(N__38013),
            .I(N__38010));
    Odrv4 I__7265 (
            .O(N__38010),
            .I(n1989));
    InMux I__7264 (
            .O(N__38007),
            .I(n12633));
    CascadeMux I__7263 (
            .O(N__38004),
            .I(N__38001));
    InMux I__7262 (
            .O(N__38001),
            .I(N__37998));
    LocalMux I__7261 (
            .O(N__37998),
            .I(N__37995));
    Odrv4 I__7260 (
            .O(N__37995),
            .I(n1988));
    InMux I__7259 (
            .O(N__37992),
            .I(n12634));
    InMux I__7258 (
            .O(N__37989),
            .I(n12635));
    CascadeMux I__7257 (
            .O(N__37986),
            .I(N__37983));
    InMux I__7256 (
            .O(N__37983),
            .I(N__37980));
    LocalMux I__7255 (
            .O(N__37980),
            .I(N__37977));
    Span4Mux_h I__7254 (
            .O(N__37977),
            .I(N__37974));
    Odrv4 I__7253 (
            .O(N__37974),
            .I(n1986));
    InMux I__7252 (
            .O(N__37971),
            .I(n12636));
    InMux I__7251 (
            .O(N__37968),
            .I(N__37965));
    LocalMux I__7250 (
            .O(N__37965),
            .I(N__37962));
    Span4Mux_h I__7249 (
            .O(N__37962),
            .I(N__37959));
    Odrv4 I__7248 (
            .O(N__37959),
            .I(n1985));
    InMux I__7247 (
            .O(N__37956),
            .I(bfn_9_18_0_));
    CascadeMux I__7246 (
            .O(N__37953),
            .I(N__37949));
    InMux I__7245 (
            .O(N__37952),
            .I(N__37946));
    InMux I__7244 (
            .O(N__37949),
            .I(N__37943));
    LocalMux I__7243 (
            .O(N__37946),
            .I(N__37940));
    LocalMux I__7242 (
            .O(N__37943),
            .I(N__37937));
    Odrv12 I__7241 (
            .O(N__37940),
            .I(n15674));
    Odrv4 I__7240 (
            .O(N__37937),
            .I(n15674));
    InMux I__7239 (
            .O(N__37932),
            .I(n12638));
    CascadeMux I__7238 (
            .O(N__37929),
            .I(N__37926));
    InMux I__7237 (
            .O(N__37926),
            .I(N__37920));
    InMux I__7236 (
            .O(N__37925),
            .I(N__37920));
    LocalMux I__7235 (
            .O(N__37920),
            .I(N__37917));
    Span4Mux_h I__7234 (
            .O(N__37917),
            .I(N__37914));
    Odrv4 I__7233 (
            .O(N__37914),
            .I(n2016));
    InMux I__7232 (
            .O(N__37911),
            .I(N__37908));
    LocalMux I__7231 (
            .O(N__37908),
            .I(N__37903));
    CascadeMux I__7230 (
            .O(N__37907),
            .I(N__37900));
    InMux I__7229 (
            .O(N__37906),
            .I(N__37897));
    Span4Mux_h I__7228 (
            .O(N__37903),
            .I(N__37894));
    InMux I__7227 (
            .O(N__37900),
            .I(N__37891));
    LocalMux I__7226 (
            .O(N__37897),
            .I(N__37888));
    Odrv4 I__7225 (
            .O(N__37894),
            .I(n1921));
    LocalMux I__7224 (
            .O(N__37891),
            .I(n1921));
    Odrv4 I__7223 (
            .O(N__37888),
            .I(n1921));
    InMux I__7222 (
            .O(N__37881),
            .I(N__37878));
    LocalMux I__7221 (
            .O(N__37878),
            .I(N__37875));
    Span4Mux_v I__7220 (
            .O(N__37875),
            .I(N__37872));
    Odrv4 I__7219 (
            .O(N__37872),
            .I(n1999));
    InMux I__7218 (
            .O(N__37869),
            .I(n12623));
    InMux I__7217 (
            .O(N__37866),
            .I(N__37863));
    LocalMux I__7216 (
            .O(N__37863),
            .I(N__37860));
    Odrv4 I__7215 (
            .O(N__37860),
            .I(n1998));
    InMux I__7214 (
            .O(N__37857),
            .I(n12624));
    CascadeMux I__7213 (
            .O(N__37854),
            .I(N__37851));
    InMux I__7212 (
            .O(N__37851),
            .I(N__37848));
    LocalMux I__7211 (
            .O(N__37848),
            .I(N__37845));
    Span4Mux_v I__7210 (
            .O(N__37845),
            .I(N__37842));
    Odrv4 I__7209 (
            .O(N__37842),
            .I(n1997));
    InMux I__7208 (
            .O(N__37839),
            .I(n12625));
    CascadeMux I__7207 (
            .O(N__37836),
            .I(N__37833));
    InMux I__7206 (
            .O(N__37833),
            .I(N__37830));
    LocalMux I__7205 (
            .O(N__37830),
            .I(N__37827));
    Span4Mux_h I__7204 (
            .O(N__37827),
            .I(N__37824));
    Odrv4 I__7203 (
            .O(N__37824),
            .I(n1996));
    InMux I__7202 (
            .O(N__37821),
            .I(n12626));
    CascadeMux I__7201 (
            .O(N__37818),
            .I(N__37815));
    InMux I__7200 (
            .O(N__37815),
            .I(N__37812));
    LocalMux I__7199 (
            .O(N__37812),
            .I(N__37809));
    Span4Mux_h I__7198 (
            .O(N__37809),
            .I(N__37806));
    Odrv4 I__7197 (
            .O(N__37806),
            .I(n1995));
    InMux I__7196 (
            .O(N__37803),
            .I(n12627));
    InMux I__7195 (
            .O(N__37800),
            .I(N__37797));
    LocalMux I__7194 (
            .O(N__37797),
            .I(N__37794));
    Span4Mux_h I__7193 (
            .O(N__37794),
            .I(N__37791));
    Odrv4 I__7192 (
            .O(N__37791),
            .I(n1994));
    InMux I__7191 (
            .O(N__37788),
            .I(n12628));
    InMux I__7190 (
            .O(N__37785),
            .I(N__37782));
    LocalMux I__7189 (
            .O(N__37782),
            .I(N__37779));
    Span4Mux_h I__7188 (
            .O(N__37779),
            .I(N__37776));
    Odrv4 I__7187 (
            .O(N__37776),
            .I(n1993));
    InMux I__7186 (
            .O(N__37773),
            .I(bfn_9_17_0_));
    InMux I__7185 (
            .O(N__37770),
            .I(N__37767));
    LocalMux I__7184 (
            .O(N__37767),
            .I(N__37764));
    Span4Mux_h I__7183 (
            .O(N__37764),
            .I(N__37761));
    Odrv4 I__7182 (
            .O(N__37761),
            .I(n1992));
    InMux I__7181 (
            .O(N__37758),
            .I(n12630));
    InMux I__7180 (
            .O(N__37755),
            .I(N__37750));
    InMux I__7179 (
            .O(N__37754),
            .I(N__37747));
    InMux I__7178 (
            .O(N__37753),
            .I(N__37744));
    LocalMux I__7177 (
            .O(N__37750),
            .I(N__37741));
    LocalMux I__7176 (
            .O(N__37747),
            .I(N__37736));
    LocalMux I__7175 (
            .O(N__37744),
            .I(N__37736));
    Odrv4 I__7174 (
            .O(N__37741),
            .I(n3209));
    Odrv4 I__7173 (
            .O(N__37736),
            .I(n3209));
    CascadeMux I__7172 (
            .O(N__37731),
            .I(N__37728));
    InMux I__7171 (
            .O(N__37728),
            .I(N__37725));
    LocalMux I__7170 (
            .O(N__37725),
            .I(N__37722));
    Odrv4 I__7169 (
            .O(N__37722),
            .I(n3276));
    InMux I__7168 (
            .O(N__37719),
            .I(n12946));
    CascadeMux I__7167 (
            .O(N__37716),
            .I(N__37711));
    InMux I__7166 (
            .O(N__37715),
            .I(N__37708));
    InMux I__7165 (
            .O(N__37714),
            .I(N__37705));
    InMux I__7164 (
            .O(N__37711),
            .I(N__37702));
    LocalMux I__7163 (
            .O(N__37708),
            .I(N__37699));
    LocalMux I__7162 (
            .O(N__37705),
            .I(N__37694));
    LocalMux I__7161 (
            .O(N__37702),
            .I(N__37694));
    Odrv4 I__7160 (
            .O(N__37699),
            .I(n3208));
    Odrv4 I__7159 (
            .O(N__37694),
            .I(n3208));
    InMux I__7158 (
            .O(N__37689),
            .I(N__37686));
    LocalMux I__7157 (
            .O(N__37686),
            .I(N__37683));
    Odrv4 I__7156 (
            .O(N__37683),
            .I(n3275));
    InMux I__7155 (
            .O(N__37680),
            .I(n12947));
    InMux I__7154 (
            .O(N__37677),
            .I(N__37674));
    LocalMux I__7153 (
            .O(N__37674),
            .I(N__37669));
    InMux I__7152 (
            .O(N__37673),
            .I(N__37664));
    InMux I__7151 (
            .O(N__37672),
            .I(N__37664));
    Span4Mux_s2_v I__7150 (
            .O(N__37669),
            .I(N__37659));
    LocalMux I__7149 (
            .O(N__37664),
            .I(N__37659));
    Span4Mux_h I__7148 (
            .O(N__37659),
            .I(N__37656));
    Odrv4 I__7147 (
            .O(N__37656),
            .I(n3207));
    InMux I__7146 (
            .O(N__37653),
            .I(N__37650));
    LocalMux I__7145 (
            .O(N__37650),
            .I(N__37647));
    Odrv4 I__7144 (
            .O(N__37647),
            .I(n3274));
    InMux I__7143 (
            .O(N__37644),
            .I(n12948));
    InMux I__7142 (
            .O(N__37641),
            .I(N__37636));
    InMux I__7141 (
            .O(N__37640),
            .I(N__37633));
    InMux I__7140 (
            .O(N__37639),
            .I(N__37630));
    LocalMux I__7139 (
            .O(N__37636),
            .I(N__37627));
    LocalMux I__7138 (
            .O(N__37633),
            .I(N__37624));
    LocalMux I__7137 (
            .O(N__37630),
            .I(N__37621));
    Span4Mux_v I__7136 (
            .O(N__37627),
            .I(N__37614));
    Span4Mux_h I__7135 (
            .O(N__37624),
            .I(N__37614));
    Span4Mux_v I__7134 (
            .O(N__37621),
            .I(N__37614));
    Odrv4 I__7133 (
            .O(N__37614),
            .I(n3206));
    InMux I__7132 (
            .O(N__37611),
            .I(N__37608));
    LocalMux I__7131 (
            .O(N__37608),
            .I(N__37605));
    Odrv4 I__7130 (
            .O(N__37605),
            .I(n3273));
    InMux I__7129 (
            .O(N__37602),
            .I(n12949));
    InMux I__7128 (
            .O(N__37599),
            .I(N__37595));
    InMux I__7127 (
            .O(N__37598),
            .I(N__37591));
    LocalMux I__7126 (
            .O(N__37595),
            .I(N__37588));
    InMux I__7125 (
            .O(N__37594),
            .I(N__37585));
    LocalMux I__7124 (
            .O(N__37591),
            .I(N__37582));
    Span4Mux_v I__7123 (
            .O(N__37588),
            .I(N__37579));
    LocalMux I__7122 (
            .O(N__37585),
            .I(N__37576));
    Span4Mux_h I__7121 (
            .O(N__37582),
            .I(N__37573));
    Odrv4 I__7120 (
            .O(N__37579),
            .I(n3205));
    Odrv12 I__7119 (
            .O(N__37576),
            .I(n3205));
    Odrv4 I__7118 (
            .O(N__37573),
            .I(n3205));
    InMux I__7117 (
            .O(N__37566),
            .I(N__37563));
    LocalMux I__7116 (
            .O(N__37563),
            .I(N__37560));
    Odrv4 I__7115 (
            .O(N__37560),
            .I(n3272));
    InMux I__7114 (
            .O(N__37557),
            .I(n12950));
    InMux I__7113 (
            .O(N__37554),
            .I(N__37551));
    LocalMux I__7112 (
            .O(N__37551),
            .I(N__37546));
    InMux I__7111 (
            .O(N__37550),
            .I(N__37543));
    InMux I__7110 (
            .O(N__37549),
            .I(N__37540));
    Span4Mux_v I__7109 (
            .O(N__37546),
            .I(N__37535));
    LocalMux I__7108 (
            .O(N__37543),
            .I(N__37535));
    LocalMux I__7107 (
            .O(N__37540),
            .I(N__37532));
    Span4Mux_h I__7106 (
            .O(N__37535),
            .I(N__37529));
    Odrv12 I__7105 (
            .O(N__37532),
            .I(n3204));
    Odrv4 I__7104 (
            .O(N__37529),
            .I(n3204));
    InMux I__7103 (
            .O(N__37524),
            .I(n12951));
    CascadeMux I__7102 (
            .O(N__37521),
            .I(N__37518));
    InMux I__7101 (
            .O(N__37518),
            .I(N__37515));
    LocalMux I__7100 (
            .O(N__37515),
            .I(N__37512));
    Span4Mux_h I__7099 (
            .O(N__37512),
            .I(N__37509));
    Odrv4 I__7098 (
            .O(N__37509),
            .I(n3271));
    InMux I__7097 (
            .O(N__37506),
            .I(N__37503));
    LocalMux I__7096 (
            .O(N__37503),
            .I(N__37500));
    Span4Mux_v I__7095 (
            .O(N__37500),
            .I(N__37497));
    Odrv4 I__7094 (
            .O(N__37497),
            .I(n2001));
    InMux I__7093 (
            .O(N__37494),
            .I(bfn_9_16_0_));
    CascadeMux I__7092 (
            .O(N__37491),
            .I(N__37488));
    InMux I__7091 (
            .O(N__37488),
            .I(N__37485));
    LocalMux I__7090 (
            .O(N__37485),
            .I(N__37482));
    Span4Mux_v I__7089 (
            .O(N__37482),
            .I(N__37479));
    Odrv4 I__7088 (
            .O(N__37479),
            .I(n2000));
    InMux I__7087 (
            .O(N__37476),
            .I(n12622));
    InMux I__7086 (
            .O(N__37473),
            .I(N__37468));
    CascadeMux I__7085 (
            .O(N__37472),
            .I(N__37465));
    InMux I__7084 (
            .O(N__37471),
            .I(N__37462));
    LocalMux I__7083 (
            .O(N__37468),
            .I(N__37459));
    InMux I__7082 (
            .O(N__37465),
            .I(N__37456));
    LocalMux I__7081 (
            .O(N__37462),
            .I(n3217));
    Odrv4 I__7080 (
            .O(N__37459),
            .I(n3217));
    LocalMux I__7079 (
            .O(N__37456),
            .I(n3217));
    InMux I__7078 (
            .O(N__37449),
            .I(N__37446));
    LocalMux I__7077 (
            .O(N__37446),
            .I(N__37443));
    Odrv4 I__7076 (
            .O(N__37443),
            .I(n3284));
    InMux I__7075 (
            .O(N__37440),
            .I(n12938));
    InMux I__7074 (
            .O(N__37437),
            .I(N__37433));
    InMux I__7073 (
            .O(N__37436),
            .I(N__37429));
    LocalMux I__7072 (
            .O(N__37433),
            .I(N__37426));
    InMux I__7071 (
            .O(N__37432),
            .I(N__37423));
    LocalMux I__7070 (
            .O(N__37429),
            .I(n3216));
    Odrv12 I__7069 (
            .O(N__37426),
            .I(n3216));
    LocalMux I__7068 (
            .O(N__37423),
            .I(n3216));
    InMux I__7067 (
            .O(N__37416),
            .I(N__37413));
    LocalMux I__7066 (
            .O(N__37413),
            .I(N__37410));
    Odrv4 I__7065 (
            .O(N__37410),
            .I(n3283));
    InMux I__7064 (
            .O(N__37407),
            .I(n12939));
    InMux I__7063 (
            .O(N__37404),
            .I(N__37400));
    InMux I__7062 (
            .O(N__37403),
            .I(N__37396));
    LocalMux I__7061 (
            .O(N__37400),
            .I(N__37393));
    InMux I__7060 (
            .O(N__37399),
            .I(N__37390));
    LocalMux I__7059 (
            .O(N__37396),
            .I(n3215));
    Odrv4 I__7058 (
            .O(N__37393),
            .I(n3215));
    LocalMux I__7057 (
            .O(N__37390),
            .I(n3215));
    InMux I__7056 (
            .O(N__37383),
            .I(N__37380));
    LocalMux I__7055 (
            .O(N__37380),
            .I(n3282));
    InMux I__7054 (
            .O(N__37377),
            .I(n12940));
    InMux I__7053 (
            .O(N__37374),
            .I(N__37370));
    InMux I__7052 (
            .O(N__37373),
            .I(N__37367));
    LocalMux I__7051 (
            .O(N__37370),
            .I(N__37361));
    LocalMux I__7050 (
            .O(N__37367),
            .I(N__37361));
    InMux I__7049 (
            .O(N__37366),
            .I(N__37358));
    Span4Mux_h I__7048 (
            .O(N__37361),
            .I(N__37353));
    LocalMux I__7047 (
            .O(N__37358),
            .I(N__37353));
    Odrv4 I__7046 (
            .O(N__37353),
            .I(n3214));
    InMux I__7045 (
            .O(N__37350),
            .I(N__37347));
    LocalMux I__7044 (
            .O(N__37347),
            .I(n3281));
    InMux I__7043 (
            .O(N__37344),
            .I(n12941));
    InMux I__7042 (
            .O(N__37341),
            .I(N__37337));
    InMux I__7041 (
            .O(N__37340),
            .I(N__37334));
    LocalMux I__7040 (
            .O(N__37337),
            .I(N__37328));
    LocalMux I__7039 (
            .O(N__37334),
            .I(N__37328));
    InMux I__7038 (
            .O(N__37333),
            .I(N__37325));
    Odrv12 I__7037 (
            .O(N__37328),
            .I(n3213));
    LocalMux I__7036 (
            .O(N__37325),
            .I(n3213));
    CascadeMux I__7035 (
            .O(N__37320),
            .I(N__37317));
    InMux I__7034 (
            .O(N__37317),
            .I(N__37314));
    LocalMux I__7033 (
            .O(N__37314),
            .I(n3280));
    InMux I__7032 (
            .O(N__37311),
            .I(n12942));
    CascadeMux I__7031 (
            .O(N__37308),
            .I(N__37304));
    InMux I__7030 (
            .O(N__37307),
            .I(N__37301));
    InMux I__7029 (
            .O(N__37304),
            .I(N__37298));
    LocalMux I__7028 (
            .O(N__37301),
            .I(N__37293));
    LocalMux I__7027 (
            .O(N__37298),
            .I(N__37293));
    Odrv4 I__7026 (
            .O(N__37293),
            .I(n3212));
    InMux I__7025 (
            .O(N__37290),
            .I(N__37287));
    LocalMux I__7024 (
            .O(N__37287),
            .I(n3279));
    InMux I__7023 (
            .O(N__37284),
            .I(n12943));
    InMux I__7022 (
            .O(N__37281),
            .I(N__37278));
    LocalMux I__7021 (
            .O(N__37278),
            .I(N__37274));
    InMux I__7020 (
            .O(N__37277),
            .I(N__37270));
    Span4Mux_s2_v I__7019 (
            .O(N__37274),
            .I(N__37267));
    InMux I__7018 (
            .O(N__37273),
            .I(N__37264));
    LocalMux I__7017 (
            .O(N__37270),
            .I(n3211));
    Odrv4 I__7016 (
            .O(N__37267),
            .I(n3211));
    LocalMux I__7015 (
            .O(N__37264),
            .I(n3211));
    InMux I__7014 (
            .O(N__37257),
            .I(N__37254));
    LocalMux I__7013 (
            .O(N__37254),
            .I(n3278));
    InMux I__7012 (
            .O(N__37251),
            .I(bfn_7_32_0_));
    InMux I__7011 (
            .O(N__37248),
            .I(N__37243));
    InMux I__7010 (
            .O(N__37247),
            .I(N__37240));
    InMux I__7009 (
            .O(N__37246),
            .I(N__37237));
    LocalMux I__7008 (
            .O(N__37243),
            .I(N__37234));
    LocalMux I__7007 (
            .O(N__37240),
            .I(N__37231));
    LocalMux I__7006 (
            .O(N__37237),
            .I(n3210));
    Odrv4 I__7005 (
            .O(N__37234),
            .I(n3210));
    Odrv4 I__7004 (
            .O(N__37231),
            .I(n3210));
    InMux I__7003 (
            .O(N__37224),
            .I(N__37221));
    LocalMux I__7002 (
            .O(N__37221),
            .I(N__37218));
    Odrv4 I__7001 (
            .O(N__37218),
            .I(n3277));
    InMux I__7000 (
            .O(N__37215),
            .I(n12945));
    CascadeMux I__6999 (
            .O(N__37212),
            .I(N__37208));
    CascadeMux I__6998 (
            .O(N__37211),
            .I(N__37204));
    InMux I__6997 (
            .O(N__37208),
            .I(N__37201));
    InMux I__6996 (
            .O(N__37207),
            .I(N__37198));
    InMux I__6995 (
            .O(N__37204),
            .I(N__37195));
    LocalMux I__6994 (
            .O(N__37201),
            .I(N__37192));
    LocalMux I__6993 (
            .O(N__37198),
            .I(n3225));
    LocalMux I__6992 (
            .O(N__37195),
            .I(n3225));
    Odrv4 I__6991 (
            .O(N__37192),
            .I(n3225));
    InMux I__6990 (
            .O(N__37185),
            .I(N__37182));
    LocalMux I__6989 (
            .O(N__37182),
            .I(n3292));
    InMux I__6988 (
            .O(N__37179),
            .I(n12930));
    CascadeMux I__6987 (
            .O(N__37176),
            .I(N__37173));
    InMux I__6986 (
            .O(N__37173),
            .I(N__37169));
    CascadeMux I__6985 (
            .O(N__37172),
            .I(N__37166));
    LocalMux I__6984 (
            .O(N__37169),
            .I(N__37162));
    InMux I__6983 (
            .O(N__37166),
            .I(N__37157));
    InMux I__6982 (
            .O(N__37165),
            .I(N__37157));
    Odrv4 I__6981 (
            .O(N__37162),
            .I(n3224));
    LocalMux I__6980 (
            .O(N__37157),
            .I(n3224));
    InMux I__6979 (
            .O(N__37152),
            .I(N__37149));
    LocalMux I__6978 (
            .O(N__37149),
            .I(N__37146));
    Odrv4 I__6977 (
            .O(N__37146),
            .I(n3291));
    InMux I__6976 (
            .O(N__37143),
            .I(n12931));
    CascadeMux I__6975 (
            .O(N__37140),
            .I(N__37136));
    InMux I__6974 (
            .O(N__37139),
            .I(N__37133));
    InMux I__6973 (
            .O(N__37136),
            .I(N__37130));
    LocalMux I__6972 (
            .O(N__37133),
            .I(N__37126));
    LocalMux I__6971 (
            .O(N__37130),
            .I(N__37123));
    InMux I__6970 (
            .O(N__37129),
            .I(N__37120));
    Odrv4 I__6969 (
            .O(N__37126),
            .I(n3223));
    Odrv4 I__6968 (
            .O(N__37123),
            .I(n3223));
    LocalMux I__6967 (
            .O(N__37120),
            .I(n3223));
    InMux I__6966 (
            .O(N__37113),
            .I(N__37110));
    LocalMux I__6965 (
            .O(N__37110),
            .I(N__37107));
    Span4Mux_s2_v I__6964 (
            .O(N__37107),
            .I(N__37104));
    Odrv4 I__6963 (
            .O(N__37104),
            .I(n3290));
    InMux I__6962 (
            .O(N__37101),
            .I(n12932));
    CascadeMux I__6961 (
            .O(N__37098),
            .I(N__37095));
    InMux I__6960 (
            .O(N__37095),
            .I(N__37091));
    InMux I__6959 (
            .O(N__37094),
            .I(N__37087));
    LocalMux I__6958 (
            .O(N__37091),
            .I(N__37084));
    InMux I__6957 (
            .O(N__37090),
            .I(N__37081));
    LocalMux I__6956 (
            .O(N__37087),
            .I(n3222));
    Odrv4 I__6955 (
            .O(N__37084),
            .I(n3222));
    LocalMux I__6954 (
            .O(N__37081),
            .I(n3222));
    InMux I__6953 (
            .O(N__37074),
            .I(N__37071));
    LocalMux I__6952 (
            .O(N__37071),
            .I(N__37068));
    Span4Mux_s2_v I__6951 (
            .O(N__37068),
            .I(N__37065));
    Odrv4 I__6950 (
            .O(N__37065),
            .I(n3289));
    InMux I__6949 (
            .O(N__37062),
            .I(n12933));
    CascadeMux I__6948 (
            .O(N__37059),
            .I(N__37055));
    CascadeMux I__6947 (
            .O(N__37058),
            .I(N__37052));
    InMux I__6946 (
            .O(N__37055),
            .I(N__37049));
    InMux I__6945 (
            .O(N__37052),
            .I(N__37045));
    LocalMux I__6944 (
            .O(N__37049),
            .I(N__37042));
    InMux I__6943 (
            .O(N__37048),
            .I(N__37039));
    LocalMux I__6942 (
            .O(N__37045),
            .I(n3221));
    Odrv4 I__6941 (
            .O(N__37042),
            .I(n3221));
    LocalMux I__6940 (
            .O(N__37039),
            .I(n3221));
    InMux I__6939 (
            .O(N__37032),
            .I(N__37029));
    LocalMux I__6938 (
            .O(N__37029),
            .I(n3288));
    InMux I__6937 (
            .O(N__37026),
            .I(n12934));
    CascadeMux I__6936 (
            .O(N__37023),
            .I(N__37020));
    InMux I__6935 (
            .O(N__37020),
            .I(N__37016));
    InMux I__6934 (
            .O(N__37019),
            .I(N__37012));
    LocalMux I__6933 (
            .O(N__37016),
            .I(N__37009));
    InMux I__6932 (
            .O(N__37015),
            .I(N__37006));
    LocalMux I__6931 (
            .O(N__37012),
            .I(n3220));
    Odrv4 I__6930 (
            .O(N__37009),
            .I(n3220));
    LocalMux I__6929 (
            .O(N__37006),
            .I(n3220));
    InMux I__6928 (
            .O(N__36999),
            .I(N__36996));
    LocalMux I__6927 (
            .O(N__36996),
            .I(N__36993));
    Odrv12 I__6926 (
            .O(N__36993),
            .I(n3287));
    InMux I__6925 (
            .O(N__36990),
            .I(n12935));
    CascadeMux I__6924 (
            .O(N__36987),
            .I(N__36983));
    InMux I__6923 (
            .O(N__36986),
            .I(N__36980));
    InMux I__6922 (
            .O(N__36983),
            .I(N__36977));
    LocalMux I__6921 (
            .O(N__36980),
            .I(N__36973));
    LocalMux I__6920 (
            .O(N__36977),
            .I(N__36970));
    InMux I__6919 (
            .O(N__36976),
            .I(N__36967));
    Span4Mux_s1_v I__6918 (
            .O(N__36973),
            .I(N__36960));
    Span4Mux_h I__6917 (
            .O(N__36970),
            .I(N__36960));
    LocalMux I__6916 (
            .O(N__36967),
            .I(N__36960));
    Span4Mux_h I__6915 (
            .O(N__36960),
            .I(N__36957));
    Odrv4 I__6914 (
            .O(N__36957),
            .I(n3219));
    CascadeMux I__6913 (
            .O(N__36954),
            .I(N__36951));
    InMux I__6912 (
            .O(N__36951),
            .I(N__36948));
    LocalMux I__6911 (
            .O(N__36948),
            .I(N__36945));
    Span4Mux_s1_v I__6910 (
            .O(N__36945),
            .I(N__36942));
    Odrv4 I__6909 (
            .O(N__36942),
            .I(n3286));
    InMux I__6908 (
            .O(N__36939),
            .I(bfn_7_31_0_));
    CascadeMux I__6907 (
            .O(N__36936),
            .I(N__36933));
    InMux I__6906 (
            .O(N__36933),
            .I(N__36929));
    InMux I__6905 (
            .O(N__36932),
            .I(N__36926));
    LocalMux I__6904 (
            .O(N__36929),
            .I(N__36923));
    LocalMux I__6903 (
            .O(N__36926),
            .I(n3218));
    Odrv4 I__6902 (
            .O(N__36923),
            .I(n3218));
    CascadeMux I__6901 (
            .O(N__36918),
            .I(N__36915));
    InMux I__6900 (
            .O(N__36915),
            .I(N__36912));
    LocalMux I__6899 (
            .O(N__36912),
            .I(N__36909));
    Odrv4 I__6898 (
            .O(N__36909),
            .I(n3285));
    InMux I__6897 (
            .O(N__36906),
            .I(n12937));
    CascadeMux I__6896 (
            .O(N__36903),
            .I(N__36900));
    InMux I__6895 (
            .O(N__36900),
            .I(N__36896));
    InMux I__6894 (
            .O(N__36899),
            .I(N__36892));
    LocalMux I__6893 (
            .O(N__36896),
            .I(N__36889));
    InMux I__6892 (
            .O(N__36895),
            .I(N__36886));
    LocalMux I__6891 (
            .O(N__36892),
            .I(n3232));
    Odrv4 I__6890 (
            .O(N__36889),
            .I(n3232));
    LocalMux I__6889 (
            .O(N__36886),
            .I(n3232));
    InMux I__6888 (
            .O(N__36879),
            .I(N__36876));
    LocalMux I__6887 (
            .O(N__36876),
            .I(n3299));
    InMux I__6886 (
            .O(N__36873),
            .I(n12923));
    CascadeMux I__6885 (
            .O(N__36870),
            .I(N__36867));
    InMux I__6884 (
            .O(N__36867),
            .I(N__36862));
    InMux I__6883 (
            .O(N__36866),
            .I(N__36859));
    InMux I__6882 (
            .O(N__36865),
            .I(N__36856));
    LocalMux I__6881 (
            .O(N__36862),
            .I(N__36853));
    LocalMux I__6880 (
            .O(N__36859),
            .I(n3231));
    LocalMux I__6879 (
            .O(N__36856),
            .I(n3231));
    Odrv4 I__6878 (
            .O(N__36853),
            .I(n3231));
    InMux I__6877 (
            .O(N__36846),
            .I(n12924));
    InMux I__6876 (
            .O(N__36843),
            .I(N__36840));
    LocalMux I__6875 (
            .O(N__36840),
            .I(n3298));
    CascadeMux I__6874 (
            .O(N__36837),
            .I(N__36834));
    InMux I__6873 (
            .O(N__36834),
            .I(N__36829));
    InMux I__6872 (
            .O(N__36833),
            .I(N__36826));
    InMux I__6871 (
            .O(N__36832),
            .I(N__36823));
    LocalMux I__6870 (
            .O(N__36829),
            .I(N__36820));
    LocalMux I__6869 (
            .O(N__36826),
            .I(n3230));
    LocalMux I__6868 (
            .O(N__36823),
            .I(n3230));
    Odrv4 I__6867 (
            .O(N__36820),
            .I(n3230));
    InMux I__6866 (
            .O(N__36813),
            .I(N__36810));
    LocalMux I__6865 (
            .O(N__36810),
            .I(N__36807));
    Odrv4 I__6864 (
            .O(N__36807),
            .I(n15079));
    InMux I__6863 (
            .O(N__36804),
            .I(n12925));
    InMux I__6862 (
            .O(N__36801),
            .I(N__36797));
    CascadeMux I__6861 (
            .O(N__36800),
            .I(N__36794));
    LocalMux I__6860 (
            .O(N__36797),
            .I(N__36790));
    InMux I__6859 (
            .O(N__36794),
            .I(N__36787));
    InMux I__6858 (
            .O(N__36793),
            .I(N__36784));
    Span4Mux_h I__6857 (
            .O(N__36790),
            .I(N__36779));
    LocalMux I__6856 (
            .O(N__36787),
            .I(N__36779));
    LocalMux I__6855 (
            .O(N__36784),
            .I(n3229));
    Odrv4 I__6854 (
            .O(N__36779),
            .I(n3229));
    InMux I__6853 (
            .O(N__36774),
            .I(N__36771));
    LocalMux I__6852 (
            .O(N__36771),
            .I(N__36768));
    Span4Mux_s3_v I__6851 (
            .O(N__36768),
            .I(N__36765));
    Odrv4 I__6850 (
            .O(N__36765),
            .I(n3296));
    InMux I__6849 (
            .O(N__36762),
            .I(n12926));
    CascadeMux I__6848 (
            .O(N__36759),
            .I(N__36755));
    InMux I__6847 (
            .O(N__36758),
            .I(N__36752));
    InMux I__6846 (
            .O(N__36755),
            .I(N__36749));
    LocalMux I__6845 (
            .O(N__36752),
            .I(N__36746));
    LocalMux I__6844 (
            .O(N__36749),
            .I(N__36743));
    Odrv4 I__6843 (
            .O(N__36746),
            .I(n3228));
    Odrv4 I__6842 (
            .O(N__36743),
            .I(n3228));
    InMux I__6841 (
            .O(N__36738),
            .I(N__36735));
    LocalMux I__6840 (
            .O(N__36735),
            .I(N__36732));
    Span4Mux_h I__6839 (
            .O(N__36732),
            .I(N__36729));
    Odrv4 I__6838 (
            .O(N__36729),
            .I(n3295));
    InMux I__6837 (
            .O(N__36726),
            .I(n12927));
    CascadeMux I__6836 (
            .O(N__36723),
            .I(N__36720));
    InMux I__6835 (
            .O(N__36720),
            .I(N__36717));
    LocalMux I__6834 (
            .O(N__36717),
            .I(N__36713));
    InMux I__6833 (
            .O(N__36716),
            .I(N__36709));
    Span4Mux_h I__6832 (
            .O(N__36713),
            .I(N__36706));
    InMux I__6831 (
            .O(N__36712),
            .I(N__36703));
    LocalMux I__6830 (
            .O(N__36709),
            .I(n3227));
    Odrv4 I__6829 (
            .O(N__36706),
            .I(n3227));
    LocalMux I__6828 (
            .O(N__36703),
            .I(n3227));
    InMux I__6827 (
            .O(N__36696),
            .I(N__36693));
    LocalMux I__6826 (
            .O(N__36693),
            .I(N__36690));
    Span4Mux_s2_v I__6825 (
            .O(N__36690),
            .I(N__36687));
    Odrv4 I__6824 (
            .O(N__36687),
            .I(n3294));
    InMux I__6823 (
            .O(N__36684),
            .I(bfn_7_30_0_));
    CascadeMux I__6822 (
            .O(N__36681),
            .I(N__36678));
    InMux I__6821 (
            .O(N__36678),
            .I(N__36674));
    InMux I__6820 (
            .O(N__36677),
            .I(N__36671));
    LocalMux I__6819 (
            .O(N__36674),
            .I(N__36668));
    LocalMux I__6818 (
            .O(N__36671),
            .I(n3226));
    Odrv12 I__6817 (
            .O(N__36668),
            .I(n3226));
    InMux I__6816 (
            .O(N__36663),
            .I(N__36660));
    LocalMux I__6815 (
            .O(N__36660),
            .I(N__36657));
    Odrv12 I__6814 (
            .O(N__36657),
            .I(n3293));
    InMux I__6813 (
            .O(N__36654),
            .I(n12929));
    InMux I__6812 (
            .O(N__36651),
            .I(n12974));
    CascadeMux I__6811 (
            .O(N__36648),
            .I(N__36645));
    InMux I__6810 (
            .O(N__36645),
            .I(N__36642));
    LocalMux I__6809 (
            .O(N__36642),
            .I(N__36638));
    InMux I__6808 (
            .O(N__36641),
            .I(N__36635));
    Span4Mux_v I__6807 (
            .O(N__36638),
            .I(N__36632));
    LocalMux I__6806 (
            .O(N__36635),
            .I(n12051));
    Odrv4 I__6805 (
            .O(N__36632),
            .I(n12051));
    InMux I__6804 (
            .O(N__36627),
            .I(N__36624));
    LocalMux I__6803 (
            .O(N__36624),
            .I(N__36621));
    Odrv4 I__6802 (
            .O(N__36621),
            .I(n15490));
    InMux I__6801 (
            .O(N__36618),
            .I(N__36614));
    InMux I__6800 (
            .O(N__36617),
            .I(N__36611));
    LocalMux I__6799 (
            .O(N__36614),
            .I(N__36608));
    LocalMux I__6798 (
            .O(N__36611),
            .I(N__36605));
    Sp12to4 I__6797 (
            .O(N__36608),
            .I(N__36602));
    Span4Mux_v I__6796 (
            .O(N__36605),
            .I(N__36599));
    Odrv12 I__6795 (
            .O(N__36602),
            .I(n319));
    Odrv4 I__6794 (
            .O(N__36599),
            .I(n319));
    InMux I__6793 (
            .O(N__36594),
            .I(N__36589));
    InMux I__6792 (
            .O(N__36593),
            .I(N__36586));
    InMux I__6791 (
            .O(N__36592),
            .I(N__36583));
    LocalMux I__6790 (
            .O(N__36589),
            .I(N__36576));
    LocalMux I__6789 (
            .O(N__36586),
            .I(N__36576));
    LocalMux I__6788 (
            .O(N__36583),
            .I(N__36576));
    Span4Mux_v I__6787 (
            .O(N__36576),
            .I(N__36573));
    Odrv4 I__6786 (
            .O(N__36573),
            .I(n318));
    CascadeMux I__6785 (
            .O(N__36570),
            .I(N__36567));
    InMux I__6784 (
            .O(N__36567),
            .I(N__36564));
    LocalMux I__6783 (
            .O(N__36564),
            .I(n3301));
    InMux I__6782 (
            .O(N__36561),
            .I(n12921));
    CascadeMux I__6781 (
            .O(N__36558),
            .I(N__36554));
    CascadeMux I__6780 (
            .O(N__36557),
            .I(N__36551));
    InMux I__6779 (
            .O(N__36554),
            .I(N__36548));
    InMux I__6778 (
            .O(N__36551),
            .I(N__36545));
    LocalMux I__6777 (
            .O(N__36548),
            .I(n3233));
    LocalMux I__6776 (
            .O(N__36545),
            .I(n3233));
    InMux I__6775 (
            .O(N__36540),
            .I(N__36537));
    LocalMux I__6774 (
            .O(N__36537),
            .I(n3300));
    InMux I__6773 (
            .O(N__36534),
            .I(n12922));
    InMux I__6772 (
            .O(N__36531),
            .I(n12965));
    InMux I__6771 (
            .O(N__36528),
            .I(N__36525));
    LocalMux I__6770 (
            .O(N__36525),
            .I(N__36522));
    Span4Mux_v I__6769 (
            .O(N__36522),
            .I(N__36519));
    Odrv4 I__6768 (
            .O(N__36519),
            .I(n15652));
    InMux I__6767 (
            .O(N__36516),
            .I(n12966));
    InMux I__6766 (
            .O(N__36513),
            .I(bfn_7_27_0_));
    InMux I__6765 (
            .O(N__36510),
            .I(n12968));
    InMux I__6764 (
            .O(N__36507),
            .I(n12969));
    InMux I__6763 (
            .O(N__36504),
            .I(n12970));
    InMux I__6762 (
            .O(N__36501),
            .I(n12971));
    InMux I__6761 (
            .O(N__36498),
            .I(n12972));
    InMux I__6760 (
            .O(N__36495),
            .I(n12973));
    InMux I__6759 (
            .O(N__36492),
            .I(N__36488));
    CascadeMux I__6758 (
            .O(N__36491),
            .I(N__36485));
    LocalMux I__6757 (
            .O(N__36488),
            .I(N__36482));
    InMux I__6756 (
            .O(N__36485),
            .I(N__36479));
    Span4Mux_v I__6755 (
            .O(N__36482),
            .I(N__36476));
    LocalMux I__6754 (
            .O(N__36479),
            .I(N__36473));
    Span4Mux_h I__6753 (
            .O(N__36476),
            .I(N__36468));
    Span4Mux_s2_h I__6752 (
            .O(N__36473),
            .I(N__36468));
    Odrv4 I__6751 (
            .O(N__36468),
            .I(n15322));
    InMux I__6750 (
            .O(N__36465),
            .I(N__36462));
    LocalMux I__6749 (
            .O(N__36462),
            .I(N__36459));
    Span4Mux_v I__6748 (
            .O(N__36459),
            .I(N__36450));
    InMux I__6747 (
            .O(N__36458),
            .I(N__36447));
    CascadeMux I__6746 (
            .O(N__36457),
            .I(N__36442));
    CascadeMux I__6745 (
            .O(N__36456),
            .I(N__36439));
    CascadeMux I__6744 (
            .O(N__36455),
            .I(N__36434));
    CascadeMux I__6743 (
            .O(N__36454),
            .I(N__36431));
    CascadeMux I__6742 (
            .O(N__36453),
            .I(N__36419));
    Span4Mux_h I__6741 (
            .O(N__36450),
            .I(N__36412));
    LocalMux I__6740 (
            .O(N__36447),
            .I(N__36412));
    CascadeMux I__6739 (
            .O(N__36446),
            .I(N__36405));
    CascadeMux I__6738 (
            .O(N__36445),
            .I(N__36402));
    InMux I__6737 (
            .O(N__36442),
            .I(N__36393));
    InMux I__6736 (
            .O(N__36439),
            .I(N__36393));
    InMux I__6735 (
            .O(N__36438),
            .I(N__36393));
    InMux I__6734 (
            .O(N__36437),
            .I(N__36393));
    InMux I__6733 (
            .O(N__36434),
            .I(N__36380));
    InMux I__6732 (
            .O(N__36431),
            .I(N__36380));
    InMux I__6731 (
            .O(N__36430),
            .I(N__36380));
    InMux I__6730 (
            .O(N__36429),
            .I(N__36380));
    InMux I__6729 (
            .O(N__36428),
            .I(N__36380));
    InMux I__6728 (
            .O(N__36427),
            .I(N__36380));
    InMux I__6727 (
            .O(N__36426),
            .I(N__36375));
    InMux I__6726 (
            .O(N__36425),
            .I(N__36375));
    InMux I__6725 (
            .O(N__36424),
            .I(N__36370));
    InMux I__6724 (
            .O(N__36423),
            .I(N__36370));
    InMux I__6723 (
            .O(N__36422),
            .I(N__36363));
    InMux I__6722 (
            .O(N__36419),
            .I(N__36363));
    InMux I__6721 (
            .O(N__36418),
            .I(N__36363));
    InMux I__6720 (
            .O(N__36417),
            .I(N__36360));
    Span4Mux_v I__6719 (
            .O(N__36412),
            .I(N__36357));
    InMux I__6718 (
            .O(N__36411),
            .I(N__36354));
    InMux I__6717 (
            .O(N__36410),
            .I(N__36349));
    InMux I__6716 (
            .O(N__36409),
            .I(N__36349));
    InMux I__6715 (
            .O(N__36408),
            .I(N__36342));
    InMux I__6714 (
            .O(N__36405),
            .I(N__36342));
    InMux I__6713 (
            .O(N__36402),
            .I(N__36342));
    LocalMux I__6712 (
            .O(N__36393),
            .I(N__36335));
    LocalMux I__6711 (
            .O(N__36380),
            .I(N__36335));
    LocalMux I__6710 (
            .O(N__36375),
            .I(N__36335));
    LocalMux I__6709 (
            .O(N__36370),
            .I(N__36330));
    LocalMux I__6708 (
            .O(N__36363),
            .I(N__36330));
    LocalMux I__6707 (
            .O(N__36360),
            .I(N__36327));
    Odrv4 I__6706 (
            .O(N__36357),
            .I(n2742));
    LocalMux I__6705 (
            .O(N__36354),
            .I(n2742));
    LocalMux I__6704 (
            .O(N__36349),
            .I(n2742));
    LocalMux I__6703 (
            .O(N__36342),
            .I(n2742));
    Odrv4 I__6702 (
            .O(N__36335),
            .I(n2742));
    Odrv4 I__6701 (
            .O(N__36330),
            .I(n2742));
    Odrv4 I__6700 (
            .O(N__36327),
            .I(n2742));
    InMux I__6699 (
            .O(N__36312),
            .I(n12957));
    InMux I__6698 (
            .O(N__36309),
            .I(N__36306));
    LocalMux I__6697 (
            .O(N__36306),
            .I(N__36303));
    Span4Mux_h I__6696 (
            .O(N__36303),
            .I(N__36300));
    Odrv4 I__6695 (
            .O(N__36300),
            .I(n15292));
    InMux I__6694 (
            .O(N__36297),
            .I(N__36289));
    InMux I__6693 (
            .O(N__36296),
            .I(N__36286));
    InMux I__6692 (
            .O(N__36295),
            .I(N__36283));
    CascadeMux I__6691 (
            .O(N__36294),
            .I(N__36272));
    CascadeMux I__6690 (
            .O(N__36293),
            .I(N__36269));
    CascadeMux I__6689 (
            .O(N__36292),
            .I(N__36263));
    LocalMux I__6688 (
            .O(N__36289),
            .I(N__36259));
    LocalMux I__6687 (
            .O(N__36286),
            .I(N__36255));
    LocalMux I__6686 (
            .O(N__36283),
            .I(N__36252));
    CascadeMux I__6685 (
            .O(N__36282),
            .I(N__36249));
    CascadeMux I__6684 (
            .O(N__36281),
            .I(N__36246));
    CascadeMux I__6683 (
            .O(N__36280),
            .I(N__36242));
    CascadeMux I__6682 (
            .O(N__36279),
            .I(N__36236));
    CascadeMux I__6681 (
            .O(N__36278),
            .I(N__36231));
    CascadeMux I__6680 (
            .O(N__36277),
            .I(N__36228));
    CascadeMux I__6679 (
            .O(N__36276),
            .I(N__36225));
    InMux I__6678 (
            .O(N__36275),
            .I(N__36217));
    InMux I__6677 (
            .O(N__36272),
            .I(N__36217));
    InMux I__6676 (
            .O(N__36269),
            .I(N__36217));
    InMux I__6675 (
            .O(N__36268),
            .I(N__36212));
    InMux I__6674 (
            .O(N__36267),
            .I(N__36212));
    InMux I__6673 (
            .O(N__36266),
            .I(N__36205));
    InMux I__6672 (
            .O(N__36263),
            .I(N__36205));
    InMux I__6671 (
            .O(N__36262),
            .I(N__36205));
    Span12Mux_s9_v I__6670 (
            .O(N__36259),
            .I(N__36202));
    InMux I__6669 (
            .O(N__36258),
            .I(N__36199));
    Span4Mux_h I__6668 (
            .O(N__36255),
            .I(N__36194));
    Span4Mux_s3_h I__6667 (
            .O(N__36252),
            .I(N__36194));
    InMux I__6666 (
            .O(N__36249),
            .I(N__36189));
    InMux I__6665 (
            .O(N__36246),
            .I(N__36189));
    InMux I__6664 (
            .O(N__36245),
            .I(N__36184));
    InMux I__6663 (
            .O(N__36242),
            .I(N__36184));
    InMux I__6662 (
            .O(N__36241),
            .I(N__36179));
    InMux I__6661 (
            .O(N__36240),
            .I(N__36179));
    InMux I__6660 (
            .O(N__36239),
            .I(N__36170));
    InMux I__6659 (
            .O(N__36236),
            .I(N__36170));
    InMux I__6658 (
            .O(N__36235),
            .I(N__36170));
    InMux I__6657 (
            .O(N__36234),
            .I(N__36170));
    InMux I__6656 (
            .O(N__36231),
            .I(N__36161));
    InMux I__6655 (
            .O(N__36228),
            .I(N__36161));
    InMux I__6654 (
            .O(N__36225),
            .I(N__36161));
    InMux I__6653 (
            .O(N__36224),
            .I(N__36161));
    LocalMux I__6652 (
            .O(N__36217),
            .I(N__36154));
    LocalMux I__6651 (
            .O(N__36212),
            .I(N__36154));
    LocalMux I__6650 (
            .O(N__36205),
            .I(N__36154));
    Odrv12 I__6649 (
            .O(N__36202),
            .I(n2643));
    LocalMux I__6648 (
            .O(N__36199),
            .I(n2643));
    Odrv4 I__6647 (
            .O(N__36194),
            .I(n2643));
    LocalMux I__6646 (
            .O(N__36189),
            .I(n2643));
    LocalMux I__6645 (
            .O(N__36184),
            .I(n2643));
    LocalMux I__6644 (
            .O(N__36179),
            .I(n2643));
    LocalMux I__6643 (
            .O(N__36170),
            .I(n2643));
    LocalMux I__6642 (
            .O(N__36161),
            .I(n2643));
    Odrv4 I__6641 (
            .O(N__36154),
            .I(n2643));
    InMux I__6640 (
            .O(N__36135),
            .I(N__36132));
    LocalMux I__6639 (
            .O(N__36132),
            .I(N__36129));
    Span4Mux_h I__6638 (
            .O(N__36129),
            .I(N__36126));
    Odrv4 I__6637 (
            .O(N__36126),
            .I(encoder0_position_scaled_7));
    InMux I__6636 (
            .O(N__36123),
            .I(n12958));
    InMux I__6635 (
            .O(N__36120),
            .I(N__36117));
    LocalMux I__6634 (
            .O(N__36117),
            .I(N__36114));
    Span4Mux_h I__6633 (
            .O(N__36114),
            .I(N__36110));
    InMux I__6632 (
            .O(N__36113),
            .I(N__36107));
    Odrv4 I__6631 (
            .O(N__36110),
            .I(n15830));
    LocalMux I__6630 (
            .O(N__36107),
            .I(n15830));
    CascadeMux I__6629 (
            .O(N__36102),
            .I(N__36091));
    InMux I__6628 (
            .O(N__36101),
            .I(N__36087));
    CascadeMux I__6627 (
            .O(N__36100),
            .I(N__36082));
    InMux I__6626 (
            .O(N__36099),
            .I(N__36077));
    InMux I__6625 (
            .O(N__36098),
            .I(N__36077));
    InMux I__6624 (
            .O(N__36097),
            .I(N__36074));
    InMux I__6623 (
            .O(N__36096),
            .I(N__36071));
    InMux I__6622 (
            .O(N__36095),
            .I(N__36065));
    InMux I__6621 (
            .O(N__36094),
            .I(N__36058));
    InMux I__6620 (
            .O(N__36091),
            .I(N__36058));
    InMux I__6619 (
            .O(N__36090),
            .I(N__36058));
    LocalMux I__6618 (
            .O(N__36087),
            .I(N__36054));
    CascadeMux I__6617 (
            .O(N__36086),
            .I(N__36051));
    CascadeMux I__6616 (
            .O(N__36085),
            .I(N__36045));
    InMux I__6615 (
            .O(N__36082),
            .I(N__36041));
    LocalMux I__6614 (
            .O(N__36077),
            .I(N__36038));
    LocalMux I__6613 (
            .O(N__36074),
            .I(N__36035));
    LocalMux I__6612 (
            .O(N__36071),
            .I(N__36032));
    CascadeMux I__6611 (
            .O(N__36070),
            .I(N__36027));
    CascadeMux I__6610 (
            .O(N__36069),
            .I(N__36024));
    InMux I__6609 (
            .O(N__36068),
            .I(N__36020));
    LocalMux I__6608 (
            .O(N__36065),
            .I(N__36015));
    LocalMux I__6607 (
            .O(N__36058),
            .I(N__36015));
    InMux I__6606 (
            .O(N__36057),
            .I(N__36012));
    Span4Mux_v I__6605 (
            .O(N__36054),
            .I(N__36008));
    InMux I__6604 (
            .O(N__36051),
            .I(N__35995));
    InMux I__6603 (
            .O(N__36050),
            .I(N__35995));
    InMux I__6602 (
            .O(N__36049),
            .I(N__35995));
    InMux I__6601 (
            .O(N__36048),
            .I(N__35995));
    InMux I__6600 (
            .O(N__36045),
            .I(N__35995));
    InMux I__6599 (
            .O(N__36044),
            .I(N__35995));
    LocalMux I__6598 (
            .O(N__36041),
            .I(N__35986));
    Span4Mux_h I__6597 (
            .O(N__36038),
            .I(N__35986));
    Span4Mux_v I__6596 (
            .O(N__36035),
            .I(N__35986));
    Span4Mux_h I__6595 (
            .O(N__36032),
            .I(N__35986));
    InMux I__6594 (
            .O(N__36031),
            .I(N__35975));
    InMux I__6593 (
            .O(N__36030),
            .I(N__35975));
    InMux I__6592 (
            .O(N__36027),
            .I(N__35975));
    InMux I__6591 (
            .O(N__36024),
            .I(N__35975));
    InMux I__6590 (
            .O(N__36023),
            .I(N__35975));
    LocalMux I__6589 (
            .O(N__36020),
            .I(N__35968));
    Span4Mux_h I__6588 (
            .O(N__36015),
            .I(N__35968));
    LocalMux I__6587 (
            .O(N__36012),
            .I(N__35968));
    InMux I__6586 (
            .O(N__36011),
            .I(N__35965));
    Odrv4 I__6585 (
            .O(N__36008),
            .I(n2544));
    LocalMux I__6584 (
            .O(N__35995),
            .I(n2544));
    Odrv4 I__6583 (
            .O(N__35986),
            .I(n2544));
    LocalMux I__6582 (
            .O(N__35975),
            .I(n2544));
    Odrv4 I__6581 (
            .O(N__35968),
            .I(n2544));
    LocalMux I__6580 (
            .O(N__35965),
            .I(n2544));
    InMux I__6579 (
            .O(N__35952),
            .I(bfn_7_26_0_));
    InMux I__6578 (
            .O(N__35949),
            .I(N__35945));
    CascadeMux I__6577 (
            .O(N__35948),
            .I(N__35942));
    LocalMux I__6576 (
            .O(N__35945),
            .I(N__35939));
    InMux I__6575 (
            .O(N__35942),
            .I(N__35936));
    Span4Mux_v I__6574 (
            .O(N__35939),
            .I(N__35933));
    LocalMux I__6573 (
            .O(N__35936),
            .I(N__35930));
    Span4Mux_v I__6572 (
            .O(N__35933),
            .I(N__35927));
    Span4Mux_v I__6571 (
            .O(N__35930),
            .I(N__35924));
    Span4Mux_h I__6570 (
            .O(N__35927),
            .I(N__35921));
    Span4Mux_h I__6569 (
            .O(N__35924),
            .I(N__35918));
    Odrv4 I__6568 (
            .O(N__35921),
            .I(n15802));
    Odrv4 I__6567 (
            .O(N__35918),
            .I(n15802));
    InMux I__6566 (
            .O(N__35913),
            .I(N__35908));
    CascadeMux I__6565 (
            .O(N__35912),
            .I(N__35905));
    InMux I__6564 (
            .O(N__35911),
            .I(N__35893));
    LocalMux I__6563 (
            .O(N__35908),
            .I(N__35890));
    InMux I__6562 (
            .O(N__35905),
            .I(N__35881));
    InMux I__6561 (
            .O(N__35904),
            .I(N__35881));
    InMux I__6560 (
            .O(N__35903),
            .I(N__35881));
    InMux I__6559 (
            .O(N__35902),
            .I(N__35881));
    InMux I__6558 (
            .O(N__35901),
            .I(N__35878));
    InMux I__6557 (
            .O(N__35900),
            .I(N__35875));
    CascadeMux I__6556 (
            .O(N__35899),
            .I(N__35871));
    CascadeMux I__6555 (
            .O(N__35898),
            .I(N__35863));
    CascadeMux I__6554 (
            .O(N__35897),
            .I(N__35857));
    InMux I__6553 (
            .O(N__35896),
            .I(N__35852));
    LocalMux I__6552 (
            .O(N__35893),
            .I(N__35847));
    Span4Mux_h I__6551 (
            .O(N__35890),
            .I(N__35847));
    LocalMux I__6550 (
            .O(N__35881),
            .I(N__35844));
    LocalMux I__6549 (
            .O(N__35878),
            .I(N__35839));
    LocalMux I__6548 (
            .O(N__35875),
            .I(N__35839));
    InMux I__6547 (
            .O(N__35874),
            .I(N__35832));
    InMux I__6546 (
            .O(N__35871),
            .I(N__35832));
    InMux I__6545 (
            .O(N__35870),
            .I(N__35832));
    InMux I__6544 (
            .O(N__35869),
            .I(N__35829));
    InMux I__6543 (
            .O(N__35868),
            .I(N__35822));
    InMux I__6542 (
            .O(N__35867),
            .I(N__35822));
    InMux I__6541 (
            .O(N__35866),
            .I(N__35822));
    InMux I__6540 (
            .O(N__35863),
            .I(N__35813));
    InMux I__6539 (
            .O(N__35862),
            .I(N__35813));
    InMux I__6538 (
            .O(N__35861),
            .I(N__35813));
    InMux I__6537 (
            .O(N__35860),
            .I(N__35813));
    InMux I__6536 (
            .O(N__35857),
            .I(N__35806));
    InMux I__6535 (
            .O(N__35856),
            .I(N__35806));
    InMux I__6534 (
            .O(N__35855),
            .I(N__35806));
    LocalMux I__6533 (
            .O(N__35852),
            .I(N__35801));
    Span4Mux_v I__6532 (
            .O(N__35847),
            .I(N__35801));
    Span4Mux_h I__6531 (
            .O(N__35844),
            .I(N__35796));
    Span4Mux_v I__6530 (
            .O(N__35839),
            .I(N__35796));
    LocalMux I__6529 (
            .O(N__35832),
            .I(n2445));
    LocalMux I__6528 (
            .O(N__35829),
            .I(n2445));
    LocalMux I__6527 (
            .O(N__35822),
            .I(n2445));
    LocalMux I__6526 (
            .O(N__35813),
            .I(n2445));
    LocalMux I__6525 (
            .O(N__35806),
            .I(n2445));
    Odrv4 I__6524 (
            .O(N__35801),
            .I(n2445));
    Odrv4 I__6523 (
            .O(N__35796),
            .I(n2445));
    InMux I__6522 (
            .O(N__35781),
            .I(n12960));
    InMux I__6521 (
            .O(N__35778),
            .I(N__35775));
    LocalMux I__6520 (
            .O(N__35775),
            .I(N__35772));
    Span4Mux_v I__6519 (
            .O(N__35772),
            .I(N__35769));
    Span4Mux_h I__6518 (
            .O(N__35769),
            .I(N__35766));
    Span4Mux_v I__6517 (
            .O(N__35766),
            .I(N__35762));
    InMux I__6516 (
            .O(N__35765),
            .I(N__35759));
    Odrv4 I__6515 (
            .O(N__35762),
            .I(n15775));
    LocalMux I__6514 (
            .O(N__35759),
            .I(n15775));
    InMux I__6513 (
            .O(N__35754),
            .I(N__35751));
    LocalMux I__6512 (
            .O(N__35751),
            .I(N__35748));
    Span4Mux_h I__6511 (
            .O(N__35748),
            .I(N__35735));
    InMux I__6510 (
            .O(N__35747),
            .I(N__35730));
    InMux I__6509 (
            .O(N__35746),
            .I(N__35730));
    CascadeMux I__6508 (
            .O(N__35745),
            .I(N__35727));
    InMux I__6507 (
            .O(N__35744),
            .I(N__35724));
    CascadeMux I__6506 (
            .O(N__35743),
            .I(N__35719));
    CascadeMux I__6505 (
            .O(N__35742),
            .I(N__35713));
    CascadeMux I__6504 (
            .O(N__35741),
            .I(N__35710));
    CascadeMux I__6503 (
            .O(N__35740),
            .I(N__35705));
    CascadeMux I__6502 (
            .O(N__35739),
            .I(N__35699));
    CascadeMux I__6501 (
            .O(N__35738),
            .I(N__35696));
    Span4Mux_v I__6500 (
            .O(N__35735),
            .I(N__35690));
    LocalMux I__6499 (
            .O(N__35730),
            .I(N__35690));
    InMux I__6498 (
            .O(N__35727),
            .I(N__35687));
    LocalMux I__6497 (
            .O(N__35724),
            .I(N__35684));
    InMux I__6496 (
            .O(N__35723),
            .I(N__35675));
    InMux I__6495 (
            .O(N__35722),
            .I(N__35675));
    InMux I__6494 (
            .O(N__35719),
            .I(N__35675));
    InMux I__6493 (
            .O(N__35718),
            .I(N__35675));
    InMux I__6492 (
            .O(N__35717),
            .I(N__35670));
    InMux I__6491 (
            .O(N__35716),
            .I(N__35670));
    InMux I__6490 (
            .O(N__35713),
            .I(N__35663));
    InMux I__6489 (
            .O(N__35710),
            .I(N__35663));
    InMux I__6488 (
            .O(N__35709),
            .I(N__35663));
    InMux I__6487 (
            .O(N__35708),
            .I(N__35656));
    InMux I__6486 (
            .O(N__35705),
            .I(N__35656));
    InMux I__6485 (
            .O(N__35704),
            .I(N__35656));
    InMux I__6484 (
            .O(N__35703),
            .I(N__35645));
    InMux I__6483 (
            .O(N__35702),
            .I(N__35645));
    InMux I__6482 (
            .O(N__35699),
            .I(N__35645));
    InMux I__6481 (
            .O(N__35696),
            .I(N__35645));
    InMux I__6480 (
            .O(N__35695),
            .I(N__35645));
    Odrv4 I__6479 (
            .O(N__35690),
            .I(n2346));
    LocalMux I__6478 (
            .O(N__35687),
            .I(n2346));
    Odrv4 I__6477 (
            .O(N__35684),
            .I(n2346));
    LocalMux I__6476 (
            .O(N__35675),
            .I(n2346));
    LocalMux I__6475 (
            .O(N__35670),
            .I(n2346));
    LocalMux I__6474 (
            .O(N__35663),
            .I(n2346));
    LocalMux I__6473 (
            .O(N__35656),
            .I(n2346));
    LocalMux I__6472 (
            .O(N__35645),
            .I(n2346));
    InMux I__6471 (
            .O(N__35628),
            .I(n12961));
    InMux I__6470 (
            .O(N__35625),
            .I(N__35622));
    LocalMux I__6469 (
            .O(N__35622),
            .I(N__35619));
    Span4Mux_v I__6468 (
            .O(N__35619),
            .I(N__35616));
    Span4Mux_v I__6467 (
            .O(N__35616),
            .I(N__35613));
    Span4Mux_h I__6466 (
            .O(N__35613),
            .I(N__35609));
    InMux I__6465 (
            .O(N__35612),
            .I(N__35606));
    Odrv4 I__6464 (
            .O(N__35609),
            .I(n15748));
    LocalMux I__6463 (
            .O(N__35606),
            .I(n15748));
    InMux I__6462 (
            .O(N__35601),
            .I(N__35598));
    LocalMux I__6461 (
            .O(N__35598),
            .I(N__35591));
    InMux I__6460 (
            .O(N__35597),
            .I(N__35584));
    CascadeMux I__6459 (
            .O(N__35596),
            .I(N__35581));
    CascadeMux I__6458 (
            .O(N__35595),
            .I(N__35578));
    CascadeMux I__6457 (
            .O(N__35594),
            .I(N__35575));
    Span4Mux_v I__6456 (
            .O(N__35591),
            .I(N__35570));
    CascadeMux I__6455 (
            .O(N__35590),
            .I(N__35567));
    CascadeMux I__6454 (
            .O(N__35589),
            .I(N__35563));
    CascadeMux I__6453 (
            .O(N__35588),
            .I(N__35558));
    CascadeMux I__6452 (
            .O(N__35587),
            .I(N__35555));
    LocalMux I__6451 (
            .O(N__35584),
            .I(N__35551));
    InMux I__6450 (
            .O(N__35581),
            .I(N__35542));
    InMux I__6449 (
            .O(N__35578),
            .I(N__35542));
    InMux I__6448 (
            .O(N__35575),
            .I(N__35542));
    InMux I__6447 (
            .O(N__35574),
            .I(N__35542));
    CascadeMux I__6446 (
            .O(N__35573),
            .I(N__35534));
    Span4Mux_h I__6445 (
            .O(N__35570),
            .I(N__35530));
    InMux I__6444 (
            .O(N__35567),
            .I(N__35525));
    InMux I__6443 (
            .O(N__35566),
            .I(N__35525));
    InMux I__6442 (
            .O(N__35563),
            .I(N__35518));
    InMux I__6441 (
            .O(N__35562),
            .I(N__35518));
    InMux I__6440 (
            .O(N__35561),
            .I(N__35518));
    InMux I__6439 (
            .O(N__35558),
            .I(N__35511));
    InMux I__6438 (
            .O(N__35555),
            .I(N__35511));
    InMux I__6437 (
            .O(N__35554),
            .I(N__35511));
    Span4Mux_h I__6436 (
            .O(N__35551),
            .I(N__35506));
    LocalMux I__6435 (
            .O(N__35542),
            .I(N__35506));
    InMux I__6434 (
            .O(N__35541),
            .I(N__35501));
    InMux I__6433 (
            .O(N__35540),
            .I(N__35501));
    InMux I__6432 (
            .O(N__35539),
            .I(N__35490));
    InMux I__6431 (
            .O(N__35538),
            .I(N__35490));
    InMux I__6430 (
            .O(N__35537),
            .I(N__35490));
    InMux I__6429 (
            .O(N__35534),
            .I(N__35490));
    InMux I__6428 (
            .O(N__35533),
            .I(N__35490));
    Odrv4 I__6427 (
            .O(N__35530),
            .I(n2247));
    LocalMux I__6426 (
            .O(N__35525),
            .I(n2247));
    LocalMux I__6425 (
            .O(N__35518),
            .I(n2247));
    LocalMux I__6424 (
            .O(N__35511),
            .I(n2247));
    Odrv4 I__6423 (
            .O(N__35506),
            .I(n2247));
    LocalMux I__6422 (
            .O(N__35501),
            .I(n2247));
    LocalMux I__6421 (
            .O(N__35490),
            .I(n2247));
    InMux I__6420 (
            .O(N__35475),
            .I(n12962));
    InMux I__6419 (
            .O(N__35472),
            .I(N__35469));
    LocalMux I__6418 (
            .O(N__35469),
            .I(N__35466));
    Span4Mux_h I__6417 (
            .O(N__35466),
            .I(N__35463));
    Span4Mux_v I__6416 (
            .O(N__35463),
            .I(N__35459));
    InMux I__6415 (
            .O(N__35462),
            .I(N__35456));
    Odrv4 I__6414 (
            .O(N__35459),
            .I(n15722));
    LocalMux I__6413 (
            .O(N__35456),
            .I(n15722));
    InMux I__6412 (
            .O(N__35451),
            .I(N__35448));
    LocalMux I__6411 (
            .O(N__35448),
            .I(N__35438));
    InMux I__6410 (
            .O(N__35447),
            .I(N__35433));
    CascadeMux I__6409 (
            .O(N__35446),
            .I(N__35430));
    CascadeMux I__6408 (
            .O(N__35445),
            .I(N__35427));
    CascadeMux I__6407 (
            .O(N__35444),
            .I(N__35424));
    CascadeMux I__6406 (
            .O(N__35443),
            .I(N__35421));
    CascadeMux I__6405 (
            .O(N__35442),
            .I(N__35413));
    CascadeMux I__6404 (
            .O(N__35441),
            .I(N__35410));
    Span4Mux_v I__6403 (
            .O(N__35438),
            .I(N__35405));
    InMux I__6402 (
            .O(N__35437),
            .I(N__35400));
    InMux I__6401 (
            .O(N__35436),
            .I(N__35400));
    LocalMux I__6400 (
            .O(N__35433),
            .I(N__35396));
    InMux I__6399 (
            .O(N__35430),
            .I(N__35391));
    InMux I__6398 (
            .O(N__35427),
            .I(N__35391));
    InMux I__6397 (
            .O(N__35424),
            .I(N__35380));
    InMux I__6396 (
            .O(N__35421),
            .I(N__35380));
    InMux I__6395 (
            .O(N__35420),
            .I(N__35380));
    InMux I__6394 (
            .O(N__35419),
            .I(N__35380));
    InMux I__6393 (
            .O(N__35418),
            .I(N__35380));
    InMux I__6392 (
            .O(N__35417),
            .I(N__35373));
    InMux I__6391 (
            .O(N__35416),
            .I(N__35373));
    InMux I__6390 (
            .O(N__35413),
            .I(N__35364));
    InMux I__6389 (
            .O(N__35410),
            .I(N__35364));
    InMux I__6388 (
            .O(N__35409),
            .I(N__35364));
    InMux I__6387 (
            .O(N__35408),
            .I(N__35364));
    Span4Mux_v I__6386 (
            .O(N__35405),
            .I(N__35359));
    LocalMux I__6385 (
            .O(N__35400),
            .I(N__35359));
    InMux I__6384 (
            .O(N__35399),
            .I(N__35356));
    Span4Mux_h I__6383 (
            .O(N__35396),
            .I(N__35353));
    LocalMux I__6382 (
            .O(N__35391),
            .I(N__35348));
    LocalMux I__6381 (
            .O(N__35380),
            .I(N__35348));
    InMux I__6380 (
            .O(N__35379),
            .I(N__35343));
    InMux I__6379 (
            .O(N__35378),
            .I(N__35343));
    LocalMux I__6378 (
            .O(N__35373),
            .I(n2148));
    LocalMux I__6377 (
            .O(N__35364),
            .I(n2148));
    Odrv4 I__6376 (
            .O(N__35359),
            .I(n2148));
    LocalMux I__6375 (
            .O(N__35356),
            .I(n2148));
    Odrv4 I__6374 (
            .O(N__35353),
            .I(n2148));
    Odrv4 I__6373 (
            .O(N__35348),
            .I(n2148));
    LocalMux I__6372 (
            .O(N__35343),
            .I(n2148));
    InMux I__6371 (
            .O(N__35328),
            .I(n12963));
    InMux I__6370 (
            .O(N__35325),
            .I(N__35322));
    LocalMux I__6369 (
            .O(N__35322),
            .I(N__35319));
    Span4Mux_h I__6368 (
            .O(N__35319),
            .I(N__35316));
    Span4Mux_v I__6367 (
            .O(N__35316),
            .I(N__35312));
    InMux I__6366 (
            .O(N__35315),
            .I(N__35309));
    Odrv4 I__6365 (
            .O(N__35312),
            .I(n15697));
    LocalMux I__6364 (
            .O(N__35309),
            .I(n15697));
    InMux I__6363 (
            .O(N__35304),
            .I(N__35299));
    CascadeMux I__6362 (
            .O(N__35303),
            .I(N__35293));
    CascadeMux I__6361 (
            .O(N__35302),
            .I(N__35289));
    LocalMux I__6360 (
            .O(N__35299),
            .I(N__35285));
    InMux I__6359 (
            .O(N__35298),
            .I(N__35282));
    InMux I__6358 (
            .O(N__35297),
            .I(N__35271));
    InMux I__6357 (
            .O(N__35296),
            .I(N__35271));
    InMux I__6356 (
            .O(N__35293),
            .I(N__35266));
    InMux I__6355 (
            .O(N__35292),
            .I(N__35266));
    InMux I__6354 (
            .O(N__35289),
            .I(N__35263));
    CascadeMux I__6353 (
            .O(N__35288),
            .I(N__35259));
    Span4Mux_v I__6352 (
            .O(N__35285),
            .I(N__35254));
    LocalMux I__6351 (
            .O(N__35282),
            .I(N__35251));
    CascadeMux I__6350 (
            .O(N__35281),
            .I(N__35248));
    CascadeMux I__6349 (
            .O(N__35280),
            .I(N__35245));
    InMux I__6348 (
            .O(N__35279),
            .I(N__35240));
    InMux I__6347 (
            .O(N__35278),
            .I(N__35233));
    InMux I__6346 (
            .O(N__35277),
            .I(N__35233));
    InMux I__6345 (
            .O(N__35276),
            .I(N__35233));
    LocalMux I__6344 (
            .O(N__35271),
            .I(N__35230));
    LocalMux I__6343 (
            .O(N__35266),
            .I(N__35225));
    LocalMux I__6342 (
            .O(N__35263),
            .I(N__35225));
    InMux I__6341 (
            .O(N__35262),
            .I(N__35218));
    InMux I__6340 (
            .O(N__35259),
            .I(N__35218));
    InMux I__6339 (
            .O(N__35258),
            .I(N__35218));
    InMux I__6338 (
            .O(N__35257),
            .I(N__35215));
    Span4Mux_v I__6337 (
            .O(N__35254),
            .I(N__35210));
    Span4Mux_v I__6336 (
            .O(N__35251),
            .I(N__35210));
    InMux I__6335 (
            .O(N__35248),
            .I(N__35203));
    InMux I__6334 (
            .O(N__35245),
            .I(N__35203));
    InMux I__6333 (
            .O(N__35244),
            .I(N__35203));
    InMux I__6332 (
            .O(N__35243),
            .I(N__35200));
    LocalMux I__6331 (
            .O(N__35240),
            .I(n2049));
    LocalMux I__6330 (
            .O(N__35233),
            .I(n2049));
    Odrv4 I__6329 (
            .O(N__35230),
            .I(n2049));
    Odrv4 I__6328 (
            .O(N__35225),
            .I(n2049));
    LocalMux I__6327 (
            .O(N__35218),
            .I(n2049));
    LocalMux I__6326 (
            .O(N__35215),
            .I(n2049));
    Odrv4 I__6325 (
            .O(N__35210),
            .I(n2049));
    LocalMux I__6324 (
            .O(N__35203),
            .I(n2049));
    LocalMux I__6323 (
            .O(N__35200),
            .I(n2049));
    InMux I__6322 (
            .O(N__35181),
            .I(n12964));
    InMux I__6321 (
            .O(N__35178),
            .I(N__35173));
    InMux I__6320 (
            .O(N__35177),
            .I(N__35170));
    InMux I__6319 (
            .O(N__35176),
            .I(N__35167));
    LocalMux I__6318 (
            .O(N__35173),
            .I(N__35164));
    LocalMux I__6317 (
            .O(N__35170),
            .I(N__35161));
    LocalMux I__6316 (
            .O(N__35167),
            .I(N__35158));
    Span4Mux_v I__6315 (
            .O(N__35164),
            .I(N__35153));
    Span4Mux_v I__6314 (
            .O(N__35161),
            .I(N__35153));
    Span4Mux_v I__6313 (
            .O(N__35158),
            .I(N__35148));
    Span4Mux_h I__6312 (
            .O(N__35153),
            .I(N__35148));
    Odrv4 I__6311 (
            .O(N__35148),
            .I(n315));
    InMux I__6310 (
            .O(N__35145),
            .I(N__35142));
    LocalMux I__6309 (
            .O(N__35142),
            .I(N__35138));
    InMux I__6308 (
            .O(N__35141),
            .I(N__35134));
    Span4Mux_h I__6307 (
            .O(N__35138),
            .I(N__35131));
    InMux I__6306 (
            .O(N__35137),
            .I(N__35128));
    LocalMux I__6305 (
            .O(N__35134),
            .I(N__35125));
    Odrv4 I__6304 (
            .O(N__35131),
            .I(n311));
    LocalMux I__6303 (
            .O(N__35128),
            .I(n311));
    Odrv4 I__6302 (
            .O(N__35125),
            .I(n311));
    InMux I__6301 (
            .O(N__35118),
            .I(bfn_7_25_0_));
    InMux I__6300 (
            .O(N__35115),
            .I(N__35112));
    LocalMux I__6299 (
            .O(N__35112),
            .I(N__35109));
    Span4Mux_h I__6298 (
            .O(N__35109),
            .I(N__35106));
    Odrv4 I__6297 (
            .O(N__35106),
            .I(n15485));
    InMux I__6296 (
            .O(N__35103),
            .I(N__35100));
    LocalMux I__6295 (
            .O(N__35100),
            .I(N__35096));
    InMux I__6294 (
            .O(N__35099),
            .I(N__35084));
    Span4Mux_v I__6293 (
            .O(N__35096),
            .I(N__35081));
    CascadeMux I__6292 (
            .O(N__35095),
            .I(N__35073));
    CascadeMux I__6291 (
            .O(N__35094),
            .I(N__35069));
    CascadeMux I__6290 (
            .O(N__35093),
            .I(N__35063));
    InMux I__6289 (
            .O(N__35092),
            .I(N__35058));
    InMux I__6288 (
            .O(N__35091),
            .I(N__35058));
    CascadeMux I__6287 (
            .O(N__35090),
            .I(N__35054));
    CascadeMux I__6286 (
            .O(N__35089),
            .I(N__35051));
    CascadeMux I__6285 (
            .O(N__35088),
            .I(N__35046));
    CascadeMux I__6284 (
            .O(N__35087),
            .I(N__35042));
    LocalMux I__6283 (
            .O(N__35084),
            .I(N__35032));
    Span4Mux_v I__6282 (
            .O(N__35081),
            .I(N__35029));
    InMux I__6281 (
            .O(N__35080),
            .I(N__35016));
    InMux I__6280 (
            .O(N__35079),
            .I(N__35016));
    InMux I__6279 (
            .O(N__35078),
            .I(N__35016));
    InMux I__6278 (
            .O(N__35077),
            .I(N__35016));
    InMux I__6277 (
            .O(N__35076),
            .I(N__35016));
    InMux I__6276 (
            .O(N__35073),
            .I(N__35016));
    InMux I__6275 (
            .O(N__35072),
            .I(N__35003));
    InMux I__6274 (
            .O(N__35069),
            .I(N__35003));
    InMux I__6273 (
            .O(N__35068),
            .I(N__35003));
    InMux I__6272 (
            .O(N__35067),
            .I(N__35003));
    InMux I__6271 (
            .O(N__35066),
            .I(N__35003));
    InMux I__6270 (
            .O(N__35063),
            .I(N__35003));
    LocalMux I__6269 (
            .O(N__35058),
            .I(N__35000));
    InMux I__6268 (
            .O(N__35057),
            .I(N__34987));
    InMux I__6267 (
            .O(N__35054),
            .I(N__34987));
    InMux I__6266 (
            .O(N__35051),
            .I(N__34987));
    InMux I__6265 (
            .O(N__35050),
            .I(N__34987));
    InMux I__6264 (
            .O(N__35049),
            .I(N__34987));
    InMux I__6263 (
            .O(N__35046),
            .I(N__34987));
    InMux I__6262 (
            .O(N__35045),
            .I(N__34980));
    InMux I__6261 (
            .O(N__35042),
            .I(N__34980));
    InMux I__6260 (
            .O(N__35041),
            .I(N__34980));
    InMux I__6259 (
            .O(N__35040),
            .I(N__34967));
    InMux I__6258 (
            .O(N__35039),
            .I(N__34967));
    InMux I__6257 (
            .O(N__35038),
            .I(N__34967));
    InMux I__6256 (
            .O(N__35037),
            .I(N__34967));
    InMux I__6255 (
            .O(N__35036),
            .I(N__34967));
    InMux I__6254 (
            .O(N__35035),
            .I(N__34967));
    Odrv4 I__6253 (
            .O(N__35032),
            .I(n3237));
    Odrv4 I__6252 (
            .O(N__35029),
            .I(n3237));
    LocalMux I__6251 (
            .O(N__35016),
            .I(n3237));
    LocalMux I__6250 (
            .O(N__35003),
            .I(n3237));
    Odrv4 I__6249 (
            .O(N__35000),
            .I(n3237));
    LocalMux I__6248 (
            .O(N__34987),
            .I(n3237));
    LocalMux I__6247 (
            .O(N__34980),
            .I(n3237));
    LocalMux I__6246 (
            .O(N__34967),
            .I(n3237));
    InMux I__6245 (
            .O(N__34950),
            .I(n12952));
    InMux I__6244 (
            .O(N__34947),
            .I(N__34944));
    LocalMux I__6243 (
            .O(N__34944),
            .I(N__34941));
    Span4Mux_v I__6242 (
            .O(N__34941),
            .I(N__34937));
    CascadeMux I__6241 (
            .O(N__34940),
            .I(N__34934));
    Span4Mux_h I__6240 (
            .O(N__34937),
            .I(N__34931));
    InMux I__6239 (
            .O(N__34934),
            .I(N__34928));
    Odrv4 I__6238 (
            .O(N__34931),
            .I(n15451));
    LocalMux I__6237 (
            .O(N__34928),
            .I(n15451));
    CascadeMux I__6236 (
            .O(N__34923),
            .I(N__34919));
    InMux I__6235 (
            .O(N__34922),
            .I(N__34912));
    InMux I__6234 (
            .O(N__34919),
            .I(N__34901));
    InMux I__6233 (
            .O(N__34918),
            .I(N__34901));
    InMux I__6232 (
            .O(N__34917),
            .I(N__34898));
    CascadeMux I__6231 (
            .O(N__34916),
            .I(N__34895));
    CascadeMux I__6230 (
            .O(N__34915),
            .I(N__34892));
    LocalMux I__6229 (
            .O(N__34912),
            .I(N__34885));
    InMux I__6228 (
            .O(N__34911),
            .I(N__34882));
    CascadeMux I__6227 (
            .O(N__34910),
            .I(N__34877));
    CascadeMux I__6226 (
            .O(N__34909),
            .I(N__34871));
    CascadeMux I__6225 (
            .O(N__34908),
            .I(N__34867));
    CascadeMux I__6224 (
            .O(N__34907),
            .I(N__34863));
    CascadeMux I__6223 (
            .O(N__34906),
            .I(N__34859));
    LocalMux I__6222 (
            .O(N__34901),
            .I(N__34855));
    LocalMux I__6221 (
            .O(N__34898),
            .I(N__34852));
    InMux I__6220 (
            .O(N__34895),
            .I(N__34843));
    InMux I__6219 (
            .O(N__34892),
            .I(N__34843));
    InMux I__6218 (
            .O(N__34891),
            .I(N__34843));
    InMux I__6217 (
            .O(N__34890),
            .I(N__34843));
    InMux I__6216 (
            .O(N__34889),
            .I(N__34840));
    CascadeMux I__6215 (
            .O(N__34888),
            .I(N__34836));
    Span4Mux_h I__6214 (
            .O(N__34885),
            .I(N__34832));
    LocalMux I__6213 (
            .O(N__34882),
            .I(N__34829));
    CascadeMux I__6212 (
            .O(N__34881),
            .I(N__34826));
    InMux I__6211 (
            .O(N__34880),
            .I(N__34814));
    InMux I__6210 (
            .O(N__34877),
            .I(N__34814));
    InMux I__6209 (
            .O(N__34876),
            .I(N__34814));
    InMux I__6208 (
            .O(N__34875),
            .I(N__34814));
    InMux I__6207 (
            .O(N__34874),
            .I(N__34807));
    InMux I__6206 (
            .O(N__34871),
            .I(N__34807));
    InMux I__6205 (
            .O(N__34870),
            .I(N__34807));
    InMux I__6204 (
            .O(N__34867),
            .I(N__34802));
    InMux I__6203 (
            .O(N__34866),
            .I(N__34802));
    InMux I__6202 (
            .O(N__34863),
            .I(N__34793));
    InMux I__6201 (
            .O(N__34862),
            .I(N__34793));
    InMux I__6200 (
            .O(N__34859),
            .I(N__34793));
    InMux I__6199 (
            .O(N__34858),
            .I(N__34793));
    Span4Mux_v I__6198 (
            .O(N__34855),
            .I(N__34790));
    Span4Mux_h I__6197 (
            .O(N__34852),
            .I(N__34783));
    LocalMux I__6196 (
            .O(N__34843),
            .I(N__34783));
    LocalMux I__6195 (
            .O(N__34840),
            .I(N__34783));
    InMux I__6194 (
            .O(N__34839),
            .I(N__34776));
    InMux I__6193 (
            .O(N__34836),
            .I(N__34776));
    InMux I__6192 (
            .O(N__34835),
            .I(N__34776));
    Span4Mux_v I__6191 (
            .O(N__34832),
            .I(N__34771));
    Span4Mux_s3_h I__6190 (
            .O(N__34829),
            .I(N__34771));
    InMux I__6189 (
            .O(N__34826),
            .I(N__34762));
    InMux I__6188 (
            .O(N__34825),
            .I(N__34762));
    InMux I__6187 (
            .O(N__34824),
            .I(N__34762));
    InMux I__6186 (
            .O(N__34823),
            .I(N__34762));
    LocalMux I__6185 (
            .O(N__34814),
            .I(n3138));
    LocalMux I__6184 (
            .O(N__34807),
            .I(n3138));
    LocalMux I__6183 (
            .O(N__34802),
            .I(n3138));
    LocalMux I__6182 (
            .O(N__34793),
            .I(n3138));
    Odrv4 I__6181 (
            .O(N__34790),
            .I(n3138));
    Odrv4 I__6180 (
            .O(N__34783),
            .I(n3138));
    LocalMux I__6179 (
            .O(N__34776),
            .I(n3138));
    Odrv4 I__6178 (
            .O(N__34771),
            .I(n3138));
    LocalMux I__6177 (
            .O(N__34762),
            .I(n3138));
    InMux I__6176 (
            .O(N__34743),
            .I(n12953));
    InMux I__6175 (
            .O(N__34740),
            .I(N__34736));
    InMux I__6174 (
            .O(N__34739),
            .I(N__34733));
    LocalMux I__6173 (
            .O(N__34736),
            .I(N__34730));
    LocalMux I__6172 (
            .O(N__34733),
            .I(N__34727));
    Span4Mux_h I__6171 (
            .O(N__34730),
            .I(N__34724));
    Span12Mux_s4_h I__6170 (
            .O(N__34727),
            .I(N__34721));
    Odrv4 I__6169 (
            .O(N__34724),
            .I(n15418));
    Odrv12 I__6168 (
            .O(N__34721),
            .I(n15418));
    CascadeMux I__6167 (
            .O(N__34716),
            .I(N__34711));
    InMux I__6166 (
            .O(N__34715),
            .I(N__34705));
    CascadeMux I__6165 (
            .O(N__34714),
            .I(N__34700));
    InMux I__6164 (
            .O(N__34711),
            .I(N__34690));
    InMux I__6163 (
            .O(N__34710),
            .I(N__34690));
    CascadeMux I__6162 (
            .O(N__34709),
            .I(N__34687));
    CascadeMux I__6161 (
            .O(N__34708),
            .I(N__34683));
    LocalMux I__6160 (
            .O(N__34705),
            .I(N__34678));
    InMux I__6159 (
            .O(N__34704),
            .I(N__34673));
    InMux I__6158 (
            .O(N__34703),
            .I(N__34673));
    InMux I__6157 (
            .O(N__34700),
            .I(N__34666));
    InMux I__6156 (
            .O(N__34699),
            .I(N__34666));
    InMux I__6155 (
            .O(N__34698),
            .I(N__34666));
    CascadeMux I__6154 (
            .O(N__34697),
            .I(N__34661));
    CascadeMux I__6153 (
            .O(N__34696),
            .I(N__34654));
    CascadeMux I__6152 (
            .O(N__34695),
            .I(N__34650));
    LocalMux I__6151 (
            .O(N__34690),
            .I(N__34646));
    InMux I__6150 (
            .O(N__34687),
            .I(N__34635));
    InMux I__6149 (
            .O(N__34686),
            .I(N__34635));
    InMux I__6148 (
            .O(N__34683),
            .I(N__34635));
    InMux I__6147 (
            .O(N__34682),
            .I(N__34635));
    InMux I__6146 (
            .O(N__34681),
            .I(N__34635));
    Span4Mux_v I__6145 (
            .O(N__34678),
            .I(N__34632));
    LocalMux I__6144 (
            .O(N__34673),
            .I(N__34627));
    LocalMux I__6143 (
            .O(N__34666),
            .I(N__34627));
    InMux I__6142 (
            .O(N__34665),
            .I(N__34620));
    InMux I__6141 (
            .O(N__34664),
            .I(N__34620));
    InMux I__6140 (
            .O(N__34661),
            .I(N__34620));
    InMux I__6139 (
            .O(N__34660),
            .I(N__34617));
    InMux I__6138 (
            .O(N__34659),
            .I(N__34614));
    CascadeMux I__6137 (
            .O(N__34658),
            .I(N__34608));
    CascadeMux I__6136 (
            .O(N__34657),
            .I(N__34605));
    InMux I__6135 (
            .O(N__34654),
            .I(N__34594));
    InMux I__6134 (
            .O(N__34653),
            .I(N__34594));
    InMux I__6133 (
            .O(N__34650),
            .I(N__34594));
    InMux I__6132 (
            .O(N__34649),
            .I(N__34594));
    Span4Mux_s1_h I__6131 (
            .O(N__34646),
            .I(N__34589));
    LocalMux I__6130 (
            .O(N__34635),
            .I(N__34589));
    Span4Mux_h I__6129 (
            .O(N__34632),
            .I(N__34582));
    Span4Mux_s1_v I__6128 (
            .O(N__34627),
            .I(N__34582));
    LocalMux I__6127 (
            .O(N__34620),
            .I(N__34582));
    LocalMux I__6126 (
            .O(N__34617),
            .I(N__34579));
    LocalMux I__6125 (
            .O(N__34614),
            .I(N__34576));
    InMux I__6124 (
            .O(N__34613),
            .I(N__34563));
    InMux I__6123 (
            .O(N__34612),
            .I(N__34563));
    InMux I__6122 (
            .O(N__34611),
            .I(N__34563));
    InMux I__6121 (
            .O(N__34608),
            .I(N__34563));
    InMux I__6120 (
            .O(N__34605),
            .I(N__34563));
    InMux I__6119 (
            .O(N__34604),
            .I(N__34563));
    InMux I__6118 (
            .O(N__34603),
            .I(N__34560));
    LocalMux I__6117 (
            .O(N__34594),
            .I(N__34555));
    Span4Mux_v I__6116 (
            .O(N__34589),
            .I(N__34555));
    Odrv4 I__6115 (
            .O(N__34582),
            .I(n3039));
    Odrv4 I__6114 (
            .O(N__34579),
            .I(n3039));
    Odrv4 I__6113 (
            .O(N__34576),
            .I(n3039));
    LocalMux I__6112 (
            .O(N__34563),
            .I(n3039));
    LocalMux I__6111 (
            .O(N__34560),
            .I(n3039));
    Odrv4 I__6110 (
            .O(N__34555),
            .I(n3039));
    InMux I__6109 (
            .O(N__34542),
            .I(n12954));
    InMux I__6108 (
            .O(N__34539),
            .I(N__34536));
    LocalMux I__6107 (
            .O(N__34536),
            .I(N__34533));
    Span4Mux_h I__6106 (
            .O(N__34533),
            .I(N__34529));
    CascadeMux I__6105 (
            .O(N__34532),
            .I(N__34526));
    Span4Mux_h I__6104 (
            .O(N__34529),
            .I(N__34523));
    InMux I__6103 (
            .O(N__34526),
            .I(N__34520));
    Odrv4 I__6102 (
            .O(N__34523),
            .I(n15384));
    LocalMux I__6101 (
            .O(N__34520),
            .I(n15384));
    InMux I__6100 (
            .O(N__34515),
            .I(N__34506));
    InMux I__6099 (
            .O(N__34514),
            .I(N__34499));
    InMux I__6098 (
            .O(N__34513),
            .I(N__34494));
    InMux I__6097 (
            .O(N__34512),
            .I(N__34494));
    CascadeMux I__6096 (
            .O(N__34511),
            .I(N__34490));
    CascadeMux I__6095 (
            .O(N__34510),
            .I(N__34487));
    CascadeMux I__6094 (
            .O(N__34509),
            .I(N__34484));
    LocalMux I__6093 (
            .O(N__34506),
            .I(N__34480));
    InMux I__6092 (
            .O(N__34505),
            .I(N__34476));
    CascadeMux I__6091 (
            .O(N__34504),
            .I(N__34469));
    CascadeMux I__6090 (
            .O(N__34503),
            .I(N__34463));
    CascadeMux I__6089 (
            .O(N__34502),
            .I(N__34455));
    LocalMux I__6088 (
            .O(N__34499),
            .I(N__34450));
    LocalMux I__6087 (
            .O(N__34494),
            .I(N__34447));
    InMux I__6086 (
            .O(N__34493),
            .I(N__34436));
    InMux I__6085 (
            .O(N__34490),
            .I(N__34436));
    InMux I__6084 (
            .O(N__34487),
            .I(N__34436));
    InMux I__6083 (
            .O(N__34484),
            .I(N__34436));
    InMux I__6082 (
            .O(N__34483),
            .I(N__34436));
    Span4Mux_h I__6081 (
            .O(N__34480),
            .I(N__34433));
    InMux I__6080 (
            .O(N__34479),
            .I(N__34430));
    LocalMux I__6079 (
            .O(N__34476),
            .I(N__34427));
    InMux I__6078 (
            .O(N__34475),
            .I(N__34420));
    InMux I__6077 (
            .O(N__34474),
            .I(N__34420));
    InMux I__6076 (
            .O(N__34473),
            .I(N__34420));
    InMux I__6075 (
            .O(N__34472),
            .I(N__34413));
    InMux I__6074 (
            .O(N__34469),
            .I(N__34413));
    InMux I__6073 (
            .O(N__34468),
            .I(N__34413));
    InMux I__6072 (
            .O(N__34467),
            .I(N__34406));
    InMux I__6071 (
            .O(N__34466),
            .I(N__34406));
    InMux I__6070 (
            .O(N__34463),
            .I(N__34406));
    InMux I__6069 (
            .O(N__34462),
            .I(N__34403));
    InMux I__6068 (
            .O(N__34461),
            .I(N__34398));
    InMux I__6067 (
            .O(N__34460),
            .I(N__34398));
    InMux I__6066 (
            .O(N__34459),
            .I(N__34387));
    InMux I__6065 (
            .O(N__34458),
            .I(N__34387));
    InMux I__6064 (
            .O(N__34455),
            .I(N__34387));
    InMux I__6063 (
            .O(N__34454),
            .I(N__34387));
    InMux I__6062 (
            .O(N__34453),
            .I(N__34387));
    Span4Mux_v I__6061 (
            .O(N__34450),
            .I(N__34380));
    Span4Mux_v I__6060 (
            .O(N__34447),
            .I(N__34380));
    LocalMux I__6059 (
            .O(N__34436),
            .I(N__34380));
    Odrv4 I__6058 (
            .O(N__34433),
            .I(n2940));
    LocalMux I__6057 (
            .O(N__34430),
            .I(n2940));
    Odrv4 I__6056 (
            .O(N__34427),
            .I(n2940));
    LocalMux I__6055 (
            .O(N__34420),
            .I(n2940));
    LocalMux I__6054 (
            .O(N__34413),
            .I(n2940));
    LocalMux I__6053 (
            .O(N__34406),
            .I(n2940));
    LocalMux I__6052 (
            .O(N__34403),
            .I(n2940));
    LocalMux I__6051 (
            .O(N__34398),
            .I(n2940));
    LocalMux I__6050 (
            .O(N__34387),
            .I(n2940));
    Odrv4 I__6049 (
            .O(N__34380),
            .I(n2940));
    InMux I__6048 (
            .O(N__34359),
            .I(n12955));
    InMux I__6047 (
            .O(N__34356),
            .I(N__34353));
    LocalMux I__6046 (
            .O(N__34353),
            .I(N__34349));
    InMux I__6045 (
            .O(N__34352),
            .I(N__34346));
    Span4Mux_h I__6044 (
            .O(N__34349),
            .I(N__34341));
    LocalMux I__6043 (
            .O(N__34346),
            .I(N__34341));
    Span4Mux_s3_h I__6042 (
            .O(N__34341),
            .I(N__34338));
    Odrv4 I__6041 (
            .O(N__34338),
            .I(n15352));
    CascadeMux I__6040 (
            .O(N__34335),
            .I(N__34329));
    InMux I__6039 (
            .O(N__34334),
            .I(N__34325));
    CascadeMux I__6038 (
            .O(N__34333),
            .I(N__34317));
    InMux I__6037 (
            .O(N__34332),
            .I(N__34311));
    InMux I__6036 (
            .O(N__34329),
            .I(N__34306));
    InMux I__6035 (
            .O(N__34328),
            .I(N__34306));
    LocalMux I__6034 (
            .O(N__34325),
            .I(N__34303));
    CascadeMux I__6033 (
            .O(N__34324),
            .I(N__34298));
    CascadeMux I__6032 (
            .O(N__34323),
            .I(N__34294));
    InMux I__6031 (
            .O(N__34322),
            .I(N__34286));
    CascadeMux I__6030 (
            .O(N__34321),
            .I(N__34283));
    CascadeMux I__6029 (
            .O(N__34320),
            .I(N__34279));
    InMux I__6028 (
            .O(N__34317),
            .I(N__34272));
    InMux I__6027 (
            .O(N__34316),
            .I(N__34272));
    CascadeMux I__6026 (
            .O(N__34315),
            .I(N__34268));
    CascadeMux I__6025 (
            .O(N__34314),
            .I(N__34264));
    LocalMux I__6024 (
            .O(N__34311),
            .I(N__34260));
    LocalMux I__6023 (
            .O(N__34306),
            .I(N__34257));
    Span4Mux_h I__6022 (
            .O(N__34303),
            .I(N__34254));
    InMux I__6021 (
            .O(N__34302),
            .I(N__34249));
    InMux I__6020 (
            .O(N__34301),
            .I(N__34249));
    InMux I__6019 (
            .O(N__34298),
            .I(N__34244));
    InMux I__6018 (
            .O(N__34297),
            .I(N__34244));
    InMux I__6017 (
            .O(N__34294),
            .I(N__34239));
    InMux I__6016 (
            .O(N__34293),
            .I(N__34239));
    InMux I__6015 (
            .O(N__34292),
            .I(N__34230));
    InMux I__6014 (
            .O(N__34291),
            .I(N__34230));
    InMux I__6013 (
            .O(N__34290),
            .I(N__34230));
    InMux I__6012 (
            .O(N__34289),
            .I(N__34230));
    LocalMux I__6011 (
            .O(N__34286),
            .I(N__34227));
    InMux I__6010 (
            .O(N__34283),
            .I(N__34222));
    InMux I__6009 (
            .O(N__34282),
            .I(N__34222));
    InMux I__6008 (
            .O(N__34279),
            .I(N__34215));
    InMux I__6007 (
            .O(N__34278),
            .I(N__34215));
    InMux I__6006 (
            .O(N__34277),
            .I(N__34215));
    LocalMux I__6005 (
            .O(N__34272),
            .I(N__34212));
    InMux I__6004 (
            .O(N__34271),
            .I(N__34201));
    InMux I__6003 (
            .O(N__34268),
            .I(N__34201));
    InMux I__6002 (
            .O(N__34267),
            .I(N__34201));
    InMux I__6001 (
            .O(N__34264),
            .I(N__34201));
    InMux I__6000 (
            .O(N__34263),
            .I(N__34201));
    Span4Mux_v I__5999 (
            .O(N__34260),
            .I(N__34196));
    Span4Mux_s3_h I__5998 (
            .O(N__34257),
            .I(N__34196));
    Odrv4 I__5997 (
            .O(N__34254),
            .I(n2841));
    LocalMux I__5996 (
            .O(N__34249),
            .I(n2841));
    LocalMux I__5995 (
            .O(N__34244),
            .I(n2841));
    LocalMux I__5994 (
            .O(N__34239),
            .I(n2841));
    LocalMux I__5993 (
            .O(N__34230),
            .I(n2841));
    Odrv4 I__5992 (
            .O(N__34227),
            .I(n2841));
    LocalMux I__5991 (
            .O(N__34222),
            .I(n2841));
    LocalMux I__5990 (
            .O(N__34215),
            .I(n2841));
    Odrv4 I__5989 (
            .O(N__34212),
            .I(n2841));
    LocalMux I__5988 (
            .O(N__34201),
            .I(n2841));
    Odrv4 I__5987 (
            .O(N__34196),
            .I(n2841));
    InMux I__5986 (
            .O(N__34173),
            .I(n12956));
    InMux I__5985 (
            .O(N__34170),
            .I(N__34167));
    LocalMux I__5984 (
            .O(N__34167),
            .I(N__34162));
    InMux I__5983 (
            .O(N__34166),
            .I(N__34159));
    InMux I__5982 (
            .O(N__34165),
            .I(N__34156));
    Span4Mux_s3_h I__5981 (
            .O(N__34162),
            .I(N__34151));
    LocalMux I__5980 (
            .O(N__34159),
            .I(N__34151));
    LocalMux I__5979 (
            .O(N__34156),
            .I(N__34148));
    Span4Mux_h I__5978 (
            .O(N__34151),
            .I(N__34145));
    Sp12to4 I__5977 (
            .O(N__34148),
            .I(N__34142));
    Span4Mux_v I__5976 (
            .O(N__34145),
            .I(N__34139));
    Odrv12 I__5975 (
            .O(N__34142),
            .I(n317));
    Odrv4 I__5974 (
            .O(N__34139),
            .I(n317));
    InMux I__5973 (
            .O(N__34134),
            .I(N__34131));
    LocalMux I__5972 (
            .O(N__34131),
            .I(N__34128));
    Odrv4 I__5971 (
            .O(N__34128),
            .I(n14184));
    InMux I__5970 (
            .O(N__34125),
            .I(N__34122));
    LocalMux I__5969 (
            .O(N__34122),
            .I(n2490));
    CascadeMux I__5968 (
            .O(N__34119),
            .I(N__34115));
    InMux I__5967 (
            .O(N__34118),
            .I(N__34112));
    InMux I__5966 (
            .O(N__34115),
            .I(N__34109));
    LocalMux I__5965 (
            .O(N__34112),
            .I(N__34106));
    LocalMux I__5964 (
            .O(N__34109),
            .I(N__34103));
    Span4Mux_v I__5963 (
            .O(N__34106),
            .I(N__34099));
    Span4Mux_h I__5962 (
            .O(N__34103),
            .I(N__34096));
    InMux I__5961 (
            .O(N__34102),
            .I(N__34093));
    Odrv4 I__5960 (
            .O(N__34099),
            .I(n2423));
    Odrv4 I__5959 (
            .O(N__34096),
            .I(n2423));
    LocalMux I__5958 (
            .O(N__34093),
            .I(n2423));
    InMux I__5957 (
            .O(N__34086),
            .I(N__34083));
    LocalMux I__5956 (
            .O(N__34083),
            .I(N__34079));
    CascadeMux I__5955 (
            .O(N__34082),
            .I(N__34076));
    Span4Mux_v I__5954 (
            .O(N__34079),
            .I(N__34072));
    InMux I__5953 (
            .O(N__34076),
            .I(N__34069));
    CascadeMux I__5952 (
            .O(N__34075),
            .I(N__34066));
    Span4Mux_h I__5951 (
            .O(N__34072),
            .I(N__34061));
    LocalMux I__5950 (
            .O(N__34069),
            .I(N__34061));
    InMux I__5949 (
            .O(N__34066),
            .I(N__34058));
    Odrv4 I__5948 (
            .O(N__34061),
            .I(n2522));
    LocalMux I__5947 (
            .O(N__34058),
            .I(n2522));
    InMux I__5946 (
            .O(N__34053),
            .I(N__34050));
    LocalMux I__5945 (
            .O(N__34050),
            .I(n2489));
    CascadeMux I__5944 (
            .O(N__34047),
            .I(N__34044));
    InMux I__5943 (
            .O(N__34044),
            .I(N__34040));
    CascadeMux I__5942 (
            .O(N__34043),
            .I(N__34037));
    LocalMux I__5941 (
            .O(N__34040),
            .I(N__34034));
    InMux I__5940 (
            .O(N__34037),
            .I(N__34031));
    Span4Mux_v I__5939 (
            .O(N__34034),
            .I(N__34027));
    LocalMux I__5938 (
            .O(N__34031),
            .I(N__34024));
    InMux I__5937 (
            .O(N__34030),
            .I(N__34021));
    Odrv4 I__5936 (
            .O(N__34027),
            .I(n2422));
    Odrv4 I__5935 (
            .O(N__34024),
            .I(n2422));
    LocalMux I__5934 (
            .O(N__34021),
            .I(n2422));
    CascadeMux I__5933 (
            .O(N__34014),
            .I(N__34011));
    InMux I__5932 (
            .O(N__34011),
            .I(N__34007));
    CascadeMux I__5931 (
            .O(N__34010),
            .I(N__34004));
    LocalMux I__5930 (
            .O(N__34007),
            .I(N__34001));
    InMux I__5929 (
            .O(N__34004),
            .I(N__33998));
    Span4Mux_h I__5928 (
            .O(N__34001),
            .I(N__33992));
    LocalMux I__5927 (
            .O(N__33998),
            .I(N__33992));
    InMux I__5926 (
            .O(N__33997),
            .I(N__33989));
    Odrv4 I__5925 (
            .O(N__33992),
            .I(n2521));
    LocalMux I__5924 (
            .O(N__33989),
            .I(n2521));
    CascadeMux I__5923 (
            .O(N__33984),
            .I(N__33980));
    InMux I__5922 (
            .O(N__33983),
            .I(N__33977));
    InMux I__5921 (
            .O(N__33980),
            .I(N__33974));
    LocalMux I__5920 (
            .O(N__33977),
            .I(N__33969));
    LocalMux I__5919 (
            .O(N__33974),
            .I(N__33969));
    Span4Mux_v I__5918 (
            .O(N__33969),
            .I(N__33965));
    InMux I__5917 (
            .O(N__33968),
            .I(N__33962));
    Odrv4 I__5916 (
            .O(N__33965),
            .I(n2426));
    LocalMux I__5915 (
            .O(N__33962),
            .I(n2426));
    InMux I__5914 (
            .O(N__33957),
            .I(N__33954));
    LocalMux I__5913 (
            .O(N__33954),
            .I(n2493));
    CascadeMux I__5912 (
            .O(N__33951),
            .I(N__33948));
    InMux I__5911 (
            .O(N__33948),
            .I(N__33945));
    LocalMux I__5910 (
            .O(N__33945),
            .I(N__33941));
    InMux I__5909 (
            .O(N__33944),
            .I(N__33938));
    Odrv4 I__5908 (
            .O(N__33941),
            .I(n2525));
    LocalMux I__5907 (
            .O(N__33938),
            .I(n2525));
    InMux I__5906 (
            .O(N__33933),
            .I(N__33930));
    LocalMux I__5905 (
            .O(N__33930),
            .I(N__33927));
    Odrv4 I__5904 (
            .O(N__33927),
            .I(n2592));
    CascadeMux I__5903 (
            .O(N__33924),
            .I(n2525_cascade_));
    CascadeMux I__5902 (
            .O(N__33921),
            .I(N__33918));
    InMux I__5901 (
            .O(N__33918),
            .I(N__33914));
    InMux I__5900 (
            .O(N__33917),
            .I(N__33911));
    LocalMux I__5899 (
            .O(N__33914),
            .I(N__33908));
    LocalMux I__5898 (
            .O(N__33911),
            .I(N__33904));
    Span4Mux_v I__5897 (
            .O(N__33908),
            .I(N__33901));
    InMux I__5896 (
            .O(N__33907),
            .I(N__33898));
    Span4Mux_v I__5895 (
            .O(N__33904),
            .I(N__33891));
    Span4Mux_v I__5894 (
            .O(N__33901),
            .I(N__33891));
    LocalMux I__5893 (
            .O(N__33898),
            .I(N__33891));
    Span4Mux_h I__5892 (
            .O(N__33891),
            .I(N__33888));
    Odrv4 I__5891 (
            .O(N__33888),
            .I(n2624));
    InMux I__5890 (
            .O(N__33885),
            .I(N__33882));
    LocalMux I__5889 (
            .O(N__33882),
            .I(n2486));
    CascadeMux I__5888 (
            .O(N__33879),
            .I(N__33875));
    CascadeMux I__5887 (
            .O(N__33878),
            .I(N__33872));
    InMux I__5886 (
            .O(N__33875),
            .I(N__33868));
    InMux I__5885 (
            .O(N__33872),
            .I(N__33865));
    CascadeMux I__5884 (
            .O(N__33871),
            .I(N__33862));
    LocalMux I__5883 (
            .O(N__33868),
            .I(N__33859));
    LocalMux I__5882 (
            .O(N__33865),
            .I(N__33856));
    InMux I__5881 (
            .O(N__33862),
            .I(N__33853));
    Span4Mux_v I__5880 (
            .O(N__33859),
            .I(N__33850));
    Span4Mux_h I__5879 (
            .O(N__33856),
            .I(N__33845));
    LocalMux I__5878 (
            .O(N__33853),
            .I(N__33845));
    Odrv4 I__5877 (
            .O(N__33850),
            .I(n2419));
    Odrv4 I__5876 (
            .O(N__33845),
            .I(n2419));
    InMux I__5875 (
            .O(N__33840),
            .I(N__33836));
    InMux I__5874 (
            .O(N__33839),
            .I(N__33833));
    LocalMux I__5873 (
            .O(N__33836),
            .I(N__33829));
    LocalMux I__5872 (
            .O(N__33833),
            .I(N__33826));
    InMux I__5871 (
            .O(N__33832),
            .I(N__33823));
    Odrv4 I__5870 (
            .O(N__33829),
            .I(n2518));
    Odrv4 I__5869 (
            .O(N__33826),
            .I(n2518));
    LocalMux I__5868 (
            .O(N__33823),
            .I(n2518));
    InMux I__5867 (
            .O(N__33816),
            .I(N__33813));
    LocalMux I__5866 (
            .O(N__33813),
            .I(n11981));
    InMux I__5865 (
            .O(N__33810),
            .I(N__33807));
    LocalMux I__5864 (
            .O(N__33807),
            .I(N__33802));
    CascadeMux I__5863 (
            .O(N__33806),
            .I(N__33799));
    InMux I__5862 (
            .O(N__33805),
            .I(N__33796));
    Span4Mux_h I__5861 (
            .O(N__33802),
            .I(N__33793));
    InMux I__5860 (
            .O(N__33799),
            .I(N__33790));
    LocalMux I__5859 (
            .O(N__33796),
            .I(N__33787));
    Odrv4 I__5858 (
            .O(N__33793),
            .I(n2029));
    LocalMux I__5857 (
            .O(N__33790),
            .I(n2029));
    Odrv4 I__5856 (
            .O(N__33787),
            .I(n2029));
    CascadeMux I__5855 (
            .O(N__33780),
            .I(n14550_cascade_));
    InMux I__5854 (
            .O(N__33777),
            .I(N__33772));
    CascadeMux I__5853 (
            .O(N__33776),
            .I(N__33769));
    InMux I__5852 (
            .O(N__33775),
            .I(N__33766));
    LocalMux I__5851 (
            .O(N__33772),
            .I(N__33763));
    InMux I__5850 (
            .O(N__33769),
            .I(N__33760));
    LocalMux I__5849 (
            .O(N__33766),
            .I(N__33757));
    Odrv4 I__5848 (
            .O(N__33763),
            .I(n2030));
    LocalMux I__5847 (
            .O(N__33760),
            .I(n2030));
    Odrv12 I__5846 (
            .O(N__33757),
            .I(n2030));
    InMux I__5845 (
            .O(N__33750),
            .I(N__33747));
    LocalMux I__5844 (
            .O(N__33747),
            .I(n14552));
    InMux I__5843 (
            .O(N__33744),
            .I(N__33741));
    LocalMux I__5842 (
            .O(N__33741),
            .I(N__33738));
    Span4Mux_v I__5841 (
            .O(N__33738),
            .I(N__33735));
    Odrv4 I__5840 (
            .O(N__33735),
            .I(n2100));
    CascadeMux I__5839 (
            .O(N__33732),
            .I(N__33728));
    CascadeMux I__5838 (
            .O(N__33731),
            .I(N__33725));
    InMux I__5837 (
            .O(N__33728),
            .I(N__33722));
    InMux I__5836 (
            .O(N__33725),
            .I(N__33718));
    LocalMux I__5835 (
            .O(N__33722),
            .I(N__33715));
    InMux I__5834 (
            .O(N__33721),
            .I(N__33712));
    LocalMux I__5833 (
            .O(N__33718),
            .I(n2033));
    Odrv4 I__5832 (
            .O(N__33715),
            .I(n2033));
    LocalMux I__5831 (
            .O(N__33712),
            .I(n2033));
    InMux I__5830 (
            .O(N__33705),
            .I(N__33701));
    CascadeMux I__5829 (
            .O(N__33704),
            .I(N__33698));
    LocalMux I__5828 (
            .O(N__33701),
            .I(N__33695));
    InMux I__5827 (
            .O(N__33698),
            .I(N__33692));
    Span4Mux_v I__5826 (
            .O(N__33695),
            .I(N__33687));
    LocalMux I__5825 (
            .O(N__33692),
            .I(N__33687));
    Span4Mux_v I__5824 (
            .O(N__33687),
            .I(N__33684));
    Odrv4 I__5823 (
            .O(N__33684),
            .I(n2132));
    CascadeMux I__5822 (
            .O(N__33681),
            .I(n2132_cascade_));
    CascadeMux I__5821 (
            .O(N__33678),
            .I(N__33674));
    InMux I__5820 (
            .O(N__33677),
            .I(N__33671));
    InMux I__5819 (
            .O(N__33674),
            .I(N__33668));
    LocalMux I__5818 (
            .O(N__33671),
            .I(N__33665));
    LocalMux I__5817 (
            .O(N__33668),
            .I(N__33662));
    Span12Mux_v I__5816 (
            .O(N__33665),
            .I(N__33658));
    Span4Mux_h I__5815 (
            .O(N__33662),
            .I(N__33655));
    InMux I__5814 (
            .O(N__33661),
            .I(N__33652));
    Odrv12 I__5813 (
            .O(N__33658),
            .I(n2133));
    Odrv4 I__5812 (
            .O(N__33655),
            .I(n2133));
    LocalMux I__5811 (
            .O(N__33652),
            .I(n2133));
    InMux I__5810 (
            .O(N__33645),
            .I(N__33642));
    LocalMux I__5809 (
            .O(N__33642),
            .I(N__33639));
    Span4Mux_h I__5808 (
            .O(N__33639),
            .I(N__33636));
    Odrv4 I__5807 (
            .O(N__33636),
            .I(n11909));
    InMux I__5806 (
            .O(N__33633),
            .I(N__33629));
    InMux I__5805 (
            .O(N__33632),
            .I(N__33626));
    LocalMux I__5804 (
            .O(N__33629),
            .I(N__33621));
    LocalMux I__5803 (
            .O(N__33626),
            .I(N__33621));
    Span4Mux_h I__5802 (
            .O(N__33621),
            .I(N__33617));
    InMux I__5801 (
            .O(N__33620),
            .I(N__33614));
    Odrv4 I__5800 (
            .O(N__33617),
            .I(n307));
    LocalMux I__5799 (
            .O(N__33614),
            .I(n307));
    InMux I__5798 (
            .O(N__33609),
            .I(N__33606));
    LocalMux I__5797 (
            .O(N__33606),
            .I(N__33602));
    InMux I__5796 (
            .O(N__33605),
            .I(N__33598));
    Span4Mux_h I__5795 (
            .O(N__33602),
            .I(N__33595));
    InMux I__5794 (
            .O(N__33601),
            .I(N__33592));
    LocalMux I__5793 (
            .O(N__33598),
            .I(N__33589));
    Odrv4 I__5792 (
            .O(N__33595),
            .I(n310));
    LocalMux I__5791 (
            .O(N__33592),
            .I(n310));
    Odrv12 I__5790 (
            .O(N__33589),
            .I(n310));
    InMux I__5789 (
            .O(N__33582),
            .I(N__33578));
    InMux I__5788 (
            .O(N__33581),
            .I(N__33574));
    LocalMux I__5787 (
            .O(N__33578),
            .I(N__33571));
    InMux I__5786 (
            .O(N__33577),
            .I(N__33568));
    LocalMux I__5785 (
            .O(N__33574),
            .I(N__33565));
    Span4Mux_s2_h I__5784 (
            .O(N__33571),
            .I(N__33562));
    LocalMux I__5783 (
            .O(N__33568),
            .I(N__33559));
    Span4Mux_v I__5782 (
            .O(N__33565),
            .I(N__33556));
    Span4Mux_v I__5781 (
            .O(N__33562),
            .I(N__33553));
    Span4Mux_v I__5780 (
            .O(N__33559),
            .I(N__33548));
    Span4Mux_s3_h I__5779 (
            .O(N__33556),
            .I(N__33548));
    Span4Mux_h I__5778 (
            .O(N__33553),
            .I(N__33545));
    Odrv4 I__5777 (
            .O(N__33548),
            .I(n312));
    Odrv4 I__5776 (
            .O(N__33545),
            .I(n312));
    InMux I__5775 (
            .O(N__33540),
            .I(N__33536));
    InMux I__5774 (
            .O(N__33539),
            .I(N__33533));
    LocalMux I__5773 (
            .O(N__33536),
            .I(N__33530));
    LocalMux I__5772 (
            .O(N__33533),
            .I(N__33527));
    Span4Mux_v I__5771 (
            .O(N__33530),
            .I(N__33524));
    Span4Mux_v I__5770 (
            .O(N__33527),
            .I(N__33520));
    Span4Mux_h I__5769 (
            .O(N__33524),
            .I(N__33517));
    InMux I__5768 (
            .O(N__33523),
            .I(N__33514));
    Span4Mux_h I__5767 (
            .O(N__33520),
            .I(N__33509));
    Span4Mux_v I__5766 (
            .O(N__33517),
            .I(N__33509));
    LocalMux I__5765 (
            .O(N__33514),
            .I(N__33506));
    Odrv4 I__5764 (
            .O(N__33509),
            .I(n313));
    Odrv12 I__5763 (
            .O(N__33506),
            .I(n313));
    InMux I__5762 (
            .O(N__33501),
            .I(N__33497));
    InMux I__5761 (
            .O(N__33500),
            .I(N__33493));
    LocalMux I__5760 (
            .O(N__33497),
            .I(N__33490));
    InMux I__5759 (
            .O(N__33496),
            .I(N__33487));
    LocalMux I__5758 (
            .O(N__33493),
            .I(N__33484));
    Span4Mux_s1_h I__5757 (
            .O(N__33490),
            .I(N__33481));
    LocalMux I__5756 (
            .O(N__33487),
            .I(N__33478));
    Span4Mux_v I__5755 (
            .O(N__33484),
            .I(N__33473));
    Span4Mux_h I__5754 (
            .O(N__33481),
            .I(N__33473));
    Span4Mux_h I__5753 (
            .O(N__33478),
            .I(N__33470));
    Odrv4 I__5752 (
            .O(N__33473),
            .I(n314));
    Odrv4 I__5751 (
            .O(N__33470),
            .I(n314));
    InMux I__5750 (
            .O(N__33465),
            .I(N__33461));
    CascadeMux I__5749 (
            .O(N__33464),
            .I(N__33458));
    LocalMux I__5748 (
            .O(N__33461),
            .I(N__33455));
    InMux I__5747 (
            .O(N__33458),
            .I(N__33452));
    Odrv4 I__5746 (
            .O(N__33455),
            .I(n2025));
    LocalMux I__5745 (
            .O(N__33452),
            .I(n2025));
    InMux I__5744 (
            .O(N__33447),
            .I(N__33444));
    LocalMux I__5743 (
            .O(N__33444),
            .I(N__33440));
    CascadeMux I__5742 (
            .O(N__33443),
            .I(N__33437));
    Span4Mux_v I__5741 (
            .O(N__33440),
            .I(N__33433));
    InMux I__5740 (
            .O(N__33437),
            .I(N__33430));
    InMux I__5739 (
            .O(N__33436),
            .I(N__33427));
    Odrv4 I__5738 (
            .O(N__33433),
            .I(n2028));
    LocalMux I__5737 (
            .O(N__33430),
            .I(n2028));
    LocalMux I__5736 (
            .O(N__33427),
            .I(n2028));
    InMux I__5735 (
            .O(N__33420),
            .I(N__33416));
    CascadeMux I__5734 (
            .O(N__33419),
            .I(N__33413));
    LocalMux I__5733 (
            .O(N__33416),
            .I(N__33409));
    InMux I__5732 (
            .O(N__33413),
            .I(N__33406));
    InMux I__5731 (
            .O(N__33412),
            .I(N__33403));
    Odrv4 I__5730 (
            .O(N__33409),
            .I(n2026));
    LocalMux I__5729 (
            .O(N__33406),
            .I(n2026));
    LocalMux I__5728 (
            .O(N__33403),
            .I(n2026));
    CascadeMux I__5727 (
            .O(N__33396),
            .I(n2025_cascade_));
    InMux I__5726 (
            .O(N__33393),
            .I(N__33389));
    CascadeMux I__5725 (
            .O(N__33392),
            .I(N__33386));
    LocalMux I__5724 (
            .O(N__33389),
            .I(N__33382));
    InMux I__5723 (
            .O(N__33386),
            .I(N__33379));
    InMux I__5722 (
            .O(N__33385),
            .I(N__33376));
    Odrv4 I__5721 (
            .O(N__33382),
            .I(n2027));
    LocalMux I__5720 (
            .O(N__33379),
            .I(n2027));
    LocalMux I__5719 (
            .O(N__33376),
            .I(n2027));
    InMux I__5718 (
            .O(N__33369),
            .I(N__33365));
    CascadeMux I__5717 (
            .O(N__33368),
            .I(N__33362));
    LocalMux I__5716 (
            .O(N__33365),
            .I(N__33359));
    InMux I__5715 (
            .O(N__33362),
            .I(N__33356));
    Span4Mux_h I__5714 (
            .O(N__33359),
            .I(N__33353));
    LocalMux I__5713 (
            .O(N__33356),
            .I(N__33350));
    Odrv4 I__5712 (
            .O(N__33353),
            .I(n2032));
    Odrv4 I__5711 (
            .O(N__33350),
            .I(n2032));
    InMux I__5710 (
            .O(N__33345),
            .I(N__33342));
    LocalMux I__5709 (
            .O(N__33342),
            .I(N__33338));
    CascadeMux I__5708 (
            .O(N__33341),
            .I(N__33335));
    Span4Mux_h I__5707 (
            .O(N__33338),
            .I(N__33331));
    InMux I__5706 (
            .O(N__33335),
            .I(N__33328));
    InMux I__5705 (
            .O(N__33334),
            .I(N__33325));
    Odrv4 I__5704 (
            .O(N__33331),
            .I(n2031));
    LocalMux I__5703 (
            .O(N__33328),
            .I(n2031));
    LocalMux I__5702 (
            .O(N__33325),
            .I(n2031));
    CascadeMux I__5701 (
            .O(N__33318),
            .I(n2032_cascade_));
    CascadeMux I__5700 (
            .O(N__33315),
            .I(N__33311));
    CascadeMux I__5699 (
            .O(N__33314),
            .I(N__33308));
    InMux I__5698 (
            .O(N__33311),
            .I(N__33304));
    InMux I__5697 (
            .O(N__33308),
            .I(N__33301));
    InMux I__5696 (
            .O(N__33307),
            .I(N__33298));
    LocalMux I__5695 (
            .O(N__33304),
            .I(n2022));
    LocalMux I__5694 (
            .O(N__33301),
            .I(n2022));
    LocalMux I__5693 (
            .O(N__33298),
            .I(n2022));
    CascadeMux I__5692 (
            .O(N__33291),
            .I(N__33288));
    InMux I__5691 (
            .O(N__33288),
            .I(N__33283));
    InMux I__5690 (
            .O(N__33287),
            .I(N__33280));
    InMux I__5689 (
            .O(N__33286),
            .I(N__33277));
    LocalMux I__5688 (
            .O(N__33283),
            .I(n2024));
    LocalMux I__5687 (
            .O(N__33280),
            .I(n2024));
    LocalMux I__5686 (
            .O(N__33277),
            .I(n2024));
    CascadeMux I__5685 (
            .O(N__33270),
            .I(N__33265));
    CascadeMux I__5684 (
            .O(N__33269),
            .I(N__33262));
    CascadeMux I__5683 (
            .O(N__33268),
            .I(N__33259));
    InMux I__5682 (
            .O(N__33265),
            .I(N__33256));
    InMux I__5681 (
            .O(N__33262),
            .I(N__33253));
    InMux I__5680 (
            .O(N__33259),
            .I(N__33250));
    LocalMux I__5679 (
            .O(N__33256),
            .I(n2023));
    LocalMux I__5678 (
            .O(N__33253),
            .I(n2023));
    LocalMux I__5677 (
            .O(N__33250),
            .I(n2023));
    InMux I__5676 (
            .O(N__33243),
            .I(N__33240));
    LocalMux I__5675 (
            .O(N__33240),
            .I(n14544));
    InMux I__5674 (
            .O(N__33237),
            .I(N__33234));
    LocalMux I__5673 (
            .O(N__33234),
            .I(n2087));
    CascadeMux I__5672 (
            .O(N__33231),
            .I(n2020_cascade_));
    InMux I__5671 (
            .O(N__33228),
            .I(N__33224));
    InMux I__5670 (
            .O(N__33227),
            .I(N__33221));
    LocalMux I__5669 (
            .O(N__33224),
            .I(N__33217));
    LocalMux I__5668 (
            .O(N__33221),
            .I(N__33214));
    InMux I__5667 (
            .O(N__33220),
            .I(N__33211));
    Span4Mux_h I__5666 (
            .O(N__33217),
            .I(N__33208));
    Span4Mux_h I__5665 (
            .O(N__33214),
            .I(N__33205));
    LocalMux I__5664 (
            .O(N__33211),
            .I(N__33202));
    Odrv4 I__5663 (
            .O(N__33208),
            .I(n2119));
    Odrv4 I__5662 (
            .O(N__33205),
            .I(n2119));
    Odrv4 I__5661 (
            .O(N__33202),
            .I(n2119));
    CascadeMux I__5660 (
            .O(N__33195),
            .I(n14446_cascade_));
    InMux I__5659 (
            .O(N__33192),
            .I(N__33189));
    LocalMux I__5658 (
            .O(N__33189),
            .I(n11985));
    CascadeMux I__5657 (
            .O(N__33186),
            .I(n14450_cascade_));
    CascadeMux I__5656 (
            .O(N__33183),
            .I(n1950_cascade_));
    InMux I__5655 (
            .O(N__33180),
            .I(N__33177));
    LocalMux I__5654 (
            .O(N__33177),
            .I(N__33172));
    InMux I__5653 (
            .O(N__33176),
            .I(N__33167));
    InMux I__5652 (
            .O(N__33175),
            .I(N__33167));
    Odrv12 I__5651 (
            .O(N__33172),
            .I(n2017));
    LocalMux I__5650 (
            .O(N__33167),
            .I(n2017));
    InMux I__5649 (
            .O(N__33162),
            .I(N__33159));
    LocalMux I__5648 (
            .O(N__33159),
            .I(n45_adj_720));
    InMux I__5647 (
            .O(N__33156),
            .I(N__33153));
    LocalMux I__5646 (
            .O(N__33153),
            .I(N__33150));
    IoSpan4Mux I__5645 (
            .O(N__33150),
            .I(N__33147));
    Odrv4 I__5644 (
            .O(N__33147),
            .I(ENCODER0_A_N));
    CascadeMux I__5643 (
            .O(N__33144),
            .I(n1922_cascade_));
    CascadeMux I__5642 (
            .O(N__33141),
            .I(N__33137));
    InMux I__5641 (
            .O(N__33140),
            .I(N__33134));
    InMux I__5640 (
            .O(N__33137),
            .I(N__33131));
    LocalMux I__5639 (
            .O(N__33134),
            .I(N__33128));
    LocalMux I__5638 (
            .O(N__33131),
            .I(n2021));
    Odrv4 I__5637 (
            .O(N__33128),
            .I(n2021));
    InMux I__5636 (
            .O(N__33123),
            .I(N__33120));
    LocalMux I__5635 (
            .O(N__33120),
            .I(n2088));
    CascadeMux I__5634 (
            .O(N__33117),
            .I(n2021_cascade_));
    CascadeMux I__5633 (
            .O(N__33114),
            .I(N__33111));
    InMux I__5632 (
            .O(N__33111),
            .I(N__33107));
    InMux I__5631 (
            .O(N__33110),
            .I(N__33104));
    LocalMux I__5630 (
            .O(N__33107),
            .I(N__33098));
    LocalMux I__5629 (
            .O(N__33104),
            .I(N__33098));
    InMux I__5628 (
            .O(N__33103),
            .I(N__33095));
    Span4Mux_h I__5627 (
            .O(N__33098),
            .I(N__33092));
    LocalMux I__5626 (
            .O(N__33095),
            .I(N__33089));
    Odrv4 I__5625 (
            .O(N__33092),
            .I(n2120));
    Odrv12 I__5624 (
            .O(N__33089),
            .I(n2120));
    CascadeMux I__5623 (
            .O(N__33084),
            .I(N__33080));
    InMux I__5622 (
            .O(N__33083),
            .I(N__33077));
    InMux I__5621 (
            .O(N__33080),
            .I(N__33074));
    LocalMux I__5620 (
            .O(N__33077),
            .I(N__33071));
    LocalMux I__5619 (
            .O(N__33074),
            .I(n2020));
    Odrv4 I__5618 (
            .O(N__33071),
            .I(n2020));
    CascadeMux I__5617 (
            .O(N__33066),
            .I(n14304_cascade_));
    CascadeMux I__5616 (
            .O(N__33063),
            .I(n14306_cascade_));
    InMux I__5615 (
            .O(N__33060),
            .I(N__33057));
    LocalMux I__5614 (
            .O(N__33057),
            .I(n14308));
    InMux I__5613 (
            .O(N__33054),
            .I(N__33051));
    LocalMux I__5612 (
            .O(N__33051),
            .I(n5_adj_704));
    CascadeMux I__5611 (
            .O(N__33048),
            .I(N__33045));
    InMux I__5610 (
            .O(N__33045),
            .I(N__33042));
    LocalMux I__5609 (
            .O(N__33042),
            .I(N__33039));
    Odrv4 I__5608 (
            .O(N__33039),
            .I(n12039));
    CascadeMux I__5607 (
            .O(N__33036),
            .I(n14292_cascade_));
    InMux I__5606 (
            .O(N__33033),
            .I(N__33030));
    LocalMux I__5605 (
            .O(N__33030),
            .I(n14284));
    CascadeMux I__5604 (
            .O(N__33027),
            .I(n14286_cascade_));
    InMux I__5603 (
            .O(N__33024),
            .I(N__33021));
    LocalMux I__5602 (
            .O(N__33021),
            .I(n14288));
    InMux I__5601 (
            .O(N__33018),
            .I(N__33015));
    LocalMux I__5600 (
            .O(N__33015),
            .I(n14294));
    CascadeMux I__5599 (
            .O(N__33012),
            .I(n14296_cascade_));
    InMux I__5598 (
            .O(N__33009),
            .I(N__33006));
    LocalMux I__5597 (
            .O(N__33006),
            .I(n14298));
    CascadeMux I__5596 (
            .O(N__33003),
            .I(n29_adj_717_cascade_));
    InMux I__5595 (
            .O(N__33000),
            .I(N__32997));
    LocalMux I__5594 (
            .O(N__32997),
            .I(N__32994));
    Span4Mux_h I__5593 (
            .O(N__32994),
            .I(N__32991));
    Odrv4 I__5592 (
            .O(N__32991),
            .I(n14270));
    CascadeMux I__5591 (
            .O(N__32988),
            .I(n11941_cascade_));
    InMux I__5590 (
            .O(N__32985),
            .I(N__32982));
    LocalMux I__5589 (
            .O(N__32982),
            .I(n11878));
    InMux I__5588 (
            .O(N__32979),
            .I(N__32976));
    LocalMux I__5587 (
            .O(N__32976),
            .I(n14782));
    InMux I__5586 (
            .O(N__32973),
            .I(N__32970));
    LocalMux I__5585 (
            .O(N__32970),
            .I(n14788));
    CascadeMux I__5584 (
            .O(N__32967),
            .I(n14300_cascade_));
    CascadeMux I__5583 (
            .O(N__32964),
            .I(n14302_cascade_));
    InMux I__5582 (
            .O(N__32961),
            .I(N__32958));
    LocalMux I__5581 (
            .O(N__32958),
            .I(N__32954));
    InMux I__5580 (
            .O(N__32957),
            .I(N__32951));
    Span4Mux_v I__5579 (
            .O(N__32954),
            .I(N__32946));
    LocalMux I__5578 (
            .O(N__32951),
            .I(N__32946));
    Odrv4 I__5577 (
            .O(N__32946),
            .I(n3130));
    CascadeMux I__5576 (
            .O(N__32943),
            .I(N__32940));
    InMux I__5575 (
            .O(N__32940),
            .I(N__32937));
    LocalMux I__5574 (
            .O(N__32937),
            .I(N__32934));
    Span4Mux_h I__5573 (
            .O(N__32934),
            .I(N__32931));
    Odrv4 I__5572 (
            .O(N__32931),
            .I(n3197));
    InMux I__5571 (
            .O(N__32928),
            .I(N__32925));
    LocalMux I__5570 (
            .O(N__32925),
            .I(N__32922));
    Span4Mux_h I__5569 (
            .O(N__32922),
            .I(N__32919));
    Odrv4 I__5568 (
            .O(N__32919),
            .I(n3193));
    CascadeMux I__5567 (
            .O(N__32916),
            .I(N__32912));
    InMux I__5566 (
            .O(N__32915),
            .I(N__32909));
    InMux I__5565 (
            .O(N__32912),
            .I(N__32906));
    LocalMux I__5564 (
            .O(N__32909),
            .I(N__32902));
    LocalMux I__5563 (
            .O(N__32906),
            .I(N__32899));
    InMux I__5562 (
            .O(N__32905),
            .I(N__32896));
    Odrv12 I__5561 (
            .O(N__32902),
            .I(n3126));
    Odrv4 I__5560 (
            .O(N__32899),
            .I(n3126));
    LocalMux I__5559 (
            .O(N__32896),
            .I(n3126));
    InMux I__5558 (
            .O(N__32889),
            .I(N__32886));
    LocalMux I__5557 (
            .O(N__32886),
            .I(N__32883));
    Span4Mux_v I__5556 (
            .O(N__32883),
            .I(N__32880));
    Span4Mux_h I__5555 (
            .O(N__32880),
            .I(N__32877));
    Odrv4 I__5554 (
            .O(N__32877),
            .I(n3201));
    CascadeMux I__5553 (
            .O(N__32874),
            .I(n3233_cascade_));
    CascadeMux I__5552 (
            .O(N__32871),
            .I(n11943_cascade_));
    InMux I__5551 (
            .O(N__32868),
            .I(N__32865));
    LocalMux I__5550 (
            .O(N__32865),
            .I(n13875));
    CascadeMux I__5549 (
            .O(N__32862),
            .I(N__32859));
    InMux I__5548 (
            .O(N__32859),
            .I(N__32855));
    InMux I__5547 (
            .O(N__32858),
            .I(N__32852));
    LocalMux I__5546 (
            .O(N__32855),
            .I(N__32849));
    LocalMux I__5545 (
            .O(N__32852),
            .I(n2515));
    Odrv4 I__5544 (
            .O(N__32849),
            .I(n2515));
    InMux I__5543 (
            .O(N__32844),
            .I(N__32841));
    LocalMux I__5542 (
            .O(N__32841),
            .I(N__32838));
    Span4Mux_h I__5541 (
            .O(N__32838),
            .I(N__32835));
    Odrv4 I__5540 (
            .O(N__32835),
            .I(n2582));
    InMux I__5539 (
            .O(N__32832),
            .I(n12757));
    CascadeMux I__5538 (
            .O(N__32829),
            .I(N__32826));
    InMux I__5537 (
            .O(N__32826),
            .I(N__32823));
    LocalMux I__5536 (
            .O(N__32823),
            .I(N__32819));
    InMux I__5535 (
            .O(N__32822),
            .I(N__32815));
    Span4Mux_v I__5534 (
            .O(N__32819),
            .I(N__32812));
    InMux I__5533 (
            .O(N__32818),
            .I(N__32809));
    LocalMux I__5532 (
            .O(N__32815),
            .I(n2514));
    Odrv4 I__5531 (
            .O(N__32812),
            .I(n2514));
    LocalMux I__5530 (
            .O(N__32809),
            .I(n2514));
    CascadeMux I__5529 (
            .O(N__32802),
            .I(N__32799));
    InMux I__5528 (
            .O(N__32799),
            .I(N__32796));
    LocalMux I__5527 (
            .O(N__32796),
            .I(N__32793));
    Span4Mux_v I__5526 (
            .O(N__32793),
            .I(N__32790));
    Odrv4 I__5525 (
            .O(N__32790),
            .I(n2581));
    InMux I__5524 (
            .O(N__32787),
            .I(n12758));
    CascadeMux I__5523 (
            .O(N__32784),
            .I(N__32781));
    InMux I__5522 (
            .O(N__32781),
            .I(N__32777));
    InMux I__5521 (
            .O(N__32780),
            .I(N__32774));
    LocalMux I__5520 (
            .O(N__32777),
            .I(n2513));
    LocalMux I__5519 (
            .O(N__32774),
            .I(n2513));
    InMux I__5518 (
            .O(N__32769),
            .I(N__32766));
    LocalMux I__5517 (
            .O(N__32766),
            .I(n2580));
    InMux I__5516 (
            .O(N__32763),
            .I(n12759));
    InMux I__5515 (
            .O(N__32760),
            .I(n12760));
    CascadeMux I__5514 (
            .O(N__32757),
            .I(N__32754));
    InMux I__5513 (
            .O(N__32754),
            .I(N__32751));
    LocalMux I__5512 (
            .O(N__32751),
            .I(N__32747));
    InMux I__5511 (
            .O(N__32750),
            .I(N__32744));
    Odrv12 I__5510 (
            .O(N__32747),
            .I(n2511));
    LocalMux I__5509 (
            .O(N__32744),
            .I(n2511));
    InMux I__5508 (
            .O(N__32739),
            .I(n12761));
    CascadeMux I__5507 (
            .O(N__32736),
            .I(N__32733));
    InMux I__5506 (
            .O(N__32733),
            .I(N__32729));
    InMux I__5505 (
            .O(N__32732),
            .I(N__32726));
    LocalMux I__5504 (
            .O(N__32729),
            .I(N__32723));
    LocalMux I__5503 (
            .O(N__32726),
            .I(N__32717));
    Span4Mux_v I__5502 (
            .O(N__32723),
            .I(N__32717));
    InMux I__5501 (
            .O(N__32722),
            .I(N__32714));
    Span4Mux_v I__5500 (
            .O(N__32717),
            .I(N__32709));
    LocalMux I__5499 (
            .O(N__32714),
            .I(N__32709));
    Span4Mux_h I__5498 (
            .O(N__32709),
            .I(N__32706));
    Odrv4 I__5497 (
            .O(N__32706),
            .I(n2610));
    InMux I__5496 (
            .O(N__32703),
            .I(N__32699));
    CascadeMux I__5495 (
            .O(N__32702),
            .I(N__32696));
    LocalMux I__5494 (
            .O(N__32699),
            .I(N__32692));
    InMux I__5493 (
            .O(N__32696),
            .I(N__32689));
    InMux I__5492 (
            .O(N__32695),
            .I(N__32686));
    Span4Mux_v I__5491 (
            .O(N__32692),
            .I(N__32679));
    LocalMux I__5490 (
            .O(N__32689),
            .I(N__32679));
    LocalMux I__5489 (
            .O(N__32686),
            .I(N__32679));
    Span4Mux_v I__5488 (
            .O(N__32679),
            .I(N__32676));
    Odrv4 I__5487 (
            .O(N__32676),
            .I(n2418));
    CascadeMux I__5486 (
            .O(N__32673),
            .I(N__32670));
    InMux I__5485 (
            .O(N__32670),
            .I(N__32667));
    LocalMux I__5484 (
            .O(N__32667),
            .I(N__32664));
    Odrv12 I__5483 (
            .O(N__32664),
            .I(n2485));
    InMux I__5482 (
            .O(N__32661),
            .I(N__32658));
    LocalMux I__5481 (
            .O(N__32658),
            .I(N__32654));
    CascadeMux I__5480 (
            .O(N__32657),
            .I(N__32651));
    Span4Mux_v I__5479 (
            .O(N__32654),
            .I(N__32648));
    InMux I__5478 (
            .O(N__32651),
            .I(N__32645));
    Span4Mux_v I__5477 (
            .O(N__32648),
            .I(N__32642));
    LocalMux I__5476 (
            .O(N__32645),
            .I(n2517));
    Odrv4 I__5475 (
            .O(N__32642),
            .I(n2517));
    InMux I__5474 (
            .O(N__32637),
            .I(N__32634));
    LocalMux I__5473 (
            .O(N__32634),
            .I(n2584));
    CascadeMux I__5472 (
            .O(N__32631),
            .I(n2517_cascade_));
    InMux I__5471 (
            .O(N__32628),
            .I(N__32625));
    LocalMux I__5470 (
            .O(N__32625),
            .I(N__32621));
    InMux I__5469 (
            .O(N__32624),
            .I(N__32618));
    Span4Mux_h I__5468 (
            .O(N__32621),
            .I(N__32614));
    LocalMux I__5467 (
            .O(N__32618),
            .I(N__32611));
    InMux I__5466 (
            .O(N__32617),
            .I(N__32608));
    Span4Mux_v I__5465 (
            .O(N__32614),
            .I(N__32605));
    Span4Mux_v I__5464 (
            .O(N__32611),
            .I(N__32600));
    LocalMux I__5463 (
            .O(N__32608),
            .I(N__32600));
    Span4Mux_v I__5462 (
            .O(N__32605),
            .I(N__32595));
    Span4Mux_h I__5461 (
            .O(N__32600),
            .I(N__32595));
    Odrv4 I__5460 (
            .O(N__32595),
            .I(n2616));
    InMux I__5459 (
            .O(N__32592),
            .I(N__32588));
    InMux I__5458 (
            .O(N__32591),
            .I(N__32585));
    LocalMux I__5457 (
            .O(N__32588),
            .I(N__32580));
    LocalMux I__5456 (
            .O(N__32585),
            .I(N__32580));
    Span4Mux_v I__5455 (
            .O(N__32580),
            .I(N__32576));
    InMux I__5454 (
            .O(N__32579),
            .I(N__32573));
    Odrv4 I__5453 (
            .O(N__32576),
            .I(n2512));
    LocalMux I__5452 (
            .O(N__32573),
            .I(n2512));
    CascadeMux I__5451 (
            .O(N__32568),
            .I(N__32565));
    InMux I__5450 (
            .O(N__32565),
            .I(N__32562));
    LocalMux I__5449 (
            .O(N__32562),
            .I(n2579));
    InMux I__5448 (
            .O(N__32559),
            .I(N__32556));
    LocalMux I__5447 (
            .O(N__32556),
            .I(N__32552));
    InMux I__5446 (
            .O(N__32555),
            .I(N__32549));
    Span4Mux_h I__5445 (
            .O(N__32552),
            .I(N__32545));
    LocalMux I__5444 (
            .O(N__32549),
            .I(N__32542));
    InMux I__5443 (
            .O(N__32548),
            .I(N__32539));
    Span4Mux_v I__5442 (
            .O(N__32545),
            .I(N__32536));
    Span4Mux_v I__5441 (
            .O(N__32542),
            .I(N__32531));
    LocalMux I__5440 (
            .O(N__32539),
            .I(N__32531));
    Span4Mux_v I__5439 (
            .O(N__32536),
            .I(N__32526));
    Span4Mux_h I__5438 (
            .O(N__32531),
            .I(N__32526));
    Odrv4 I__5437 (
            .O(N__32526),
            .I(n2611));
    InMux I__5436 (
            .O(N__32523),
            .I(n12748));
    CascadeMux I__5435 (
            .O(N__32520),
            .I(N__32517));
    InMux I__5434 (
            .O(N__32517),
            .I(N__32514));
    LocalMux I__5433 (
            .O(N__32514),
            .I(N__32510));
    InMux I__5432 (
            .O(N__32513),
            .I(N__32507));
    Span4Mux_h I__5431 (
            .O(N__32510),
            .I(N__32504));
    LocalMux I__5430 (
            .O(N__32507),
            .I(n2523));
    Odrv4 I__5429 (
            .O(N__32504),
            .I(n2523));
    InMux I__5428 (
            .O(N__32499),
            .I(N__32496));
    LocalMux I__5427 (
            .O(N__32496),
            .I(N__32493));
    Span4Mux_h I__5426 (
            .O(N__32493),
            .I(N__32490));
    Odrv4 I__5425 (
            .O(N__32490),
            .I(n2590));
    InMux I__5424 (
            .O(N__32487),
            .I(n12749));
    CascadeMux I__5423 (
            .O(N__32484),
            .I(N__32481));
    InMux I__5422 (
            .O(N__32481),
            .I(N__32478));
    LocalMux I__5421 (
            .O(N__32478),
            .I(N__32475));
    Span4Mux_h I__5420 (
            .O(N__32475),
            .I(N__32472));
    Odrv4 I__5419 (
            .O(N__32472),
            .I(n2589));
    InMux I__5418 (
            .O(N__32469),
            .I(n12750));
    InMux I__5417 (
            .O(N__32466),
            .I(N__32463));
    LocalMux I__5416 (
            .O(N__32463),
            .I(N__32460));
    Odrv4 I__5415 (
            .O(N__32460),
            .I(n2588));
    InMux I__5414 (
            .O(N__32457),
            .I(n12751));
    CascadeMux I__5413 (
            .O(N__32454),
            .I(N__32451));
    InMux I__5412 (
            .O(N__32451),
            .I(N__32447));
    InMux I__5411 (
            .O(N__32450),
            .I(N__32443));
    LocalMux I__5410 (
            .O(N__32447),
            .I(N__32440));
    InMux I__5409 (
            .O(N__32446),
            .I(N__32437));
    LocalMux I__5408 (
            .O(N__32443),
            .I(n2520));
    Odrv4 I__5407 (
            .O(N__32440),
            .I(n2520));
    LocalMux I__5406 (
            .O(N__32437),
            .I(n2520));
    InMux I__5405 (
            .O(N__32430),
            .I(N__32427));
    LocalMux I__5404 (
            .O(N__32427),
            .I(N__32424));
    Span4Mux_h I__5403 (
            .O(N__32424),
            .I(N__32421));
    Odrv4 I__5402 (
            .O(N__32421),
            .I(n2587));
    InMux I__5401 (
            .O(N__32418),
            .I(n12752));
    CascadeMux I__5400 (
            .O(N__32415),
            .I(N__32412));
    InMux I__5399 (
            .O(N__32412),
            .I(N__32409));
    LocalMux I__5398 (
            .O(N__32409),
            .I(N__32405));
    InMux I__5397 (
            .O(N__32408),
            .I(N__32401));
    Span4Mux_v I__5396 (
            .O(N__32405),
            .I(N__32398));
    InMux I__5395 (
            .O(N__32404),
            .I(N__32395));
    LocalMux I__5394 (
            .O(N__32401),
            .I(n2519));
    Odrv4 I__5393 (
            .O(N__32398),
            .I(n2519));
    LocalMux I__5392 (
            .O(N__32395),
            .I(n2519));
    CascadeMux I__5391 (
            .O(N__32388),
            .I(N__32385));
    InMux I__5390 (
            .O(N__32385),
            .I(N__32382));
    LocalMux I__5389 (
            .O(N__32382),
            .I(N__32379));
    Span4Mux_v I__5388 (
            .O(N__32379),
            .I(N__32376));
    Odrv4 I__5387 (
            .O(N__32376),
            .I(n2586));
    InMux I__5386 (
            .O(N__32373),
            .I(n12753));
    CascadeMux I__5385 (
            .O(N__32370),
            .I(N__32367));
    InMux I__5384 (
            .O(N__32367),
            .I(N__32364));
    LocalMux I__5383 (
            .O(N__32364),
            .I(N__32361));
    Span4Mux_h I__5382 (
            .O(N__32361),
            .I(N__32358));
    Odrv4 I__5381 (
            .O(N__32358),
            .I(n2585));
    InMux I__5380 (
            .O(N__32355),
            .I(bfn_6_26_0_));
    InMux I__5379 (
            .O(N__32352),
            .I(n12755));
    InMux I__5378 (
            .O(N__32349),
            .I(N__32345));
    CascadeMux I__5377 (
            .O(N__32348),
            .I(N__32342));
    LocalMux I__5376 (
            .O(N__32345),
            .I(N__32339));
    InMux I__5375 (
            .O(N__32342),
            .I(N__32336));
    Span4Mux_v I__5374 (
            .O(N__32339),
            .I(N__32331));
    LocalMux I__5373 (
            .O(N__32336),
            .I(N__32331));
    Span4Mux_v I__5372 (
            .O(N__32331),
            .I(N__32327));
    InMux I__5371 (
            .O(N__32330),
            .I(N__32324));
    Odrv4 I__5370 (
            .O(N__32327),
            .I(n2516));
    LocalMux I__5369 (
            .O(N__32324),
            .I(n2516));
    InMux I__5368 (
            .O(N__32319),
            .I(N__32316));
    LocalMux I__5367 (
            .O(N__32316),
            .I(n2583));
    InMux I__5366 (
            .O(N__32313),
            .I(n12756));
    CascadeMux I__5365 (
            .O(N__32310),
            .I(N__32307));
    InMux I__5364 (
            .O(N__32307),
            .I(N__32302));
    InMux I__5363 (
            .O(N__32306),
            .I(N__32299));
    InMux I__5362 (
            .O(N__32305),
            .I(N__32296));
    LocalMux I__5361 (
            .O(N__32302),
            .I(N__32293));
    LocalMux I__5360 (
            .O(N__32299),
            .I(N__32288));
    LocalMux I__5359 (
            .O(N__32296),
            .I(N__32288));
    Odrv4 I__5358 (
            .O(N__32293),
            .I(n2531));
    Odrv4 I__5357 (
            .O(N__32288),
            .I(n2531));
    InMux I__5356 (
            .O(N__32283),
            .I(N__32280));
    LocalMux I__5355 (
            .O(N__32280),
            .I(n2598));
    InMux I__5354 (
            .O(N__32277),
            .I(n12741));
    CascadeMux I__5353 (
            .O(N__32274),
            .I(N__32271));
    InMux I__5352 (
            .O(N__32271),
            .I(N__32267));
    CascadeMux I__5351 (
            .O(N__32270),
            .I(N__32264));
    LocalMux I__5350 (
            .O(N__32267),
            .I(N__32261));
    InMux I__5349 (
            .O(N__32264),
            .I(N__32258));
    Odrv4 I__5348 (
            .O(N__32261),
            .I(n2530));
    LocalMux I__5347 (
            .O(N__32258),
            .I(n2530));
    InMux I__5346 (
            .O(N__32253),
            .I(N__32250));
    LocalMux I__5345 (
            .O(N__32250),
            .I(n2597));
    InMux I__5344 (
            .O(N__32247),
            .I(n12742));
    InMux I__5343 (
            .O(N__32244),
            .I(N__32241));
    LocalMux I__5342 (
            .O(N__32241),
            .I(N__32237));
    CascadeMux I__5341 (
            .O(N__32240),
            .I(N__32234));
    Span4Mux_h I__5340 (
            .O(N__32237),
            .I(N__32230));
    InMux I__5339 (
            .O(N__32234),
            .I(N__32227));
    InMux I__5338 (
            .O(N__32233),
            .I(N__32224));
    Odrv4 I__5337 (
            .O(N__32230),
            .I(n2529));
    LocalMux I__5336 (
            .O(N__32227),
            .I(n2529));
    LocalMux I__5335 (
            .O(N__32224),
            .I(n2529));
    CascadeMux I__5334 (
            .O(N__32217),
            .I(N__32214));
    InMux I__5333 (
            .O(N__32214),
            .I(N__32211));
    LocalMux I__5332 (
            .O(N__32211),
            .I(N__32208));
    Span4Mux_v I__5331 (
            .O(N__32208),
            .I(N__32205));
    Odrv4 I__5330 (
            .O(N__32205),
            .I(n2596));
    InMux I__5329 (
            .O(N__32202),
            .I(n12743));
    CascadeMux I__5328 (
            .O(N__32199),
            .I(N__32196));
    InMux I__5327 (
            .O(N__32196),
            .I(N__32193));
    LocalMux I__5326 (
            .O(N__32193),
            .I(N__32190));
    Span4Mux_h I__5325 (
            .O(N__32190),
            .I(N__32186));
    InMux I__5324 (
            .O(N__32189),
            .I(N__32183));
    Odrv4 I__5323 (
            .O(N__32186),
            .I(n2528));
    LocalMux I__5322 (
            .O(N__32183),
            .I(n2528));
    InMux I__5321 (
            .O(N__32178),
            .I(N__32175));
    LocalMux I__5320 (
            .O(N__32175),
            .I(N__32172));
    Odrv4 I__5319 (
            .O(N__32172),
            .I(n2595));
    InMux I__5318 (
            .O(N__32169),
            .I(n12744));
    CascadeMux I__5317 (
            .O(N__32166),
            .I(N__32163));
    InMux I__5316 (
            .O(N__32163),
            .I(N__32160));
    LocalMux I__5315 (
            .O(N__32160),
            .I(N__32157));
    Span4Mux_h I__5314 (
            .O(N__32157),
            .I(N__32153));
    InMux I__5313 (
            .O(N__32156),
            .I(N__32150));
    Odrv4 I__5312 (
            .O(N__32153),
            .I(n2527));
    LocalMux I__5311 (
            .O(N__32150),
            .I(n2527));
    InMux I__5310 (
            .O(N__32145),
            .I(N__32142));
    LocalMux I__5309 (
            .O(N__32142),
            .I(N__32139));
    Span4Mux_h I__5308 (
            .O(N__32139),
            .I(N__32136));
    Odrv4 I__5307 (
            .O(N__32136),
            .I(n2594));
    InMux I__5306 (
            .O(N__32133),
            .I(n12745));
    CascadeMux I__5305 (
            .O(N__32130),
            .I(N__32127));
    InMux I__5304 (
            .O(N__32127),
            .I(N__32124));
    LocalMux I__5303 (
            .O(N__32124),
            .I(N__32121));
    Span4Mux_v I__5302 (
            .O(N__32121),
            .I(N__32117));
    InMux I__5301 (
            .O(N__32120),
            .I(N__32114));
    Odrv4 I__5300 (
            .O(N__32117),
            .I(n2526));
    LocalMux I__5299 (
            .O(N__32114),
            .I(n2526));
    InMux I__5298 (
            .O(N__32109),
            .I(N__32106));
    LocalMux I__5297 (
            .O(N__32106),
            .I(N__32103));
    Span4Mux_h I__5296 (
            .O(N__32103),
            .I(N__32100));
    Odrv4 I__5295 (
            .O(N__32100),
            .I(n2593));
    InMux I__5294 (
            .O(N__32097),
            .I(bfn_6_25_0_));
    InMux I__5293 (
            .O(N__32094),
            .I(n12747));
    InMux I__5292 (
            .O(N__32091),
            .I(N__32087));
    CascadeMux I__5291 (
            .O(N__32090),
            .I(N__32084));
    LocalMux I__5290 (
            .O(N__32087),
            .I(N__32081));
    InMux I__5289 (
            .O(N__32084),
            .I(N__32078));
    Span4Mux_v I__5288 (
            .O(N__32081),
            .I(N__32075));
    LocalMux I__5287 (
            .O(N__32078),
            .I(n2524));
    Odrv4 I__5286 (
            .O(N__32075),
            .I(n2524));
    InMux I__5285 (
            .O(N__32070),
            .I(N__32067));
    LocalMux I__5284 (
            .O(N__32067),
            .I(N__32064));
    Span4Mux_h I__5283 (
            .O(N__32064),
            .I(N__32061));
    Odrv4 I__5282 (
            .O(N__32061),
            .I(n2591));
    InMux I__5281 (
            .O(N__32058),
            .I(n12734));
    CascadeMux I__5280 (
            .O(N__32055),
            .I(N__32050));
    InMux I__5279 (
            .O(N__32054),
            .I(N__32047));
    InMux I__5278 (
            .O(N__32053),
            .I(N__32042));
    InMux I__5277 (
            .O(N__32050),
            .I(N__32042));
    LocalMux I__5276 (
            .O(N__32047),
            .I(N__32037));
    LocalMux I__5275 (
            .O(N__32042),
            .I(N__32037));
    Span4Mux_h I__5274 (
            .O(N__32037),
            .I(N__32034));
    Odrv4 I__5273 (
            .O(N__32034),
            .I(n2415));
    InMux I__5272 (
            .O(N__32031),
            .I(N__32028));
    LocalMux I__5271 (
            .O(N__32028),
            .I(n2482));
    InMux I__5270 (
            .O(N__32025),
            .I(n12735));
    CascadeMux I__5269 (
            .O(N__32022),
            .I(N__32019));
    InMux I__5268 (
            .O(N__32019),
            .I(N__32016));
    LocalMux I__5267 (
            .O(N__32016),
            .I(N__32012));
    InMux I__5266 (
            .O(N__32015),
            .I(N__32009));
    Span4Mux_v I__5265 (
            .O(N__32012),
            .I(N__32003));
    LocalMux I__5264 (
            .O(N__32009),
            .I(N__32003));
    InMux I__5263 (
            .O(N__32008),
            .I(N__32000));
    Span4Mux_h I__5262 (
            .O(N__32003),
            .I(N__31995));
    LocalMux I__5261 (
            .O(N__32000),
            .I(N__31995));
    Odrv4 I__5260 (
            .O(N__31995),
            .I(n2414));
    InMux I__5259 (
            .O(N__31992),
            .I(N__31989));
    LocalMux I__5258 (
            .O(N__31989),
            .I(N__31986));
    Odrv4 I__5257 (
            .O(N__31986),
            .I(n2481));
    InMux I__5256 (
            .O(N__31983),
            .I(n12736));
    InMux I__5255 (
            .O(N__31980),
            .I(N__31976));
    InMux I__5254 (
            .O(N__31979),
            .I(N__31973));
    LocalMux I__5253 (
            .O(N__31976),
            .I(N__31969));
    LocalMux I__5252 (
            .O(N__31973),
            .I(N__31966));
    InMux I__5251 (
            .O(N__31972),
            .I(N__31963));
    Span4Mux_v I__5250 (
            .O(N__31969),
            .I(N__31956));
    Span4Mux_h I__5249 (
            .O(N__31966),
            .I(N__31956));
    LocalMux I__5248 (
            .O(N__31963),
            .I(N__31956));
    Odrv4 I__5247 (
            .O(N__31956),
            .I(n2413));
    InMux I__5246 (
            .O(N__31953),
            .I(N__31950));
    LocalMux I__5245 (
            .O(N__31950),
            .I(n2480));
    InMux I__5244 (
            .O(N__31947),
            .I(n12737));
    InMux I__5243 (
            .O(N__31944),
            .I(N__31941));
    LocalMux I__5242 (
            .O(N__31941),
            .I(N__31937));
    InMux I__5241 (
            .O(N__31940),
            .I(N__31934));
    Span4Mux_h I__5240 (
            .O(N__31937),
            .I(N__31929));
    LocalMux I__5239 (
            .O(N__31934),
            .I(N__31929));
    Span4Mux_h I__5238 (
            .O(N__31929),
            .I(N__31926));
    Odrv4 I__5237 (
            .O(N__31926),
            .I(n2412));
    InMux I__5236 (
            .O(N__31923),
            .I(n12738));
    InMux I__5235 (
            .O(N__31920),
            .I(N__31917));
    LocalMux I__5234 (
            .O(N__31917),
            .I(N__31913));
    CascadeMux I__5233 (
            .O(N__31916),
            .I(N__31910));
    Span4Mux_v I__5232 (
            .O(N__31913),
            .I(N__31906));
    InMux I__5231 (
            .O(N__31910),
            .I(N__31903));
    InMux I__5230 (
            .O(N__31909),
            .I(N__31900));
    Odrv4 I__5229 (
            .O(N__31906),
            .I(n2433));
    LocalMux I__5228 (
            .O(N__31903),
            .I(n2433));
    LocalMux I__5227 (
            .O(N__31900),
            .I(n2433));
    CascadeMux I__5226 (
            .O(N__31893),
            .I(N__31890));
    InMux I__5225 (
            .O(N__31890),
            .I(N__31887));
    LocalMux I__5224 (
            .O(N__31887),
            .I(N__31884));
    Odrv4 I__5223 (
            .O(N__31884),
            .I(n2500));
    InMux I__5222 (
            .O(N__31881),
            .I(N__31878));
    LocalMux I__5221 (
            .O(N__31878),
            .I(N__31875));
    Span4Mux_v I__5220 (
            .O(N__31875),
            .I(N__31872));
    Odrv4 I__5219 (
            .O(N__31872),
            .I(n2601));
    InMux I__5218 (
            .O(N__31869),
            .I(bfn_6_24_0_));
    CascadeMux I__5217 (
            .O(N__31866),
            .I(N__31862));
    InMux I__5216 (
            .O(N__31865),
            .I(N__31859));
    InMux I__5215 (
            .O(N__31862),
            .I(N__31856));
    LocalMux I__5214 (
            .O(N__31859),
            .I(n2533));
    LocalMux I__5213 (
            .O(N__31856),
            .I(n2533));
    CascadeMux I__5212 (
            .O(N__31851),
            .I(N__31848));
    InMux I__5211 (
            .O(N__31848),
            .I(N__31845));
    LocalMux I__5210 (
            .O(N__31845),
            .I(n2600));
    InMux I__5209 (
            .O(N__31842),
            .I(n12739));
    CascadeMux I__5208 (
            .O(N__31839),
            .I(N__31836));
    InMux I__5207 (
            .O(N__31836),
            .I(N__31831));
    InMux I__5206 (
            .O(N__31835),
            .I(N__31826));
    InMux I__5205 (
            .O(N__31834),
            .I(N__31826));
    LocalMux I__5204 (
            .O(N__31831),
            .I(n2532));
    LocalMux I__5203 (
            .O(N__31826),
            .I(n2532));
    InMux I__5202 (
            .O(N__31821),
            .I(N__31818));
    LocalMux I__5201 (
            .O(N__31818),
            .I(n2599));
    InMux I__5200 (
            .O(N__31815),
            .I(n12740));
    CascadeMux I__5199 (
            .O(N__31812),
            .I(N__31809));
    InMux I__5198 (
            .O(N__31809),
            .I(N__31805));
    InMux I__5197 (
            .O(N__31808),
            .I(N__31802));
    LocalMux I__5196 (
            .O(N__31805),
            .I(N__31799));
    LocalMux I__5195 (
            .O(N__31802),
            .I(N__31793));
    Span4Mux_h I__5194 (
            .O(N__31799),
            .I(N__31793));
    InMux I__5193 (
            .O(N__31798),
            .I(N__31790));
    Odrv4 I__5192 (
            .O(N__31793),
            .I(n2424));
    LocalMux I__5191 (
            .O(N__31790),
            .I(n2424));
    CascadeMux I__5190 (
            .O(N__31785),
            .I(N__31782));
    InMux I__5189 (
            .O(N__31782),
            .I(N__31779));
    LocalMux I__5188 (
            .O(N__31779),
            .I(N__31776));
    Odrv4 I__5187 (
            .O(N__31776),
            .I(n2491));
    InMux I__5186 (
            .O(N__31773),
            .I(n12726));
    InMux I__5185 (
            .O(N__31770),
            .I(n12727));
    InMux I__5184 (
            .O(N__31767),
            .I(n12728));
    CascadeMux I__5183 (
            .O(N__31764),
            .I(N__31761));
    InMux I__5182 (
            .O(N__31761),
            .I(N__31757));
    InMux I__5181 (
            .O(N__31760),
            .I(N__31754));
    LocalMux I__5180 (
            .O(N__31757),
            .I(N__31750));
    LocalMux I__5179 (
            .O(N__31754),
            .I(N__31747));
    InMux I__5178 (
            .O(N__31753),
            .I(N__31744));
    Odrv12 I__5177 (
            .O(N__31750),
            .I(n2421));
    Odrv4 I__5176 (
            .O(N__31747),
            .I(n2421));
    LocalMux I__5175 (
            .O(N__31744),
            .I(n2421));
    InMux I__5174 (
            .O(N__31737),
            .I(N__31734));
    LocalMux I__5173 (
            .O(N__31734),
            .I(n2488));
    InMux I__5172 (
            .O(N__31731),
            .I(n12729));
    CascadeMux I__5171 (
            .O(N__31728),
            .I(N__31724));
    CascadeMux I__5170 (
            .O(N__31727),
            .I(N__31721));
    InMux I__5169 (
            .O(N__31724),
            .I(N__31718));
    InMux I__5168 (
            .O(N__31721),
            .I(N__31715));
    LocalMux I__5167 (
            .O(N__31718),
            .I(n2420));
    LocalMux I__5166 (
            .O(N__31715),
            .I(n2420));
    InMux I__5165 (
            .O(N__31710),
            .I(N__31707));
    LocalMux I__5164 (
            .O(N__31707),
            .I(N__31704));
    Odrv4 I__5163 (
            .O(N__31704),
            .I(n2487));
    InMux I__5162 (
            .O(N__31701),
            .I(n12730));
    InMux I__5161 (
            .O(N__31698),
            .I(n12731));
    InMux I__5160 (
            .O(N__31695),
            .I(bfn_6_23_0_));
    InMux I__5159 (
            .O(N__31692),
            .I(N__31688));
    InMux I__5158 (
            .O(N__31691),
            .I(N__31685));
    LocalMux I__5157 (
            .O(N__31688),
            .I(n2417));
    LocalMux I__5156 (
            .O(N__31685),
            .I(n2417));
    InMux I__5155 (
            .O(N__31680),
            .I(N__31677));
    LocalMux I__5154 (
            .O(N__31677),
            .I(n2484));
    InMux I__5153 (
            .O(N__31674),
            .I(n12733));
    InMux I__5152 (
            .O(N__31671),
            .I(N__31668));
    LocalMux I__5151 (
            .O(N__31668),
            .I(N__31663));
    InMux I__5150 (
            .O(N__31667),
            .I(N__31660));
    InMux I__5149 (
            .O(N__31666),
            .I(N__31657));
    Odrv4 I__5148 (
            .O(N__31663),
            .I(n2416));
    LocalMux I__5147 (
            .O(N__31660),
            .I(n2416));
    LocalMux I__5146 (
            .O(N__31657),
            .I(n2416));
    CascadeMux I__5145 (
            .O(N__31650),
            .I(N__31647));
    InMux I__5144 (
            .O(N__31647),
            .I(N__31644));
    LocalMux I__5143 (
            .O(N__31644),
            .I(n2483));
    CascadeMux I__5142 (
            .O(N__31641),
            .I(N__31637));
    CascadeMux I__5141 (
            .O(N__31640),
            .I(N__31634));
    InMux I__5140 (
            .O(N__31637),
            .I(N__31631));
    InMux I__5139 (
            .O(N__31634),
            .I(N__31628));
    LocalMux I__5138 (
            .O(N__31631),
            .I(n2432));
    LocalMux I__5137 (
            .O(N__31628),
            .I(n2432));
    InMux I__5136 (
            .O(N__31623),
            .I(N__31620));
    LocalMux I__5135 (
            .O(N__31620),
            .I(N__31617));
    Odrv4 I__5134 (
            .O(N__31617),
            .I(n2499));
    InMux I__5133 (
            .O(N__31614),
            .I(n12718));
    InMux I__5132 (
            .O(N__31611),
            .I(N__31607));
    CascadeMux I__5131 (
            .O(N__31610),
            .I(N__31603));
    LocalMux I__5130 (
            .O(N__31607),
            .I(N__31600));
    InMux I__5129 (
            .O(N__31606),
            .I(N__31597));
    InMux I__5128 (
            .O(N__31603),
            .I(N__31594));
    Odrv4 I__5127 (
            .O(N__31600),
            .I(n2431));
    LocalMux I__5126 (
            .O(N__31597),
            .I(n2431));
    LocalMux I__5125 (
            .O(N__31594),
            .I(n2431));
    CascadeMux I__5124 (
            .O(N__31587),
            .I(N__31584));
    InMux I__5123 (
            .O(N__31584),
            .I(N__31581));
    LocalMux I__5122 (
            .O(N__31581),
            .I(N__31578));
    Odrv4 I__5121 (
            .O(N__31578),
            .I(n2498));
    InMux I__5120 (
            .O(N__31575),
            .I(n12719));
    InMux I__5119 (
            .O(N__31572),
            .I(N__31568));
    CascadeMux I__5118 (
            .O(N__31571),
            .I(N__31565));
    LocalMux I__5117 (
            .O(N__31568),
            .I(N__31562));
    InMux I__5116 (
            .O(N__31565),
            .I(N__31559));
    Odrv12 I__5115 (
            .O(N__31562),
            .I(n2430));
    LocalMux I__5114 (
            .O(N__31559),
            .I(n2430));
    InMux I__5113 (
            .O(N__31554),
            .I(N__31551));
    LocalMux I__5112 (
            .O(N__31551),
            .I(N__31548));
    Odrv4 I__5111 (
            .O(N__31548),
            .I(n2497));
    InMux I__5110 (
            .O(N__31545),
            .I(n12720));
    CascadeMux I__5109 (
            .O(N__31542),
            .I(N__31539));
    InMux I__5108 (
            .O(N__31539),
            .I(N__31535));
    CascadeMux I__5107 (
            .O(N__31538),
            .I(N__31532));
    LocalMux I__5106 (
            .O(N__31535),
            .I(N__31528));
    InMux I__5105 (
            .O(N__31532),
            .I(N__31525));
    InMux I__5104 (
            .O(N__31531),
            .I(N__31522));
    Odrv4 I__5103 (
            .O(N__31528),
            .I(n2429));
    LocalMux I__5102 (
            .O(N__31525),
            .I(n2429));
    LocalMux I__5101 (
            .O(N__31522),
            .I(n2429));
    InMux I__5100 (
            .O(N__31515),
            .I(N__31512));
    LocalMux I__5099 (
            .O(N__31512),
            .I(n2496));
    InMux I__5098 (
            .O(N__31509),
            .I(n12721));
    CascadeMux I__5097 (
            .O(N__31506),
            .I(N__31503));
    InMux I__5096 (
            .O(N__31503),
            .I(N__31499));
    InMux I__5095 (
            .O(N__31502),
            .I(N__31495));
    LocalMux I__5094 (
            .O(N__31499),
            .I(N__31492));
    InMux I__5093 (
            .O(N__31498),
            .I(N__31489));
    LocalMux I__5092 (
            .O(N__31495),
            .I(n2428));
    Odrv4 I__5091 (
            .O(N__31492),
            .I(n2428));
    LocalMux I__5090 (
            .O(N__31489),
            .I(n2428));
    CascadeMux I__5089 (
            .O(N__31482),
            .I(N__31479));
    InMux I__5088 (
            .O(N__31479),
            .I(N__31476));
    LocalMux I__5087 (
            .O(N__31476),
            .I(N__31473));
    Span4Mux_h I__5086 (
            .O(N__31473),
            .I(N__31470));
    Odrv4 I__5085 (
            .O(N__31470),
            .I(n2495));
    InMux I__5084 (
            .O(N__31467),
            .I(n12722));
    InMux I__5083 (
            .O(N__31464),
            .I(N__31460));
    InMux I__5082 (
            .O(N__31463),
            .I(N__31457));
    LocalMux I__5081 (
            .O(N__31460),
            .I(N__31452));
    LocalMux I__5080 (
            .O(N__31457),
            .I(N__31452));
    Odrv4 I__5079 (
            .O(N__31452),
            .I(n2427));
    CascadeMux I__5078 (
            .O(N__31449),
            .I(N__31446));
    InMux I__5077 (
            .O(N__31446),
            .I(N__31443));
    LocalMux I__5076 (
            .O(N__31443),
            .I(N__31440));
    Odrv4 I__5075 (
            .O(N__31440),
            .I(n2494));
    InMux I__5074 (
            .O(N__31437),
            .I(n12723));
    InMux I__5073 (
            .O(N__31434),
            .I(bfn_6_22_0_));
    CascadeMux I__5072 (
            .O(N__31431),
            .I(N__31427));
    InMux I__5071 (
            .O(N__31430),
            .I(N__31424));
    InMux I__5070 (
            .O(N__31427),
            .I(N__31421));
    LocalMux I__5069 (
            .O(N__31424),
            .I(N__31417));
    LocalMux I__5068 (
            .O(N__31421),
            .I(N__31414));
    InMux I__5067 (
            .O(N__31420),
            .I(N__31411));
    Odrv4 I__5066 (
            .O(N__31417),
            .I(n2425));
    Odrv4 I__5065 (
            .O(N__31414),
            .I(n2425));
    LocalMux I__5064 (
            .O(N__31411),
            .I(n2425));
    InMux I__5063 (
            .O(N__31404),
            .I(N__31401));
    LocalMux I__5062 (
            .O(N__31401),
            .I(N__31398));
    Odrv4 I__5061 (
            .O(N__31398),
            .I(n2492));
    InMux I__5060 (
            .O(N__31395),
            .I(n12725));
    CascadeMux I__5059 (
            .O(N__31392),
            .I(n14558_cascade_));
    InMux I__5058 (
            .O(N__31389),
            .I(N__31386));
    LocalMux I__5057 (
            .O(N__31386),
            .I(N__31383));
    Odrv4 I__5056 (
            .O(N__31383),
            .I(n2101));
    CascadeMux I__5055 (
            .O(N__31380),
            .I(n2049_cascade_));
    InMux I__5054 (
            .O(N__31377),
            .I(N__31371));
    InMux I__5053 (
            .O(N__31376),
            .I(N__31371));
    LocalMux I__5052 (
            .O(N__31371),
            .I(N__31368));
    Odrv4 I__5051 (
            .O(N__31368),
            .I(n2018));
    InMux I__5050 (
            .O(N__31365),
            .I(N__31362));
    LocalMux I__5049 (
            .O(N__31362),
            .I(n2085));
    CascadeMux I__5048 (
            .O(N__31359),
            .I(n2018_cascade_));
    InMux I__5047 (
            .O(N__31356),
            .I(N__31352));
    InMux I__5046 (
            .O(N__31355),
            .I(N__31349));
    LocalMux I__5045 (
            .O(N__31352),
            .I(N__31346));
    LocalMux I__5044 (
            .O(N__31349),
            .I(N__31342));
    Span4Mux_v I__5043 (
            .O(N__31346),
            .I(N__31339));
    InMux I__5042 (
            .O(N__31345),
            .I(N__31336));
    Span4Mux_h I__5041 (
            .O(N__31342),
            .I(N__31333));
    Span4Mux_h I__5040 (
            .O(N__31339),
            .I(N__31330));
    LocalMux I__5039 (
            .O(N__31336),
            .I(n2117));
    Odrv4 I__5038 (
            .O(N__31333),
            .I(n2117));
    Odrv4 I__5037 (
            .O(N__31330),
            .I(n2117));
    InMux I__5036 (
            .O(N__31323),
            .I(N__31320));
    LocalMux I__5035 (
            .O(N__31320),
            .I(N__31317));
    Odrv4 I__5034 (
            .O(N__31317),
            .I(n2089));
    InMux I__5033 (
            .O(N__31314),
            .I(N__31309));
    InMux I__5032 (
            .O(N__31313),
            .I(N__31306));
    CascadeMux I__5031 (
            .O(N__31312),
            .I(N__31303));
    LocalMux I__5030 (
            .O(N__31309),
            .I(N__31300));
    LocalMux I__5029 (
            .O(N__31306),
            .I(N__31297));
    InMux I__5028 (
            .O(N__31303),
            .I(N__31294));
    Span4Mux_h I__5027 (
            .O(N__31300),
            .I(N__31291));
    Span4Mux_h I__5026 (
            .O(N__31297),
            .I(N__31288));
    LocalMux I__5025 (
            .O(N__31294),
            .I(N__31285));
    Odrv4 I__5024 (
            .O(N__31291),
            .I(n2121));
    Odrv4 I__5023 (
            .O(N__31288),
            .I(n2121));
    Odrv4 I__5022 (
            .O(N__31285),
            .I(n2121));
    InMux I__5021 (
            .O(N__31278),
            .I(N__31275));
    LocalMux I__5020 (
            .O(N__31275),
            .I(N__31272));
    Span4Mux_v I__5019 (
            .O(N__31272),
            .I(N__31269));
    Odrv4 I__5018 (
            .O(N__31269),
            .I(n2501));
    InMux I__5017 (
            .O(N__31266),
            .I(bfn_6_21_0_));
    InMux I__5016 (
            .O(N__31263),
            .I(n12717));
    InMux I__5015 (
            .O(N__31260),
            .I(n12651));
    InMux I__5014 (
            .O(N__31257),
            .I(n12652));
    InMux I__5013 (
            .O(N__31254),
            .I(N__31251));
    LocalMux I__5012 (
            .O(N__31251),
            .I(N__31248));
    Odrv4 I__5011 (
            .O(N__31248),
            .I(n2086));
    InMux I__5010 (
            .O(N__31245),
            .I(n12653));
    InMux I__5009 (
            .O(N__31242),
            .I(bfn_6_19_0_));
    CascadeMux I__5008 (
            .O(N__31239),
            .I(N__31236));
    InMux I__5007 (
            .O(N__31236),
            .I(N__31233));
    LocalMux I__5006 (
            .O(N__31233),
            .I(n2084));
    InMux I__5005 (
            .O(N__31230),
            .I(n12655));
    InMux I__5004 (
            .O(N__31227),
            .I(n12656));
    CascadeMux I__5003 (
            .O(N__31224),
            .I(N__31221));
    InMux I__5002 (
            .O(N__31221),
            .I(N__31218));
    LocalMux I__5001 (
            .O(N__31218),
            .I(N__31214));
    InMux I__5000 (
            .O(N__31217),
            .I(N__31211));
    Odrv4 I__4999 (
            .O(N__31214),
            .I(n2115));
    LocalMux I__4998 (
            .O(N__31211),
            .I(n2115));
    InMux I__4997 (
            .O(N__31206),
            .I(N__31203));
    LocalMux I__4996 (
            .O(N__31203),
            .I(n2091));
    CascadeMux I__4995 (
            .O(N__31200),
            .I(N__31196));
    CascadeMux I__4994 (
            .O(N__31199),
            .I(N__31193));
    InMux I__4993 (
            .O(N__31196),
            .I(N__31190));
    InMux I__4992 (
            .O(N__31193),
            .I(N__31187));
    LocalMux I__4991 (
            .O(N__31190),
            .I(N__31182));
    LocalMux I__4990 (
            .O(N__31187),
            .I(N__31182));
    Span4Mux_h I__4989 (
            .O(N__31182),
            .I(N__31178));
    InMux I__4988 (
            .O(N__31181),
            .I(N__31175));
    Odrv4 I__4987 (
            .O(N__31178),
            .I(n2123));
    LocalMux I__4986 (
            .O(N__31175),
            .I(n2123));
    CascadeMux I__4985 (
            .O(N__31170),
            .I(N__31167));
    InMux I__4984 (
            .O(N__31167),
            .I(N__31164));
    LocalMux I__4983 (
            .O(N__31164),
            .I(N__31161));
    Span4Mux_h I__4982 (
            .O(N__31161),
            .I(N__31158));
    Odrv4 I__4981 (
            .O(N__31158),
            .I(n2097));
    InMux I__4980 (
            .O(N__31155),
            .I(n12642));
    InMux I__4979 (
            .O(N__31152),
            .I(N__31149));
    LocalMux I__4978 (
            .O(N__31149),
            .I(n2096));
    InMux I__4977 (
            .O(N__31146),
            .I(n12643));
    InMux I__4976 (
            .O(N__31143),
            .I(N__31140));
    LocalMux I__4975 (
            .O(N__31140),
            .I(n2095));
    InMux I__4974 (
            .O(N__31137),
            .I(n12644));
    CascadeMux I__4973 (
            .O(N__31134),
            .I(N__31131));
    InMux I__4972 (
            .O(N__31131),
            .I(N__31128));
    LocalMux I__4971 (
            .O(N__31128),
            .I(n2094));
    InMux I__4970 (
            .O(N__31125),
            .I(n12645));
    InMux I__4969 (
            .O(N__31122),
            .I(N__31119));
    LocalMux I__4968 (
            .O(N__31119),
            .I(n2093));
    InMux I__4967 (
            .O(N__31116),
            .I(bfn_6_18_0_));
    InMux I__4966 (
            .O(N__31113),
            .I(N__31110));
    LocalMux I__4965 (
            .O(N__31110),
            .I(n2092));
    InMux I__4964 (
            .O(N__31107),
            .I(n12647));
    InMux I__4963 (
            .O(N__31104),
            .I(n12648));
    InMux I__4962 (
            .O(N__31101),
            .I(N__31098));
    LocalMux I__4961 (
            .O(N__31098),
            .I(n2090));
    InMux I__4960 (
            .O(N__31095),
            .I(n12649));
    InMux I__4959 (
            .O(N__31092),
            .I(n12650));
    InMux I__4958 (
            .O(N__31089),
            .I(N__31086));
    LocalMux I__4957 (
            .O(N__31086),
            .I(n14272));
    InMux I__4956 (
            .O(N__31083),
            .I(N__31080));
    LocalMux I__4955 (
            .O(N__31080),
            .I(n14268));
    CascadeMux I__4954 (
            .O(N__31077),
            .I(n14262_cascade_));
    InMux I__4953 (
            .O(N__31074),
            .I(N__31071));
    LocalMux I__4952 (
            .O(N__31071),
            .I(n14282));
    InMux I__4951 (
            .O(N__31068),
            .I(N__31065));
    LocalMux I__4950 (
            .O(N__31065),
            .I(N__31060));
    InMux I__4949 (
            .O(N__31064),
            .I(N__31057));
    InMux I__4948 (
            .O(N__31063),
            .I(N__31054));
    Odrv4 I__4947 (
            .O(N__31060),
            .I(n3111));
    LocalMux I__4946 (
            .O(N__31057),
            .I(n3111));
    LocalMux I__4945 (
            .O(N__31054),
            .I(n3111));
    CascadeMux I__4944 (
            .O(N__31047),
            .I(N__31044));
    InMux I__4943 (
            .O(N__31044),
            .I(N__31041));
    LocalMux I__4942 (
            .O(N__31041),
            .I(N__31038));
    Span4Mux_s1_v I__4941 (
            .O(N__31038),
            .I(N__31035));
    Odrv4 I__4940 (
            .O(N__31035),
            .I(n3178));
    InMux I__4939 (
            .O(N__31032),
            .I(N__31029));
    LocalMux I__4938 (
            .O(N__31029),
            .I(N__31024));
    InMux I__4937 (
            .O(N__31028),
            .I(N__31021));
    InMux I__4936 (
            .O(N__31027),
            .I(N__31018));
    Odrv4 I__4935 (
            .O(N__31024),
            .I(n3110));
    LocalMux I__4934 (
            .O(N__31021),
            .I(n3110));
    LocalMux I__4933 (
            .O(N__31018),
            .I(n3110));
    InMux I__4932 (
            .O(N__31011),
            .I(N__31008));
    LocalMux I__4931 (
            .O(N__31008),
            .I(N__31005));
    Odrv4 I__4930 (
            .O(N__31005),
            .I(n3177));
    InMux I__4929 (
            .O(N__31002),
            .I(N__30999));
    LocalMux I__4928 (
            .O(N__30999),
            .I(N__30996));
    Odrv4 I__4927 (
            .O(N__30996),
            .I(n2283));
    CascadeMux I__4926 (
            .O(N__30993),
            .I(N__30989));
    InMux I__4925 (
            .O(N__30992),
            .I(N__30986));
    InMux I__4924 (
            .O(N__30989),
            .I(N__30982));
    LocalMux I__4923 (
            .O(N__30986),
            .I(N__30979));
    InMux I__4922 (
            .O(N__30985),
            .I(N__30976));
    LocalMux I__4921 (
            .O(N__30982),
            .I(N__30973));
    Span4Mux_v I__4920 (
            .O(N__30979),
            .I(N__30968));
    LocalMux I__4919 (
            .O(N__30976),
            .I(N__30968));
    Odrv4 I__4918 (
            .O(N__30973),
            .I(n2216));
    Odrv4 I__4917 (
            .O(N__30968),
            .I(n2216));
    InMux I__4916 (
            .O(N__30963),
            .I(N__30959));
    InMux I__4915 (
            .O(N__30962),
            .I(N__30956));
    LocalMux I__4914 (
            .O(N__30959),
            .I(N__30953));
    LocalMux I__4913 (
            .O(N__30956),
            .I(N__30949));
    Span4Mux_v I__4912 (
            .O(N__30953),
            .I(N__30946));
    InMux I__4911 (
            .O(N__30952),
            .I(N__30943));
    Span4Mux_v I__4910 (
            .O(N__30949),
            .I(N__30936));
    Span4Mux_h I__4909 (
            .O(N__30946),
            .I(N__30936));
    LocalMux I__4908 (
            .O(N__30943),
            .I(N__30936));
    Span4Mux_v I__4907 (
            .O(N__30936),
            .I(N__30933));
    Odrv4 I__4906 (
            .O(N__30933),
            .I(n2315));
    InMux I__4905 (
            .O(N__30930),
            .I(bfn_6_17_0_));
    InMux I__4904 (
            .O(N__30927),
            .I(n12639));
    CascadeMux I__4903 (
            .O(N__30924),
            .I(N__30921));
    InMux I__4902 (
            .O(N__30921),
            .I(N__30918));
    LocalMux I__4901 (
            .O(N__30918),
            .I(n2099));
    InMux I__4900 (
            .O(N__30915),
            .I(n12640));
    InMux I__4899 (
            .O(N__30912),
            .I(N__30909));
    LocalMux I__4898 (
            .O(N__30909),
            .I(n2098));
    InMux I__4897 (
            .O(N__30906),
            .I(n12641));
    InMux I__4896 (
            .O(N__30903),
            .I(N__30900));
    LocalMux I__4895 (
            .O(N__30900),
            .I(N__30897));
    Odrv12 I__4894 (
            .O(N__30897),
            .I(n3185));
    InMux I__4893 (
            .O(N__30894),
            .I(N__30891));
    LocalMux I__4892 (
            .O(N__30891),
            .I(N__30887));
    InMux I__4891 (
            .O(N__30890),
            .I(N__30884));
    Span4Mux_h I__4890 (
            .O(N__30887),
            .I(N__30878));
    LocalMux I__4889 (
            .O(N__30884),
            .I(N__30878));
    InMux I__4888 (
            .O(N__30883),
            .I(N__30875));
    Odrv4 I__4887 (
            .O(N__30878),
            .I(n3118));
    LocalMux I__4886 (
            .O(N__30875),
            .I(n3118));
    CascadeMux I__4885 (
            .O(N__30870),
            .I(n27_adj_716_cascade_));
    InMux I__4884 (
            .O(N__30867),
            .I(N__30864));
    LocalMux I__4883 (
            .O(N__30864),
            .I(n14266));
    InMux I__4882 (
            .O(N__30861),
            .I(N__30858));
    LocalMux I__4881 (
            .O(N__30858),
            .I(n35_adj_719));
    CascadeMux I__4880 (
            .O(N__30855),
            .I(n17_adj_714_cascade_));
    InMux I__4879 (
            .O(N__30852),
            .I(N__30848));
    InMux I__4878 (
            .O(N__30851),
            .I(N__30844));
    LocalMux I__4877 (
            .O(N__30848),
            .I(N__30841));
    InMux I__4876 (
            .O(N__30847),
            .I(N__30838));
    LocalMux I__4875 (
            .O(N__30844),
            .I(n3109));
    Odrv4 I__4874 (
            .O(N__30841),
            .I(n3109));
    LocalMux I__4873 (
            .O(N__30838),
            .I(n3109));
    CascadeMux I__4872 (
            .O(N__30831),
            .I(N__30828));
    InMux I__4871 (
            .O(N__30828),
            .I(N__30825));
    LocalMux I__4870 (
            .O(N__30825),
            .I(N__30822));
    Odrv4 I__4869 (
            .O(N__30822),
            .I(n3176));
    CascadeMux I__4868 (
            .O(N__30819),
            .I(n33_adj_718_cascade_));
    InMux I__4867 (
            .O(N__30816),
            .I(N__30813));
    LocalMux I__4866 (
            .O(N__30813),
            .I(N__30808));
    CascadeMux I__4865 (
            .O(N__30812),
            .I(N__30805));
    CascadeMux I__4864 (
            .O(N__30811),
            .I(N__30802));
    Span4Mux_h I__4863 (
            .O(N__30808),
            .I(N__30799));
    InMux I__4862 (
            .O(N__30805),
            .I(N__30796));
    InMux I__4861 (
            .O(N__30802),
            .I(N__30793));
    Odrv4 I__4860 (
            .O(N__30799),
            .I(n3124));
    LocalMux I__4859 (
            .O(N__30796),
            .I(n3124));
    LocalMux I__4858 (
            .O(N__30793),
            .I(n3124));
    CascadeMux I__4857 (
            .O(N__30786),
            .I(N__30783));
    InMux I__4856 (
            .O(N__30783),
            .I(N__30780));
    LocalMux I__4855 (
            .O(N__30780),
            .I(N__30777));
    Odrv4 I__4854 (
            .O(N__30777),
            .I(n3191));
    InMux I__4853 (
            .O(N__30774),
            .I(N__30771));
    LocalMux I__4852 (
            .O(N__30771),
            .I(n14804));
    CascadeMux I__4851 (
            .O(N__30768),
            .I(N__30765));
    InMux I__4850 (
            .O(N__30765),
            .I(N__30762));
    LocalMux I__4849 (
            .O(N__30762),
            .I(n14025));
    CascadeMux I__4848 (
            .O(N__30759),
            .I(n3237_cascade_));
    InMux I__4847 (
            .O(N__30756),
            .I(N__30753));
    LocalMux I__4846 (
            .O(N__30753),
            .I(n13_adj_713));
    InMux I__4845 (
            .O(N__30750),
            .I(N__30747));
    LocalMux I__4844 (
            .O(N__30747),
            .I(N__30744));
    Span4Mux_h I__4843 (
            .O(N__30744),
            .I(N__30741));
    Odrv4 I__4842 (
            .O(N__30741),
            .I(n3179));
    InMux I__4841 (
            .O(N__30738),
            .I(N__30734));
    InMux I__4840 (
            .O(N__30737),
            .I(N__30731));
    LocalMux I__4839 (
            .O(N__30734),
            .I(N__30727));
    LocalMux I__4838 (
            .O(N__30731),
            .I(N__30724));
    InMux I__4837 (
            .O(N__30730),
            .I(N__30721));
    Span4Mux_s3_h I__4836 (
            .O(N__30727),
            .I(N__30716));
    Span4Mux_s1_v I__4835 (
            .O(N__30724),
            .I(N__30716));
    LocalMux I__4834 (
            .O(N__30721),
            .I(n3112));
    Odrv4 I__4833 (
            .O(N__30716),
            .I(n3112));
    InMux I__4832 (
            .O(N__30711),
            .I(N__30708));
    LocalMux I__4831 (
            .O(N__30708),
            .I(n14770));
    CascadeMux I__4830 (
            .O(N__30705),
            .I(n14776_cascade_));
    InMux I__4829 (
            .O(N__30702),
            .I(N__30699));
    LocalMux I__4828 (
            .O(N__30699),
            .I(N__30696));
    Span4Mux_s3_v I__4827 (
            .O(N__30696),
            .I(N__30693));
    Span4Mux_h I__4826 (
            .O(N__30693),
            .I(N__30689));
    InMux I__4825 (
            .O(N__30692),
            .I(N__30686));
    Odrv4 I__4824 (
            .O(N__30689),
            .I(n3122));
    LocalMux I__4823 (
            .O(N__30686),
            .I(n3122));
    CascadeMux I__4822 (
            .O(N__30681),
            .I(N__30678));
    InMux I__4821 (
            .O(N__30678),
            .I(N__30675));
    LocalMux I__4820 (
            .O(N__30675),
            .I(N__30672));
    Odrv4 I__4819 (
            .O(N__30672),
            .I(n3189));
    InMux I__4818 (
            .O(N__30669),
            .I(N__30666));
    LocalMux I__4817 (
            .O(N__30666),
            .I(N__30662));
    InMux I__4816 (
            .O(N__30665),
            .I(N__30659));
    Span4Mux_h I__4815 (
            .O(N__30662),
            .I(N__30653));
    LocalMux I__4814 (
            .O(N__30659),
            .I(N__30653));
    InMux I__4813 (
            .O(N__30658),
            .I(N__30650));
    Odrv4 I__4812 (
            .O(N__30653),
            .I(n3116));
    LocalMux I__4811 (
            .O(N__30650),
            .I(n3116));
    CascadeMux I__4810 (
            .O(N__30645),
            .I(N__30642));
    InMux I__4809 (
            .O(N__30642),
            .I(N__30639));
    LocalMux I__4808 (
            .O(N__30639),
            .I(N__30636));
    Odrv4 I__4807 (
            .O(N__30636),
            .I(n3183));
    CascadeMux I__4806 (
            .O(N__30633),
            .I(n3030_cascade_));
    InMux I__4805 (
            .O(N__30630),
            .I(N__30627));
    LocalMux I__4804 (
            .O(N__30627),
            .I(n11947));
    CascadeMux I__4803 (
            .O(N__30624),
            .I(N__30620));
    InMux I__4802 (
            .O(N__30623),
            .I(N__30617));
    InMux I__4801 (
            .O(N__30620),
            .I(N__30614));
    LocalMux I__4800 (
            .O(N__30617),
            .I(N__30609));
    LocalMux I__4799 (
            .O(N__30614),
            .I(N__30609));
    Span4Mux_h I__4798 (
            .O(N__30609),
            .I(N__30605));
    InMux I__4797 (
            .O(N__30608),
            .I(N__30602));
    Odrv4 I__4796 (
            .O(N__30605),
            .I(n3019));
    LocalMux I__4795 (
            .O(N__30602),
            .I(n3019));
    CascadeMux I__4794 (
            .O(N__30597),
            .I(N__30594));
    InMux I__4793 (
            .O(N__30594),
            .I(N__30591));
    LocalMux I__4792 (
            .O(N__30591),
            .I(N__30588));
    Span4Mux_v I__4791 (
            .O(N__30588),
            .I(N__30584));
    CascadeMux I__4790 (
            .O(N__30587),
            .I(N__30581));
    Span4Mux_s0_h I__4789 (
            .O(N__30584),
            .I(N__30577));
    InMux I__4788 (
            .O(N__30581),
            .I(N__30574));
    InMux I__4787 (
            .O(N__30580),
            .I(N__30571));
    Odrv4 I__4786 (
            .O(N__30577),
            .I(n3027));
    LocalMux I__4785 (
            .O(N__30574),
            .I(n3027));
    LocalMux I__4784 (
            .O(N__30571),
            .I(n3027));
    CascadeMux I__4783 (
            .O(N__30564),
            .I(n13871_cascade_));
    CascadeMux I__4782 (
            .O(N__30561),
            .I(N__30557));
    InMux I__4781 (
            .O(N__30560),
            .I(N__30554));
    InMux I__4780 (
            .O(N__30557),
            .I(N__30551));
    LocalMux I__4779 (
            .O(N__30554),
            .I(N__30548));
    LocalMux I__4778 (
            .O(N__30551),
            .I(N__30545));
    Span4Mux_v I__4777 (
            .O(N__30548),
            .I(N__30541));
    Span4Mux_v I__4776 (
            .O(N__30545),
            .I(N__30538));
    InMux I__4775 (
            .O(N__30544),
            .I(N__30535));
    Odrv4 I__4774 (
            .O(N__30541),
            .I(n3023));
    Odrv4 I__4773 (
            .O(N__30538),
            .I(n3023));
    LocalMux I__4772 (
            .O(N__30535),
            .I(n3023));
    CascadeMux I__4771 (
            .O(N__30528),
            .I(N__30525));
    InMux I__4770 (
            .O(N__30525),
            .I(N__30522));
    LocalMux I__4769 (
            .O(N__30522),
            .I(n14078));
    InMux I__4768 (
            .O(N__30519),
            .I(N__30516));
    LocalMux I__4767 (
            .O(N__30516),
            .I(N__30513));
    Odrv4 I__4766 (
            .O(N__30513),
            .I(n3199));
    CascadeMux I__4765 (
            .O(N__30510),
            .I(N__30507));
    InMux I__4764 (
            .O(N__30507),
            .I(N__30503));
    InMux I__4763 (
            .O(N__30506),
            .I(N__30500));
    LocalMux I__4762 (
            .O(N__30503),
            .I(N__30497));
    LocalMux I__4761 (
            .O(N__30500),
            .I(n3132));
    Odrv4 I__4760 (
            .O(N__30497),
            .I(n3132));
    CascadeMux I__4759 (
            .O(N__30492),
            .I(N__30489));
    InMux I__4758 (
            .O(N__30489),
            .I(N__30485));
    InMux I__4757 (
            .O(N__30488),
            .I(N__30481));
    LocalMux I__4756 (
            .O(N__30485),
            .I(N__30478));
    InMux I__4755 (
            .O(N__30484),
            .I(N__30475));
    LocalMux I__4754 (
            .O(N__30481),
            .I(n3129));
    Odrv4 I__4753 (
            .O(N__30478),
            .I(n3129));
    LocalMux I__4752 (
            .O(N__30475),
            .I(n3129));
    CascadeMux I__4751 (
            .O(N__30468),
            .I(N__30465));
    InMux I__4750 (
            .O(N__30465),
            .I(N__30462));
    LocalMux I__4749 (
            .O(N__30462),
            .I(N__30459));
    Span4Mux_h I__4748 (
            .O(N__30459),
            .I(N__30456));
    Odrv4 I__4747 (
            .O(N__30456),
            .I(n3196));
    CascadeMux I__4746 (
            .O(N__30453),
            .I(n3228_cascade_));
    InMux I__4745 (
            .O(N__30450),
            .I(N__30447));
    LocalMux I__4744 (
            .O(N__30447),
            .I(n14768));
    InMux I__4743 (
            .O(N__30444),
            .I(N__30441));
    LocalMux I__4742 (
            .O(N__30441),
            .I(N__30438));
    Span4Mux_h I__4741 (
            .O(N__30438),
            .I(N__30435));
    Odrv4 I__4740 (
            .O(N__30435),
            .I(n3200));
    CascadeMux I__4739 (
            .O(N__30432),
            .I(N__30428));
    CascadeMux I__4738 (
            .O(N__30431),
            .I(N__30425));
    InMux I__4737 (
            .O(N__30428),
            .I(N__30422));
    InMux I__4736 (
            .O(N__30425),
            .I(N__30418));
    LocalMux I__4735 (
            .O(N__30422),
            .I(N__30415));
    InMux I__4734 (
            .O(N__30421),
            .I(N__30412));
    LocalMux I__4733 (
            .O(N__30418),
            .I(n3133));
    Odrv4 I__4732 (
            .O(N__30415),
            .I(n3133));
    LocalMux I__4731 (
            .O(N__30412),
            .I(n3133));
    InMux I__4730 (
            .O(N__30405),
            .I(N__30402));
    LocalMux I__4729 (
            .O(N__30402),
            .I(N__30399));
    Odrv4 I__4728 (
            .O(N__30399),
            .I(n3198));
    CascadeMux I__4727 (
            .O(N__30396),
            .I(N__30393));
    InMux I__4726 (
            .O(N__30393),
            .I(N__30390));
    LocalMux I__4725 (
            .O(N__30390),
            .I(N__30386));
    InMux I__4724 (
            .O(N__30389),
            .I(N__30382));
    Span4Mux_v I__4723 (
            .O(N__30386),
            .I(N__30379));
    InMux I__4722 (
            .O(N__30385),
            .I(N__30376));
    LocalMux I__4721 (
            .O(N__30382),
            .I(n3131));
    Odrv4 I__4720 (
            .O(N__30379),
            .I(n3131));
    LocalMux I__4719 (
            .O(N__30376),
            .I(n3131));
    InMux I__4718 (
            .O(N__30369),
            .I(N__30365));
    InMux I__4717 (
            .O(N__30368),
            .I(N__30362));
    LocalMux I__4716 (
            .O(N__30365),
            .I(N__30359));
    LocalMux I__4715 (
            .O(N__30362),
            .I(N__30356));
    Span4Mux_v I__4714 (
            .O(N__30359),
            .I(N__30352));
    Span4Mux_s3_h I__4713 (
            .O(N__30356),
            .I(N__30349));
    InMux I__4712 (
            .O(N__30355),
            .I(N__30346));
    Odrv4 I__4711 (
            .O(N__30352),
            .I(n2917));
    Odrv4 I__4710 (
            .O(N__30349),
            .I(n2917));
    LocalMux I__4709 (
            .O(N__30346),
            .I(n2917));
    CascadeMux I__4708 (
            .O(N__30339),
            .I(N__30336));
    InMux I__4707 (
            .O(N__30336),
            .I(N__30333));
    LocalMux I__4706 (
            .O(N__30333),
            .I(N__30330));
    Span4Mux_v I__4705 (
            .O(N__30330),
            .I(N__30327));
    Odrv4 I__4704 (
            .O(N__30327),
            .I(n2984));
    InMux I__4703 (
            .O(N__30324),
            .I(N__30320));
    InMux I__4702 (
            .O(N__30323),
            .I(N__30317));
    LocalMux I__4701 (
            .O(N__30320),
            .I(N__30314));
    LocalMux I__4700 (
            .O(N__30317),
            .I(N__30311));
    Span4Mux_s1_v I__4699 (
            .O(N__30314),
            .I(N__30307));
    Span4Mux_s3_v I__4698 (
            .O(N__30311),
            .I(N__30304));
    InMux I__4697 (
            .O(N__30310),
            .I(N__30301));
    Odrv4 I__4696 (
            .O(N__30307),
            .I(n3016));
    Odrv4 I__4695 (
            .O(N__30304),
            .I(n3016));
    LocalMux I__4694 (
            .O(N__30301),
            .I(n3016));
    InMux I__4693 (
            .O(N__30294),
            .I(N__30291));
    LocalMux I__4692 (
            .O(N__30291),
            .I(N__30287));
    InMux I__4691 (
            .O(N__30290),
            .I(N__30283));
    Span4Mux_h I__4690 (
            .O(N__30287),
            .I(N__30280));
    InMux I__4689 (
            .O(N__30286),
            .I(N__30277));
    LocalMux I__4688 (
            .O(N__30283),
            .I(n2913));
    Odrv4 I__4687 (
            .O(N__30280),
            .I(n2913));
    LocalMux I__4686 (
            .O(N__30277),
            .I(n2913));
    CascadeMux I__4685 (
            .O(N__30270),
            .I(N__30267));
    InMux I__4684 (
            .O(N__30267),
            .I(N__30264));
    LocalMux I__4683 (
            .O(N__30264),
            .I(N__30261));
    Odrv4 I__4682 (
            .O(N__30261),
            .I(n2980));
    CascadeMux I__4681 (
            .O(N__30258),
            .I(N__30255));
    InMux I__4680 (
            .O(N__30255),
            .I(N__30252));
    LocalMux I__4679 (
            .O(N__30252),
            .I(N__30248));
    InMux I__4678 (
            .O(N__30251),
            .I(N__30245));
    Span4Mux_s1_v I__4677 (
            .O(N__30248),
            .I(N__30242));
    LocalMux I__4676 (
            .O(N__30245),
            .I(N__30239));
    Span4Mux_v I__4675 (
            .O(N__30242),
            .I(N__30235));
    Span4Mux_h I__4674 (
            .O(N__30239),
            .I(N__30232));
    InMux I__4673 (
            .O(N__30238),
            .I(N__30229));
    Odrv4 I__4672 (
            .O(N__30235),
            .I(n3012));
    Odrv4 I__4671 (
            .O(N__30232),
            .I(n3012));
    LocalMux I__4670 (
            .O(N__30229),
            .I(n3012));
    InMux I__4669 (
            .O(N__30222),
            .I(N__30217));
    InMux I__4668 (
            .O(N__30221),
            .I(N__30214));
    InMux I__4667 (
            .O(N__30220),
            .I(N__30211));
    LocalMux I__4666 (
            .O(N__30217),
            .I(N__30208));
    LocalMux I__4665 (
            .O(N__30214),
            .I(N__30203));
    LocalMux I__4664 (
            .O(N__30211),
            .I(N__30203));
    Odrv4 I__4663 (
            .O(N__30208),
            .I(n2933));
    Odrv4 I__4662 (
            .O(N__30203),
            .I(n2933));
    InMux I__4661 (
            .O(N__30198),
            .I(N__30195));
    LocalMux I__4660 (
            .O(N__30195),
            .I(n12053));
    InMux I__4659 (
            .O(N__30192),
            .I(N__30189));
    LocalMux I__4658 (
            .O(N__30189),
            .I(N__30186));
    Span4Mux_h I__4657 (
            .O(N__30186),
            .I(N__30183));
    Odrv4 I__4656 (
            .O(N__30183),
            .I(n2987));
    CascadeMux I__4655 (
            .O(N__30180),
            .I(N__30176));
    InMux I__4654 (
            .O(N__30179),
            .I(N__30173));
    InMux I__4653 (
            .O(N__30176),
            .I(N__30169));
    LocalMux I__4652 (
            .O(N__30173),
            .I(N__30166));
    InMux I__4651 (
            .O(N__30172),
            .I(N__30163));
    LocalMux I__4650 (
            .O(N__30169),
            .I(n2920));
    Odrv4 I__4649 (
            .O(N__30166),
            .I(n2920));
    LocalMux I__4648 (
            .O(N__30163),
            .I(n2920));
    InMux I__4647 (
            .O(N__30156),
            .I(N__30153));
    LocalMux I__4646 (
            .O(N__30153),
            .I(N__30150));
    Span4Mux_h I__4645 (
            .O(N__30150),
            .I(N__30147));
    Odrv4 I__4644 (
            .O(N__30147),
            .I(n2999));
    CascadeMux I__4643 (
            .O(N__30144),
            .I(N__30141));
    InMux I__4642 (
            .O(N__30141),
            .I(N__30137));
    InMux I__4641 (
            .O(N__30140),
            .I(N__30134));
    LocalMux I__4640 (
            .O(N__30137),
            .I(N__30131));
    LocalMux I__4639 (
            .O(N__30134),
            .I(N__30127));
    Span4Mux_h I__4638 (
            .O(N__30131),
            .I(N__30124));
    InMux I__4637 (
            .O(N__30130),
            .I(N__30121));
    Span4Mux_h I__4636 (
            .O(N__30127),
            .I(N__30118));
    Odrv4 I__4635 (
            .O(N__30124),
            .I(n2932));
    LocalMux I__4634 (
            .O(N__30121),
            .I(n2932));
    Odrv4 I__4633 (
            .O(N__30118),
            .I(n2932));
    InMux I__4632 (
            .O(N__30111),
            .I(N__30108));
    LocalMux I__4631 (
            .O(N__30108),
            .I(N__30105));
    Span4Mux_v I__4630 (
            .O(N__30105),
            .I(N__30102));
    Odrv4 I__4629 (
            .O(N__30102),
            .I(n3001));
    CascadeMux I__4628 (
            .O(N__30099),
            .I(N__30096));
    InMux I__4627 (
            .O(N__30096),
            .I(N__30092));
    InMux I__4626 (
            .O(N__30095),
            .I(N__30089));
    LocalMux I__4625 (
            .O(N__30092),
            .I(N__30086));
    LocalMux I__4624 (
            .O(N__30089),
            .I(n3033));
    Odrv4 I__4623 (
            .O(N__30086),
            .I(n3033));
    CascadeMux I__4622 (
            .O(N__30081),
            .I(n3033_cascade_));
    CascadeMux I__4621 (
            .O(N__30078),
            .I(N__30074));
    InMux I__4620 (
            .O(N__30077),
            .I(N__30070));
    InMux I__4619 (
            .O(N__30074),
            .I(N__30067));
    InMux I__4618 (
            .O(N__30073),
            .I(N__30064));
    LocalMux I__4617 (
            .O(N__30070),
            .I(n3032));
    LocalMux I__4616 (
            .O(N__30067),
            .I(n3032));
    LocalMux I__4615 (
            .O(N__30064),
            .I(n3032));
    InMux I__4614 (
            .O(N__30057),
            .I(N__30054));
    LocalMux I__4613 (
            .O(N__30054),
            .I(N__30051));
    Span4Mux_h I__4612 (
            .O(N__30051),
            .I(N__30048));
    Odrv4 I__4611 (
            .O(N__30048),
            .I(n3182));
    CascadeMux I__4610 (
            .O(N__30045),
            .I(N__30042));
    InMux I__4609 (
            .O(N__30042),
            .I(N__30039));
    LocalMux I__4608 (
            .O(N__30039),
            .I(N__30035));
    InMux I__4607 (
            .O(N__30038),
            .I(N__30032));
    Span4Mux_h I__4606 (
            .O(N__30035),
            .I(N__30027));
    LocalMux I__4605 (
            .O(N__30032),
            .I(N__30027));
    Span4Mux_v I__4604 (
            .O(N__30027),
            .I(N__30024));
    Odrv4 I__4603 (
            .O(N__30024),
            .I(n3115));
    InMux I__4602 (
            .O(N__30021),
            .I(N__30018));
    LocalMux I__4601 (
            .O(N__30018),
            .I(N__30015));
    Span4Mux_h I__4600 (
            .O(N__30015),
            .I(N__30012));
    Odrv4 I__4599 (
            .O(N__30012),
            .I(n2998));
    CascadeMux I__4598 (
            .O(N__30009),
            .I(N__30004));
    CascadeMux I__4597 (
            .O(N__30008),
            .I(N__30001));
    InMux I__4596 (
            .O(N__30007),
            .I(N__29998));
    InMux I__4595 (
            .O(N__30004),
            .I(N__29995));
    InMux I__4594 (
            .O(N__30001),
            .I(N__29992));
    LocalMux I__4593 (
            .O(N__29998),
            .I(N__29989));
    LocalMux I__4592 (
            .O(N__29995),
            .I(N__29984));
    LocalMux I__4591 (
            .O(N__29992),
            .I(N__29984));
    Odrv4 I__4590 (
            .O(N__29989),
            .I(n2931));
    Odrv4 I__4589 (
            .O(N__29984),
            .I(n2931));
    CascadeMux I__4588 (
            .O(N__29979),
            .I(N__29975));
    CascadeMux I__4587 (
            .O(N__29978),
            .I(N__29972));
    InMux I__4586 (
            .O(N__29975),
            .I(N__29969));
    InMux I__4585 (
            .O(N__29972),
            .I(N__29966));
    LocalMux I__4584 (
            .O(N__29969),
            .I(N__29963));
    LocalMux I__4583 (
            .O(N__29966),
            .I(n3030));
    Odrv4 I__4582 (
            .O(N__29963),
            .I(n3030));
    InMux I__4581 (
            .O(N__29958),
            .I(N__29955));
    LocalMux I__4580 (
            .O(N__29955),
            .I(N__29951));
    CascadeMux I__4579 (
            .O(N__29954),
            .I(N__29948));
    Span4Mux_v I__4578 (
            .O(N__29951),
            .I(N__29944));
    InMux I__4577 (
            .O(N__29948),
            .I(N__29941));
    InMux I__4576 (
            .O(N__29947),
            .I(N__29938));
    Odrv4 I__4575 (
            .O(N__29944),
            .I(n3029));
    LocalMux I__4574 (
            .O(N__29941),
            .I(n3029));
    LocalMux I__4573 (
            .O(N__29938),
            .I(n3029));
    CascadeMux I__4572 (
            .O(N__29931),
            .I(N__29928));
    InMux I__4571 (
            .O(N__29928),
            .I(N__29923));
    InMux I__4570 (
            .O(N__29927),
            .I(N__29920));
    InMux I__4569 (
            .O(N__29926),
            .I(N__29917));
    LocalMux I__4568 (
            .O(N__29923),
            .I(N__29914));
    LocalMux I__4567 (
            .O(N__29920),
            .I(n3031));
    LocalMux I__4566 (
            .O(N__29917),
            .I(n3031));
    Odrv4 I__4565 (
            .O(N__29914),
            .I(n3031));
    InMux I__4564 (
            .O(N__29907),
            .I(N__29904));
    LocalMux I__4563 (
            .O(N__29904),
            .I(N__29901));
    Span4Mux_v I__4562 (
            .O(N__29901),
            .I(N__29898));
    Odrv4 I__4561 (
            .O(N__29898),
            .I(n2896));
    CascadeMux I__4560 (
            .O(N__29895),
            .I(N__29892));
    InMux I__4559 (
            .O(N__29892),
            .I(N__29889));
    LocalMux I__4558 (
            .O(N__29889),
            .I(N__29885));
    InMux I__4557 (
            .O(N__29888),
            .I(N__29881));
    Span4Mux_v I__4556 (
            .O(N__29885),
            .I(N__29878));
    CascadeMux I__4555 (
            .O(N__29884),
            .I(N__29875));
    LocalMux I__4554 (
            .O(N__29881),
            .I(N__29872));
    Span4Mux_h I__4553 (
            .O(N__29878),
            .I(N__29869));
    InMux I__4552 (
            .O(N__29875),
            .I(N__29866));
    Span4Mux_v I__4551 (
            .O(N__29872),
            .I(N__29863));
    Odrv4 I__4550 (
            .O(N__29869),
            .I(n2829));
    LocalMux I__4549 (
            .O(N__29866),
            .I(n2829));
    Odrv4 I__4548 (
            .O(N__29863),
            .I(n2829));
    InMux I__4547 (
            .O(N__29856),
            .I(N__29853));
    LocalMux I__4546 (
            .O(N__29853),
            .I(N__29849));
    InMux I__4545 (
            .O(N__29852),
            .I(N__29845));
    Span4Mux_h I__4544 (
            .O(N__29849),
            .I(N__29842));
    InMux I__4543 (
            .O(N__29848),
            .I(N__29839));
    LocalMux I__4542 (
            .O(N__29845),
            .I(n2928));
    Odrv4 I__4541 (
            .O(N__29842),
            .I(n2928));
    LocalMux I__4540 (
            .O(N__29839),
            .I(n2928));
    InMux I__4539 (
            .O(N__29832),
            .I(N__29828));
    CascadeMux I__4538 (
            .O(N__29831),
            .I(N__29824));
    LocalMux I__4537 (
            .O(N__29828),
            .I(N__29821));
    InMux I__4536 (
            .O(N__29827),
            .I(N__29818));
    InMux I__4535 (
            .O(N__29824),
            .I(N__29815));
    Span4Mux_h I__4534 (
            .O(N__29821),
            .I(N__29810));
    LocalMux I__4533 (
            .O(N__29818),
            .I(N__29810));
    LocalMux I__4532 (
            .O(N__29815),
            .I(n2821));
    Odrv4 I__4531 (
            .O(N__29810),
            .I(n2821));
    InMux I__4530 (
            .O(N__29805),
            .I(N__29802));
    LocalMux I__4529 (
            .O(N__29802),
            .I(N__29799));
    Span4Mux_h I__4528 (
            .O(N__29799),
            .I(N__29796));
    Odrv4 I__4527 (
            .O(N__29796),
            .I(n2888));
    InMux I__4526 (
            .O(N__29793),
            .I(N__29790));
    LocalMux I__4525 (
            .O(N__29790),
            .I(N__29787));
    Span4Mux_v I__4524 (
            .O(N__29787),
            .I(N__29784));
    Odrv4 I__4523 (
            .O(N__29784),
            .I(n2881));
    CascadeMux I__4522 (
            .O(N__29781),
            .I(N__29778));
    InMux I__4521 (
            .O(N__29778),
            .I(N__29775));
    LocalMux I__4520 (
            .O(N__29775),
            .I(N__29771));
    InMux I__4519 (
            .O(N__29774),
            .I(N__29768));
    Span4Mux_v I__4518 (
            .O(N__29771),
            .I(N__29762));
    LocalMux I__4517 (
            .O(N__29768),
            .I(N__29762));
    InMux I__4516 (
            .O(N__29767),
            .I(N__29759));
    Span4Mux_h I__4515 (
            .O(N__29762),
            .I(N__29756));
    LocalMux I__4514 (
            .O(N__29759),
            .I(n2814));
    Odrv4 I__4513 (
            .O(N__29756),
            .I(n2814));
    InMux I__4512 (
            .O(N__29751),
            .I(N__29748));
    LocalMux I__4511 (
            .O(N__29748),
            .I(N__29745));
    Span4Mux_v I__4510 (
            .O(N__29745),
            .I(N__29742));
    Odrv4 I__4509 (
            .O(N__29742),
            .I(n2893));
    CascadeMux I__4508 (
            .O(N__29739),
            .I(N__29736));
    InMux I__4507 (
            .O(N__29736),
            .I(N__29733));
    LocalMux I__4506 (
            .O(N__29733),
            .I(N__29729));
    CascadeMux I__4505 (
            .O(N__29732),
            .I(N__29726));
    Span4Mux_v I__4504 (
            .O(N__29729),
            .I(N__29723));
    InMux I__4503 (
            .O(N__29726),
            .I(N__29720));
    Odrv4 I__4502 (
            .O(N__29723),
            .I(n2826));
    LocalMux I__4501 (
            .O(N__29720),
            .I(n2826));
    CascadeMux I__4500 (
            .O(N__29715),
            .I(N__29712));
    InMux I__4499 (
            .O(N__29712),
            .I(N__29709));
    LocalMux I__4498 (
            .O(N__29709),
            .I(N__29705));
    InMux I__4497 (
            .O(N__29708),
            .I(N__29702));
    Span4Mux_v I__4496 (
            .O(N__29705),
            .I(N__29696));
    LocalMux I__4495 (
            .O(N__29702),
            .I(N__29696));
    InMux I__4494 (
            .O(N__29701),
            .I(N__29693));
    Odrv4 I__4493 (
            .O(N__29696),
            .I(n2925));
    LocalMux I__4492 (
            .O(N__29693),
            .I(n2925));
    CascadeMux I__4491 (
            .O(N__29688),
            .I(N__29685));
    InMux I__4490 (
            .O(N__29685),
            .I(N__29680));
    InMux I__4489 (
            .O(N__29684),
            .I(N__29677));
    InMux I__4488 (
            .O(N__29683),
            .I(N__29674));
    LocalMux I__4487 (
            .O(N__29680),
            .I(N__29671));
    LocalMux I__4486 (
            .O(N__29677),
            .I(N__29668));
    LocalMux I__4485 (
            .O(N__29674),
            .I(N__29665));
    Span4Mux_h I__4484 (
            .O(N__29671),
            .I(N__29662));
    Span12Mux_s4_h I__4483 (
            .O(N__29668),
            .I(N__29659));
    Span4Mux_h I__4482 (
            .O(N__29665),
            .I(N__29656));
    Odrv4 I__4481 (
            .O(N__29662),
            .I(n2615));
    Odrv12 I__4480 (
            .O(N__29659),
            .I(n2615));
    Odrv4 I__4479 (
            .O(N__29656),
            .I(n2615));
    CascadeMux I__4478 (
            .O(N__29649),
            .I(N__29645));
    InMux I__4477 (
            .O(N__29648),
            .I(N__29642));
    InMux I__4476 (
            .O(N__29645),
            .I(N__29639));
    LocalMux I__4475 (
            .O(N__29642),
            .I(N__29636));
    LocalMux I__4474 (
            .O(N__29639),
            .I(N__29632));
    Span4Mux_v I__4473 (
            .O(N__29636),
            .I(N__29629));
    InMux I__4472 (
            .O(N__29635),
            .I(N__29626));
    Span4Mux_s2_h I__4471 (
            .O(N__29632),
            .I(N__29623));
    Odrv4 I__4470 (
            .O(N__29629),
            .I(n2831));
    LocalMux I__4469 (
            .O(N__29626),
            .I(n2831));
    Odrv4 I__4468 (
            .O(N__29623),
            .I(n2831));
    CascadeMux I__4467 (
            .O(N__29616),
            .I(N__29613));
    InMux I__4466 (
            .O(N__29613),
            .I(N__29610));
    LocalMux I__4465 (
            .O(N__29610),
            .I(N__29607));
    Span4Mux_v I__4464 (
            .O(N__29607),
            .I(N__29604));
    Span4Mux_h I__4463 (
            .O(N__29604),
            .I(N__29601));
    Odrv4 I__4462 (
            .O(N__29601),
            .I(n2898));
    CascadeMux I__4461 (
            .O(N__29598),
            .I(N__29595));
    InMux I__4460 (
            .O(N__29595),
            .I(N__29592));
    LocalMux I__4459 (
            .O(N__29592),
            .I(N__29587));
    InMux I__4458 (
            .O(N__29591),
            .I(N__29582));
    InMux I__4457 (
            .O(N__29590),
            .I(N__29582));
    Span4Mux_v I__4456 (
            .O(N__29587),
            .I(N__29579));
    LocalMux I__4455 (
            .O(N__29582),
            .I(n2930));
    Odrv4 I__4454 (
            .O(N__29579),
            .I(n2930));
    InMux I__4453 (
            .O(N__29574),
            .I(N__29571));
    LocalMux I__4452 (
            .O(N__29571),
            .I(N__29568));
    Span4Mux_h I__4451 (
            .O(N__29568),
            .I(N__29565));
    Odrv4 I__4450 (
            .O(N__29565),
            .I(n2991));
    InMux I__4449 (
            .O(N__29562),
            .I(N__29558));
    InMux I__4448 (
            .O(N__29561),
            .I(N__29555));
    LocalMux I__4447 (
            .O(N__29558),
            .I(N__29552));
    LocalMux I__4446 (
            .O(N__29555),
            .I(n2924));
    Odrv4 I__4445 (
            .O(N__29552),
            .I(n2924));
    CascadeMux I__4444 (
            .O(N__29547),
            .I(n2513_cascade_));
    InMux I__4443 (
            .O(N__29544),
            .I(N__29541));
    LocalMux I__4442 (
            .O(N__29541),
            .I(N__29537));
    InMux I__4441 (
            .O(N__29540),
            .I(N__29534));
    Span4Mux_h I__4440 (
            .O(N__29537),
            .I(N__29530));
    LocalMux I__4439 (
            .O(N__29534),
            .I(N__29527));
    InMux I__4438 (
            .O(N__29533),
            .I(N__29524));
    Span4Mux_v I__4437 (
            .O(N__29530),
            .I(N__29521));
    Span4Mux_v I__4436 (
            .O(N__29527),
            .I(N__29516));
    LocalMux I__4435 (
            .O(N__29524),
            .I(N__29516));
    Span4Mux_v I__4434 (
            .O(N__29521),
            .I(N__29511));
    Span4Mux_h I__4433 (
            .O(N__29516),
            .I(N__29511));
    Odrv4 I__4432 (
            .O(N__29511),
            .I(n2612));
    CascadeMux I__4431 (
            .O(N__29508),
            .I(N__29505));
    InMux I__4430 (
            .O(N__29505),
            .I(N__29502));
    LocalMux I__4429 (
            .O(N__29502),
            .I(N__29497));
    InMux I__4428 (
            .O(N__29501),
            .I(N__29494));
    InMux I__4427 (
            .O(N__29500),
            .I(N__29491));
    Span4Mux_h I__4426 (
            .O(N__29497),
            .I(N__29488));
    LocalMux I__4425 (
            .O(N__29494),
            .I(N__29483));
    LocalMux I__4424 (
            .O(N__29491),
            .I(N__29483));
    Span4Mux_v I__4423 (
            .O(N__29488),
            .I(N__29480));
    Span4Mux_h I__4422 (
            .O(N__29483),
            .I(N__29475));
    Span4Mux_v I__4421 (
            .O(N__29480),
            .I(N__29475));
    Odrv4 I__4420 (
            .O(N__29475),
            .I(n2629));
    InMux I__4419 (
            .O(N__29472),
            .I(N__29469));
    LocalMux I__4418 (
            .O(N__29469),
            .I(N__29466));
    Span4Mux_v I__4417 (
            .O(N__29466),
            .I(N__29463));
    Odrv4 I__4416 (
            .O(N__29463),
            .I(n2899));
    CascadeMux I__4415 (
            .O(N__29460),
            .I(N__29457));
    InMux I__4414 (
            .O(N__29457),
            .I(N__29454));
    LocalMux I__4413 (
            .O(N__29454),
            .I(N__29450));
    InMux I__4412 (
            .O(N__29453),
            .I(N__29447));
    Span4Mux_s3_h I__4411 (
            .O(N__29450),
            .I(N__29444));
    LocalMux I__4410 (
            .O(N__29447),
            .I(n2832));
    Odrv4 I__4409 (
            .O(N__29444),
            .I(n2832));
    CascadeMux I__4408 (
            .O(N__29439),
            .I(N__29435));
    CascadeMux I__4407 (
            .O(N__29438),
            .I(N__29431));
    InMux I__4406 (
            .O(N__29435),
            .I(N__29428));
    InMux I__4405 (
            .O(N__29434),
            .I(N__29425));
    InMux I__4404 (
            .O(N__29431),
            .I(N__29422));
    LocalMux I__4403 (
            .O(N__29428),
            .I(N__29419));
    LocalMux I__4402 (
            .O(N__29425),
            .I(N__29416));
    LocalMux I__4401 (
            .O(N__29422),
            .I(N__29413));
    Span12Mux_s3_h I__4400 (
            .O(N__29419),
            .I(N__29410));
    Span4Mux_v I__4399 (
            .O(N__29416),
            .I(N__29407));
    Span4Mux_h I__4398 (
            .O(N__29413),
            .I(N__29404));
    Span12Mux_v I__4397 (
            .O(N__29410),
            .I(N__29401));
    Odrv4 I__4396 (
            .O(N__29407),
            .I(n2630));
    Odrv4 I__4395 (
            .O(N__29404),
            .I(n2630));
    Odrv12 I__4394 (
            .O(N__29401),
            .I(n2630));
    CascadeMux I__4393 (
            .O(N__29394),
            .I(N__29391));
    InMux I__4392 (
            .O(N__29391),
            .I(N__29388));
    LocalMux I__4391 (
            .O(N__29388),
            .I(N__29384));
    InMux I__4390 (
            .O(N__29387),
            .I(N__29380));
    Span4Mux_h I__4389 (
            .O(N__29384),
            .I(N__29377));
    InMux I__4388 (
            .O(N__29383),
            .I(N__29374));
    LocalMux I__4387 (
            .O(N__29380),
            .I(N__29371));
    Span4Mux_v I__4386 (
            .O(N__29377),
            .I(N__29368));
    LocalMux I__4385 (
            .O(N__29374),
            .I(N__29365));
    Span4Mux_h I__4384 (
            .O(N__29371),
            .I(N__29362));
    Span4Mux_v I__4383 (
            .O(N__29368),
            .I(N__29357));
    Span4Mux_h I__4382 (
            .O(N__29365),
            .I(N__29357));
    Odrv4 I__4381 (
            .O(N__29362),
            .I(n2620));
    Odrv4 I__4380 (
            .O(N__29357),
            .I(n2620));
    InMux I__4379 (
            .O(N__29352),
            .I(N__29349));
    LocalMux I__4378 (
            .O(N__29349),
            .I(N__29346));
    Span4Mux_v I__4377 (
            .O(N__29346),
            .I(N__29343));
    Odrv4 I__4376 (
            .O(N__29343),
            .I(n2901));
    InMux I__4375 (
            .O(N__29340),
            .I(N__29337));
    LocalMux I__4374 (
            .O(N__29337),
            .I(N__29333));
    CascadeMux I__4373 (
            .O(N__29336),
            .I(N__29330));
    Span4Mux_h I__4372 (
            .O(N__29333),
            .I(N__29326));
    InMux I__4371 (
            .O(N__29330),
            .I(N__29323));
    InMux I__4370 (
            .O(N__29329),
            .I(N__29320));
    Odrv4 I__4369 (
            .O(N__29326),
            .I(n2824));
    LocalMux I__4368 (
            .O(N__29323),
            .I(n2824));
    LocalMux I__4367 (
            .O(N__29320),
            .I(n2824));
    InMux I__4366 (
            .O(N__29313),
            .I(N__29310));
    LocalMux I__4365 (
            .O(N__29310),
            .I(N__29307));
    Span4Mux_h I__4364 (
            .O(N__29307),
            .I(N__29304));
    Odrv4 I__4363 (
            .O(N__29304),
            .I(n2891));
    InMux I__4362 (
            .O(N__29301),
            .I(N__29297));
    CascadeMux I__4361 (
            .O(N__29300),
            .I(N__29294));
    LocalMux I__4360 (
            .O(N__29297),
            .I(N__29291));
    InMux I__4359 (
            .O(N__29294),
            .I(N__29288));
    Span12Mux_s6_v I__4358 (
            .O(N__29291),
            .I(N__29283));
    LocalMux I__4357 (
            .O(N__29288),
            .I(N__29283));
    Odrv12 I__4356 (
            .O(N__29283),
            .I(n2923));
    CascadeMux I__4355 (
            .O(N__29280),
            .I(n2923_cascade_));
    InMux I__4354 (
            .O(N__29277),
            .I(N__29274));
    LocalMux I__4353 (
            .O(N__29274),
            .I(n14214));
    CascadeMux I__4352 (
            .O(N__29271),
            .I(n2533_cascade_));
    CascadeMux I__4351 (
            .O(N__29268),
            .I(N__29265));
    InMux I__4350 (
            .O(N__29265),
            .I(N__29262));
    LocalMux I__4349 (
            .O(N__29262),
            .I(n12063));
    CascadeMux I__4348 (
            .O(N__29259),
            .I(N__29256));
    InMux I__4347 (
            .O(N__29256),
            .I(N__29253));
    LocalMux I__4346 (
            .O(N__29253),
            .I(N__29249));
    InMux I__4345 (
            .O(N__29252),
            .I(N__29246));
    Span4Mux_h I__4344 (
            .O(N__29249),
            .I(N__29243));
    LocalMux I__4343 (
            .O(N__29246),
            .I(N__29240));
    Span4Mux_v I__4342 (
            .O(N__29243),
            .I(N__29236));
    Span12Mux_s4_h I__4341 (
            .O(N__29240),
            .I(N__29233));
    InMux I__4340 (
            .O(N__29239),
            .I(N__29230));
    Span4Mux_v I__4339 (
            .O(N__29236),
            .I(N__29227));
    Odrv12 I__4338 (
            .O(N__29233),
            .I(n2632));
    LocalMux I__4337 (
            .O(N__29230),
            .I(n2632));
    Odrv4 I__4336 (
            .O(N__29227),
            .I(n2632));
    InMux I__4335 (
            .O(N__29220),
            .I(N__29217));
    LocalMux I__4334 (
            .O(N__29217),
            .I(n14188));
    CascadeMux I__4333 (
            .O(N__29214),
            .I(n2515_cascade_));
    InMux I__4332 (
            .O(N__29211),
            .I(N__29208));
    LocalMux I__4331 (
            .O(N__29208),
            .I(N__29205));
    Odrv4 I__4330 (
            .O(N__29205),
            .I(n14117));
    CascadeMux I__4329 (
            .O(N__29202),
            .I(n14194_cascade_));
    CascadeMux I__4328 (
            .O(N__29199),
            .I(n2544_cascade_));
    CascadeMux I__4327 (
            .O(N__29196),
            .I(N__29192));
    InMux I__4326 (
            .O(N__29195),
            .I(N__29189));
    InMux I__4325 (
            .O(N__29192),
            .I(N__29186));
    LocalMux I__4324 (
            .O(N__29189),
            .I(N__29183));
    LocalMux I__4323 (
            .O(N__29186),
            .I(N__29179));
    Span4Mux_v I__4322 (
            .O(N__29183),
            .I(N__29176));
    InMux I__4321 (
            .O(N__29182),
            .I(N__29173));
    Span12Mux_v I__4320 (
            .O(N__29179),
            .I(N__29170));
    Odrv4 I__4319 (
            .O(N__29176),
            .I(n2631));
    LocalMux I__4318 (
            .O(N__29173),
            .I(n2631));
    Odrv12 I__4317 (
            .O(N__29170),
            .I(n2631));
    CascadeMux I__4316 (
            .O(N__29163),
            .I(n2417_cascade_));
    InMux I__4315 (
            .O(N__29160),
            .I(N__29157));
    LocalMux I__4314 (
            .O(N__29157),
            .I(n14634));
    CascadeMux I__4313 (
            .O(N__29154),
            .I(n14640_cascade_));
    CascadeMux I__4312 (
            .O(N__29151),
            .I(n2445_cascade_));
    CascadeMux I__4311 (
            .O(N__29148),
            .I(n2530_cascade_));
    InMux I__4310 (
            .O(N__29145),
            .I(N__29142));
    LocalMux I__4309 (
            .O(N__29142),
            .I(n14646));
    CascadeMux I__4308 (
            .O(N__29139),
            .I(n2430_cascade_));
    InMux I__4307 (
            .O(N__29136),
            .I(N__29133));
    LocalMux I__4306 (
            .O(N__29133),
            .I(N__29130));
    Span4Mux_v I__4305 (
            .O(N__29130),
            .I(N__29127));
    Odrv4 I__4304 (
            .O(N__29127),
            .I(n2400));
    CascadeMux I__4303 (
            .O(N__29124),
            .I(N__29120));
    CascadeMux I__4302 (
            .O(N__29123),
            .I(N__29117));
    InMux I__4301 (
            .O(N__29120),
            .I(N__29114));
    InMux I__4300 (
            .O(N__29117),
            .I(N__29111));
    LocalMux I__4299 (
            .O(N__29114),
            .I(N__29108));
    LocalMux I__4298 (
            .O(N__29111),
            .I(N__29105));
    Span4Mux_v I__4297 (
            .O(N__29108),
            .I(N__29101));
    Span4Mux_s2_h I__4296 (
            .O(N__29105),
            .I(N__29098));
    InMux I__4295 (
            .O(N__29104),
            .I(N__29095));
    Odrv4 I__4294 (
            .O(N__29101),
            .I(n2333));
    Odrv4 I__4293 (
            .O(N__29098),
            .I(n2333));
    LocalMux I__4292 (
            .O(N__29095),
            .I(n2333));
    CascadeMux I__4291 (
            .O(N__29088),
            .I(n2432_cascade_));
    InMux I__4290 (
            .O(N__29085),
            .I(N__29082));
    LocalMux I__4289 (
            .O(N__29082),
            .I(n11967));
    CascadeMux I__4288 (
            .O(N__29079),
            .I(n2528_cascade_));
    CascadeMux I__4287 (
            .O(N__29076),
            .I(N__29073));
    InMux I__4286 (
            .O(N__29073),
            .I(N__29070));
    LocalMux I__4285 (
            .O(N__29070),
            .I(N__29066));
    InMux I__4284 (
            .O(N__29069),
            .I(N__29063));
    Span4Mux_h I__4283 (
            .O(N__29066),
            .I(N__29060));
    LocalMux I__4282 (
            .O(N__29063),
            .I(N__29056));
    Span4Mux_v I__4281 (
            .O(N__29060),
            .I(N__29053));
    InMux I__4280 (
            .O(N__29059),
            .I(N__29050));
    Span4Mux_h I__4279 (
            .O(N__29056),
            .I(N__29045));
    Span4Mux_v I__4278 (
            .O(N__29053),
            .I(N__29045));
    LocalMux I__4277 (
            .O(N__29050),
            .I(n2627));
    Odrv4 I__4276 (
            .O(N__29045),
            .I(n2627));
    InMux I__4275 (
            .O(N__29040),
            .I(N__29037));
    LocalMux I__4274 (
            .O(N__29037),
            .I(N__29034));
    Span4Mux_h I__4273 (
            .O(N__29034),
            .I(N__29031));
    Odrv4 I__4272 (
            .O(N__29031),
            .I(n2384));
    CascadeMux I__4271 (
            .O(N__29028),
            .I(N__29025));
    InMux I__4270 (
            .O(N__29025),
            .I(N__29021));
    InMux I__4269 (
            .O(N__29024),
            .I(N__29018));
    LocalMux I__4268 (
            .O(N__29021),
            .I(N__29014));
    LocalMux I__4267 (
            .O(N__29018),
            .I(N__29011));
    CascadeMux I__4266 (
            .O(N__29017),
            .I(N__29008));
    Span4Mux_h I__4265 (
            .O(N__29014),
            .I(N__29005));
    Span4Mux_s3_h I__4264 (
            .O(N__29011),
            .I(N__29002));
    InMux I__4263 (
            .O(N__29008),
            .I(N__28999));
    Odrv4 I__4262 (
            .O(N__29005),
            .I(n2317));
    Odrv4 I__4261 (
            .O(N__29002),
            .I(n2317));
    LocalMux I__4260 (
            .O(N__28999),
            .I(n2317));
    InMux I__4259 (
            .O(N__28992),
            .I(N__28989));
    LocalMux I__4258 (
            .O(N__28989),
            .I(n13828));
    InMux I__4257 (
            .O(N__28986),
            .I(N__28983));
    LocalMux I__4256 (
            .O(N__28983),
            .I(n14628));
    InMux I__4255 (
            .O(N__28980),
            .I(N__28976));
    InMux I__4254 (
            .O(N__28979),
            .I(N__28973));
    LocalMux I__4253 (
            .O(N__28976),
            .I(N__28969));
    LocalMux I__4252 (
            .O(N__28973),
            .I(N__28966));
    InMux I__4251 (
            .O(N__28972),
            .I(N__28963));
    Span4Mux_v I__4250 (
            .O(N__28969),
            .I(N__28960));
    Span4Mux_s2_h I__4249 (
            .O(N__28966),
            .I(N__28957));
    LocalMux I__4248 (
            .O(N__28963),
            .I(N__28954));
    Odrv4 I__4247 (
            .O(N__28960),
            .I(n2318));
    Odrv4 I__4246 (
            .O(N__28957),
            .I(n2318));
    Odrv4 I__4245 (
            .O(N__28954),
            .I(n2318));
    CascadeMux I__4244 (
            .O(N__28947),
            .I(N__28944));
    InMux I__4243 (
            .O(N__28944),
            .I(N__28941));
    LocalMux I__4242 (
            .O(N__28941),
            .I(N__28938));
    Span4Mux_h I__4241 (
            .O(N__28938),
            .I(N__28935));
    Odrv4 I__4240 (
            .O(N__28935),
            .I(n2385));
    InMux I__4239 (
            .O(N__28932),
            .I(N__28929));
    LocalMux I__4238 (
            .O(N__28929),
            .I(N__28926));
    Odrv12 I__4237 (
            .O(N__28926),
            .I(n2390));
    CascadeMux I__4236 (
            .O(N__28923),
            .I(N__28919));
    CascadeMux I__4235 (
            .O(N__28922),
            .I(N__28916));
    InMux I__4234 (
            .O(N__28919),
            .I(N__28913));
    InMux I__4233 (
            .O(N__28916),
            .I(N__28910));
    LocalMux I__4232 (
            .O(N__28913),
            .I(N__28907));
    LocalMux I__4231 (
            .O(N__28910),
            .I(N__28904));
    Span4Mux_v I__4230 (
            .O(N__28907),
            .I(N__28899));
    Span4Mux_v I__4229 (
            .O(N__28904),
            .I(N__28899));
    Odrv4 I__4228 (
            .O(N__28899),
            .I(n2323));
    CascadeMux I__4227 (
            .O(N__28896),
            .I(N__28892));
    InMux I__4226 (
            .O(N__28895),
            .I(N__28888));
    InMux I__4225 (
            .O(N__28892),
            .I(N__28885));
    InMux I__4224 (
            .O(N__28891),
            .I(N__28882));
    LocalMux I__4223 (
            .O(N__28888),
            .I(N__28879));
    LocalMux I__4222 (
            .O(N__28885),
            .I(n2118));
    LocalMux I__4221 (
            .O(N__28882),
            .I(n2118));
    Odrv4 I__4220 (
            .O(N__28879),
            .I(n2118));
    InMux I__4219 (
            .O(N__28872),
            .I(N__28869));
    LocalMux I__4218 (
            .O(N__28869),
            .I(N__28866));
    Odrv12 I__4217 (
            .O(N__28866),
            .I(n2393));
    CascadeMux I__4216 (
            .O(N__28863),
            .I(N__28860));
    InMux I__4215 (
            .O(N__28860),
            .I(N__28856));
    CascadeMux I__4214 (
            .O(N__28859),
            .I(N__28853));
    LocalMux I__4213 (
            .O(N__28856),
            .I(N__28850));
    InMux I__4212 (
            .O(N__28853),
            .I(N__28846));
    Span4Mux_v I__4211 (
            .O(N__28850),
            .I(N__28843));
    InMux I__4210 (
            .O(N__28849),
            .I(N__28840));
    LocalMux I__4209 (
            .O(N__28846),
            .I(n2326));
    Odrv4 I__4208 (
            .O(N__28843),
            .I(n2326));
    LocalMux I__4207 (
            .O(N__28840),
            .I(n2326));
    InMux I__4206 (
            .O(N__28833),
            .I(N__28828));
    CascadeMux I__4205 (
            .O(N__28832),
            .I(N__28825));
    CascadeMux I__4204 (
            .O(N__28831),
            .I(N__28822));
    LocalMux I__4203 (
            .O(N__28828),
            .I(N__28819));
    InMux I__4202 (
            .O(N__28825),
            .I(N__28816));
    InMux I__4201 (
            .O(N__28822),
            .I(N__28813));
    Span4Mux_v I__4200 (
            .O(N__28819),
            .I(N__28808));
    LocalMux I__4199 (
            .O(N__28816),
            .I(N__28808));
    LocalMux I__4198 (
            .O(N__28813),
            .I(n2330));
    Odrv4 I__4197 (
            .O(N__28808),
            .I(n2330));
    InMux I__4196 (
            .O(N__28803),
            .I(N__28800));
    LocalMux I__4195 (
            .O(N__28800),
            .I(N__28797));
    Span12Mux_v I__4194 (
            .O(N__28797),
            .I(N__28794));
    Odrv12 I__4193 (
            .O(N__28794),
            .I(n2397));
    CascadeMux I__4192 (
            .O(N__28791),
            .I(N__28787));
    InMux I__4191 (
            .O(N__28790),
            .I(N__28784));
    InMux I__4190 (
            .O(N__28787),
            .I(N__28781));
    LocalMux I__4189 (
            .O(N__28784),
            .I(N__28778));
    LocalMux I__4188 (
            .O(N__28781),
            .I(N__28775));
    Span4Mux_h I__4187 (
            .O(N__28778),
            .I(N__28769));
    Span4Mux_s2_h I__4186 (
            .O(N__28775),
            .I(N__28769));
    InMux I__4185 (
            .O(N__28774),
            .I(N__28766));
    Odrv4 I__4184 (
            .O(N__28769),
            .I(n2322));
    LocalMux I__4183 (
            .O(N__28766),
            .I(n2322));
    CascadeMux I__4182 (
            .O(N__28761),
            .I(N__28758));
    InMux I__4181 (
            .O(N__28758),
            .I(N__28755));
    LocalMux I__4180 (
            .O(N__28755),
            .I(N__28752));
    Odrv12 I__4179 (
            .O(N__28752),
            .I(n2389));
    InMux I__4178 (
            .O(N__28749),
            .I(N__28746));
    LocalMux I__4177 (
            .O(N__28746),
            .I(N__28743));
    Span4Mux_v I__4176 (
            .O(N__28743),
            .I(N__28740));
    Odrv4 I__4175 (
            .O(N__28740),
            .I(n2399));
    CascadeMux I__4174 (
            .O(N__28737),
            .I(N__28733));
    InMux I__4173 (
            .O(N__28736),
            .I(N__28730));
    InMux I__4172 (
            .O(N__28733),
            .I(N__28727));
    LocalMux I__4171 (
            .O(N__28730),
            .I(N__28724));
    LocalMux I__4170 (
            .O(N__28727),
            .I(N__28721));
    Span4Mux_v I__4169 (
            .O(N__28724),
            .I(N__28717));
    Span4Mux_s2_h I__4168 (
            .O(N__28721),
            .I(N__28714));
    InMux I__4167 (
            .O(N__28720),
            .I(N__28711));
    Odrv4 I__4166 (
            .O(N__28717),
            .I(n2332));
    Odrv4 I__4165 (
            .O(N__28714),
            .I(n2332));
    LocalMux I__4164 (
            .O(N__28711),
            .I(n2332));
    InMux I__4163 (
            .O(N__28704),
            .I(N__28701));
    LocalMux I__4162 (
            .O(N__28701),
            .I(N__28698));
    Span4Mux_v I__4161 (
            .O(N__28698),
            .I(N__28695));
    Odrv4 I__4160 (
            .O(N__28695),
            .I(n2388));
    CascadeMux I__4159 (
            .O(N__28692),
            .I(N__28689));
    InMux I__4158 (
            .O(N__28689),
            .I(N__28685));
    InMux I__4157 (
            .O(N__28688),
            .I(N__28682));
    LocalMux I__4156 (
            .O(N__28685),
            .I(N__28678));
    LocalMux I__4155 (
            .O(N__28682),
            .I(N__28675));
    InMux I__4154 (
            .O(N__28681),
            .I(N__28672));
    Span4Mux_v I__4153 (
            .O(N__28678),
            .I(N__28669));
    Span4Mux_s3_h I__4152 (
            .O(N__28675),
            .I(N__28664));
    LocalMux I__4151 (
            .O(N__28672),
            .I(N__28664));
    Odrv4 I__4150 (
            .O(N__28669),
            .I(n2321));
    Odrv4 I__4149 (
            .O(N__28664),
            .I(n2321));
    CascadeMux I__4148 (
            .O(N__28659),
            .I(n2420_cascade_));
    InMux I__4147 (
            .O(N__28656),
            .I(N__28653));
    LocalMux I__4146 (
            .O(N__28653),
            .I(n14622));
    InMux I__4145 (
            .O(N__28650),
            .I(N__28647));
    LocalMux I__4144 (
            .O(N__28647),
            .I(N__28644));
    Span4Mux_v I__4143 (
            .O(N__28644),
            .I(N__28641));
    Odrv4 I__4142 (
            .O(N__28641),
            .I(n2398));
    CascadeMux I__4141 (
            .O(N__28638),
            .I(N__28634));
    CascadeMux I__4140 (
            .O(N__28637),
            .I(N__28631));
    InMux I__4139 (
            .O(N__28634),
            .I(N__28628));
    InMux I__4138 (
            .O(N__28631),
            .I(N__28625));
    LocalMux I__4137 (
            .O(N__28628),
            .I(N__28622));
    LocalMux I__4136 (
            .O(N__28625),
            .I(N__28619));
    Span4Mux_v I__4135 (
            .O(N__28622),
            .I(N__28614));
    Span4Mux_v I__4134 (
            .O(N__28619),
            .I(N__28614));
    Odrv4 I__4133 (
            .O(N__28614),
            .I(n2331));
    CascadeMux I__4132 (
            .O(N__28611),
            .I(N__28608));
    InMux I__4131 (
            .O(N__28608),
            .I(N__28604));
    CascadeMux I__4130 (
            .O(N__28607),
            .I(N__28601));
    LocalMux I__4129 (
            .O(N__28604),
            .I(N__28597));
    InMux I__4128 (
            .O(N__28601),
            .I(N__28594));
    InMux I__4127 (
            .O(N__28600),
            .I(N__28591));
    Odrv4 I__4126 (
            .O(N__28597),
            .I(n2126));
    LocalMux I__4125 (
            .O(N__28594),
            .I(n2126));
    LocalMux I__4124 (
            .O(N__28591),
            .I(n2126));
    CascadeMux I__4123 (
            .O(N__28584),
            .I(n2128_cascade_));
    InMux I__4122 (
            .O(N__28581),
            .I(N__28578));
    LocalMux I__4121 (
            .O(N__28578),
            .I(n14316));
    CascadeMux I__4120 (
            .O(N__28575),
            .I(N__28570));
    CascadeMux I__4119 (
            .O(N__28574),
            .I(N__28567));
    InMux I__4118 (
            .O(N__28573),
            .I(N__28564));
    InMux I__4117 (
            .O(N__28570),
            .I(N__28561));
    InMux I__4116 (
            .O(N__28567),
            .I(N__28558));
    LocalMux I__4115 (
            .O(N__28564),
            .I(N__28555));
    LocalMux I__4114 (
            .O(N__28561),
            .I(n2125));
    LocalMux I__4113 (
            .O(N__28558),
            .I(n2125));
    Odrv4 I__4112 (
            .O(N__28555),
            .I(n2125));
    InMux I__4111 (
            .O(N__28548),
            .I(N__28545));
    LocalMux I__4110 (
            .O(N__28545),
            .I(N__28542));
    Odrv4 I__4109 (
            .O(N__28542),
            .I(n2185));
    CascadeMux I__4108 (
            .O(N__28539),
            .I(N__28536));
    InMux I__4107 (
            .O(N__28536),
            .I(N__28532));
    CascadeMux I__4106 (
            .O(N__28535),
            .I(N__28528));
    LocalMux I__4105 (
            .O(N__28532),
            .I(N__28525));
    InMux I__4104 (
            .O(N__28531),
            .I(N__28522));
    InMux I__4103 (
            .O(N__28528),
            .I(N__28519));
    Span4Mux_h I__4102 (
            .O(N__28525),
            .I(N__28516));
    LocalMux I__4101 (
            .O(N__28522),
            .I(N__28513));
    LocalMux I__4100 (
            .O(N__28519),
            .I(n2217));
    Odrv4 I__4099 (
            .O(N__28516),
            .I(n2217));
    Odrv4 I__4098 (
            .O(N__28513),
            .I(n2217));
    InMux I__4097 (
            .O(N__28506),
            .I(N__28503));
    LocalMux I__4096 (
            .O(N__28503),
            .I(n2183));
    InMux I__4095 (
            .O(N__28500),
            .I(N__28496));
    InMux I__4094 (
            .O(N__28499),
            .I(N__28493));
    LocalMux I__4093 (
            .O(N__28496),
            .I(n2116));
    LocalMux I__4092 (
            .O(N__28493),
            .I(n2116));
    InMux I__4091 (
            .O(N__28488),
            .I(N__28485));
    LocalMux I__4090 (
            .O(N__28485),
            .I(N__28480));
    InMux I__4089 (
            .O(N__28484),
            .I(N__28477));
    InMux I__4088 (
            .O(N__28483),
            .I(N__28474));
    Span4Mux_h I__4087 (
            .O(N__28480),
            .I(N__28471));
    LocalMux I__4086 (
            .O(N__28477),
            .I(N__28468));
    LocalMux I__4085 (
            .O(N__28474),
            .I(n2215));
    Odrv4 I__4084 (
            .O(N__28471),
            .I(n2215));
    Odrv4 I__4083 (
            .O(N__28468),
            .I(n2215));
    InMux I__4082 (
            .O(N__28461),
            .I(N__28458));
    LocalMux I__4081 (
            .O(N__28458),
            .I(n2184));
    InMux I__4080 (
            .O(N__28455),
            .I(N__28452));
    LocalMux I__4079 (
            .O(N__28452),
            .I(N__28447));
    CascadeMux I__4078 (
            .O(N__28451),
            .I(N__28444));
    InMux I__4077 (
            .O(N__28450),
            .I(N__28441));
    Span4Mux_v I__4076 (
            .O(N__28447),
            .I(N__28438));
    InMux I__4075 (
            .O(N__28444),
            .I(N__28435));
    LocalMux I__4074 (
            .O(N__28441),
            .I(N__28432));
    Odrv4 I__4073 (
            .O(N__28438),
            .I(n2122));
    LocalMux I__4072 (
            .O(N__28435),
            .I(n2122));
    Odrv4 I__4071 (
            .O(N__28432),
            .I(n2122));
    CascadeMux I__4070 (
            .O(N__28425),
            .I(N__28422));
    InMux I__4069 (
            .O(N__28422),
            .I(N__28417));
    InMux I__4068 (
            .O(N__28421),
            .I(N__28412));
    InMux I__4067 (
            .O(N__28420),
            .I(N__28412));
    LocalMux I__4066 (
            .O(N__28417),
            .I(n2124));
    LocalMux I__4065 (
            .O(N__28412),
            .I(n2124));
    InMux I__4064 (
            .O(N__28407),
            .I(N__28404));
    LocalMux I__4063 (
            .O(N__28404),
            .I(N__28401));
    Span4Mux_h I__4062 (
            .O(N__28401),
            .I(N__28398));
    Odrv4 I__4061 (
            .O(N__28398),
            .I(n2401));
    InMux I__4060 (
            .O(N__28395),
            .I(N__28392));
    LocalMux I__4059 (
            .O(N__28392),
            .I(n2198));
    CascadeMux I__4058 (
            .O(N__28389),
            .I(n2131_cascade_));
    CascadeMux I__4057 (
            .O(N__28386),
            .I(N__28381));
    InMux I__4056 (
            .O(N__28385),
            .I(N__28376));
    InMux I__4055 (
            .O(N__28384),
            .I(N__28376));
    InMux I__4054 (
            .O(N__28381),
            .I(N__28373));
    LocalMux I__4053 (
            .O(N__28376),
            .I(N__28370));
    LocalMux I__4052 (
            .O(N__28373),
            .I(N__28367));
    Span4Mux_h I__4051 (
            .O(N__28370),
            .I(N__28364));
    Span4Mux_h I__4050 (
            .O(N__28367),
            .I(N__28361));
    Odrv4 I__4049 (
            .O(N__28364),
            .I(n2230));
    Odrv4 I__4048 (
            .O(N__28361),
            .I(n2230));
    InMux I__4047 (
            .O(N__28356),
            .I(N__28353));
    LocalMux I__4046 (
            .O(N__28353),
            .I(n14584));
    CascadeMux I__4045 (
            .O(N__28350),
            .I(N__28347));
    InMux I__4044 (
            .O(N__28347),
            .I(N__28344));
    LocalMux I__4043 (
            .O(N__28344),
            .I(n2191));
    CascadeMux I__4042 (
            .O(N__28341),
            .I(N__28337));
    CascadeMux I__4041 (
            .O(N__28340),
            .I(N__28333));
    InMux I__4040 (
            .O(N__28337),
            .I(N__28330));
    InMux I__4039 (
            .O(N__28336),
            .I(N__28327));
    InMux I__4038 (
            .O(N__28333),
            .I(N__28324));
    LocalMux I__4037 (
            .O(N__28330),
            .I(N__28319));
    LocalMux I__4036 (
            .O(N__28327),
            .I(N__28319));
    LocalMux I__4035 (
            .O(N__28324),
            .I(N__28314));
    Span4Mux_v I__4034 (
            .O(N__28319),
            .I(N__28314));
    Odrv4 I__4033 (
            .O(N__28314),
            .I(n2223));
    InMux I__4032 (
            .O(N__28311),
            .I(N__28308));
    LocalMux I__4031 (
            .O(N__28308),
            .I(n2192));
    CascadeMux I__4030 (
            .O(N__28305),
            .I(N__28301));
    CascadeMux I__4029 (
            .O(N__28304),
            .I(N__28298));
    InMux I__4028 (
            .O(N__28301),
            .I(N__28295));
    InMux I__4027 (
            .O(N__28298),
            .I(N__28292));
    LocalMux I__4026 (
            .O(N__28295),
            .I(N__28289));
    LocalMux I__4025 (
            .O(N__28292),
            .I(N__28285));
    Span4Mux_h I__4024 (
            .O(N__28289),
            .I(N__28282));
    InMux I__4023 (
            .O(N__28288),
            .I(N__28279));
    Odrv4 I__4022 (
            .O(N__28285),
            .I(n2224));
    Odrv4 I__4021 (
            .O(N__28282),
            .I(n2224));
    LocalMux I__4020 (
            .O(N__28279),
            .I(n2224));
    InMux I__4019 (
            .O(N__28272),
            .I(N__28269));
    LocalMux I__4018 (
            .O(N__28269),
            .I(n14330));
    CascadeMux I__4017 (
            .O(N__28266),
            .I(n2116_cascade_));
    CascadeMux I__4016 (
            .O(N__28263),
            .I(n2148_cascade_));
    InMux I__4015 (
            .O(N__28260),
            .I(N__28257));
    LocalMux I__4014 (
            .O(N__28257),
            .I(n2195));
    CascadeMux I__4013 (
            .O(N__28254),
            .I(N__28251));
    InMux I__4012 (
            .O(N__28251),
            .I(N__28248));
    LocalMux I__4011 (
            .O(N__28248),
            .I(N__28243));
    CascadeMux I__4010 (
            .O(N__28247),
            .I(N__28240));
    InMux I__4009 (
            .O(N__28246),
            .I(N__28237));
    Span4Mux_h I__4008 (
            .O(N__28243),
            .I(N__28234));
    InMux I__4007 (
            .O(N__28240),
            .I(N__28231));
    LocalMux I__4006 (
            .O(N__28237),
            .I(n2227));
    Odrv4 I__4005 (
            .O(N__28234),
            .I(n2227));
    LocalMux I__4004 (
            .O(N__28231),
            .I(n2227));
    CascadeMux I__4003 (
            .O(N__28224),
            .I(N__28220));
    InMux I__4002 (
            .O(N__28223),
            .I(N__28217));
    InMux I__4001 (
            .O(N__28220),
            .I(N__28214));
    LocalMux I__4000 (
            .O(N__28217),
            .I(n2128));
    LocalMux I__3999 (
            .O(N__28214),
            .I(n2128));
    InMux I__3998 (
            .O(N__28209),
            .I(N__28205));
    InMux I__3997 (
            .O(N__28208),
            .I(N__28202));
    LocalMux I__3996 (
            .O(N__28205),
            .I(N__28197));
    LocalMux I__3995 (
            .O(N__28202),
            .I(N__28197));
    Span4Mux_s3_v I__3994 (
            .O(N__28197),
            .I(N__28193));
    InMux I__3993 (
            .O(N__28196),
            .I(N__28190));
    Odrv4 I__3992 (
            .O(N__28193),
            .I(n3010));
    LocalMux I__3991 (
            .O(N__28190),
            .I(n3010));
    CascadeMux I__3990 (
            .O(N__28185),
            .I(N__28182));
    InMux I__3989 (
            .O(N__28182),
            .I(N__28179));
    LocalMux I__3988 (
            .O(N__28179),
            .I(n3077));
    InMux I__3987 (
            .O(N__28176),
            .I(N__28173));
    LocalMux I__3986 (
            .O(N__28173),
            .I(N__28170));
    Odrv4 I__3985 (
            .O(N__28170),
            .I(n14264));
    CascadeMux I__3984 (
            .O(N__28167),
            .I(N__28164));
    InMux I__3983 (
            .O(N__28164),
            .I(N__28161));
    LocalMux I__3982 (
            .O(N__28161),
            .I(N__28158));
    Odrv4 I__3981 (
            .O(N__28158),
            .I(n14260));
    CascadeMux I__3980 (
            .O(N__28155),
            .I(N__28152));
    InMux I__3979 (
            .O(N__28152),
            .I(N__28147));
    InMux I__3978 (
            .O(N__28151),
            .I(N__28142));
    InMux I__3977 (
            .O(N__28150),
            .I(N__28142));
    LocalMux I__3976 (
            .O(N__28147),
            .I(n2130));
    LocalMux I__3975 (
            .O(N__28142),
            .I(n2130));
    CascadeMux I__3974 (
            .O(N__28137),
            .I(n14324_cascade_));
    InMux I__3973 (
            .O(N__28134),
            .I(N__28131));
    LocalMux I__3972 (
            .O(N__28131),
            .I(n13787));
    CascadeMux I__3971 (
            .O(N__28128),
            .I(N__28124));
    CascadeMux I__3970 (
            .O(N__28127),
            .I(N__28121));
    InMux I__3969 (
            .O(N__28124),
            .I(N__28118));
    InMux I__3968 (
            .O(N__28121),
            .I(N__28115));
    LocalMux I__3967 (
            .O(N__28118),
            .I(n2127));
    LocalMux I__3966 (
            .O(N__28115),
            .I(n2127));
    CascadeMux I__3965 (
            .O(N__28110),
            .I(n2127_cascade_));
    InMux I__3964 (
            .O(N__28107),
            .I(N__28104));
    LocalMux I__3963 (
            .O(N__28104),
            .I(n14318));
    CascadeMux I__3962 (
            .O(N__28101),
            .I(N__28098));
    InMux I__3961 (
            .O(N__28098),
            .I(N__28094));
    InMux I__3960 (
            .O(N__28097),
            .I(N__28091));
    LocalMux I__3959 (
            .O(N__28094),
            .I(n2131));
    LocalMux I__3958 (
            .O(N__28091),
            .I(n2131));
    CascadeMux I__3957 (
            .O(N__28086),
            .I(n3212_cascade_));
    InMux I__3956 (
            .O(N__28083),
            .I(N__28080));
    LocalMux I__3955 (
            .O(N__28080),
            .I(n14798));
    InMux I__3954 (
            .O(N__28077),
            .I(N__28072));
    InMux I__3953 (
            .O(N__28076),
            .I(N__28069));
    InMux I__3952 (
            .O(N__28075),
            .I(N__28066));
    LocalMux I__3951 (
            .O(N__28072),
            .I(n3107));
    LocalMux I__3950 (
            .O(N__28069),
            .I(n3107));
    LocalMux I__3949 (
            .O(N__28066),
            .I(n3107));
    InMux I__3948 (
            .O(N__28059),
            .I(N__28054));
    InMux I__3947 (
            .O(N__28058),
            .I(N__28051));
    InMux I__3946 (
            .O(N__28057),
            .I(N__28048));
    LocalMux I__3945 (
            .O(N__28054),
            .I(n3106));
    LocalMux I__3944 (
            .O(N__28051),
            .I(n3106));
    LocalMux I__3943 (
            .O(N__28048),
            .I(n3106));
    CascadeMux I__3942 (
            .O(N__28041),
            .I(N__28037));
    InMux I__3941 (
            .O(N__28040),
            .I(N__28034));
    InMux I__3940 (
            .O(N__28037),
            .I(N__28031));
    LocalMux I__3939 (
            .O(N__28034),
            .I(n3105));
    LocalMux I__3938 (
            .O(N__28031),
            .I(n3105));
    InMux I__3937 (
            .O(N__28026),
            .I(N__28023));
    LocalMux I__3936 (
            .O(N__28023),
            .I(N__28020));
    Span4Mux_h I__3935 (
            .O(N__28020),
            .I(N__28017));
    Odrv4 I__3934 (
            .O(N__28017),
            .I(n3195));
    CascadeMux I__3933 (
            .O(N__28014),
            .I(n3138_cascade_));
    InMux I__3932 (
            .O(N__28011),
            .I(N__28008));
    LocalMux I__3931 (
            .O(N__28008),
            .I(N__28004));
    CascadeMux I__3930 (
            .O(N__28007),
            .I(N__28001));
    Span4Mux_h I__3929 (
            .O(N__28004),
            .I(N__27998));
    InMux I__3928 (
            .O(N__28001),
            .I(N__27995));
    Odrv4 I__3927 (
            .O(N__27998),
            .I(n3128));
    LocalMux I__3926 (
            .O(N__27995),
            .I(n3128));
    CascadeMux I__3925 (
            .O(N__27990),
            .I(N__27987));
    InMux I__3924 (
            .O(N__27987),
            .I(N__27984));
    LocalMux I__3923 (
            .O(N__27984),
            .I(N__27981));
    Odrv4 I__3922 (
            .O(N__27981),
            .I(n3181));
    InMux I__3921 (
            .O(N__27978),
            .I(N__27975));
    LocalMux I__3920 (
            .O(N__27975),
            .I(N__27972));
    Odrv4 I__3919 (
            .O(N__27972),
            .I(n3184));
    InMux I__3918 (
            .O(N__27969),
            .I(N__27964));
    InMux I__3917 (
            .O(N__27968),
            .I(N__27961));
    InMux I__3916 (
            .O(N__27967),
            .I(N__27958));
    LocalMux I__3915 (
            .O(N__27964),
            .I(N__27955));
    LocalMux I__3914 (
            .O(N__27961),
            .I(N__27952));
    LocalMux I__3913 (
            .O(N__27958),
            .I(N__27949));
    Span4Mux_s3_v I__3912 (
            .O(N__27955),
            .I(N__27944));
    Span4Mux_v I__3911 (
            .O(N__27952),
            .I(N__27944));
    Odrv4 I__3910 (
            .O(N__27949),
            .I(n3117));
    Odrv4 I__3909 (
            .O(N__27944),
            .I(n3117));
    CascadeMux I__3908 (
            .O(N__27939),
            .I(N__27936));
    InMux I__3907 (
            .O(N__27936),
            .I(N__27933));
    LocalMux I__3906 (
            .O(N__27933),
            .I(N__27930));
    Span4Mux_s2_v I__3905 (
            .O(N__27930),
            .I(N__27927));
    Odrv4 I__3904 (
            .O(N__27927),
            .I(n3083));
    InMux I__3903 (
            .O(N__27924),
            .I(N__27921));
    LocalMux I__3902 (
            .O(N__27921),
            .I(N__27918));
    Odrv4 I__3901 (
            .O(N__27918),
            .I(n13831));
    InMux I__3900 (
            .O(N__27915),
            .I(N__27910));
    InMux I__3899 (
            .O(N__27914),
            .I(N__27907));
    InMux I__3898 (
            .O(N__27913),
            .I(N__27904));
    LocalMux I__3897 (
            .O(N__27910),
            .I(n3114));
    LocalMux I__3896 (
            .O(N__27907),
            .I(n3114));
    LocalMux I__3895 (
            .O(N__27904),
            .I(n3114));
    CascadeMux I__3894 (
            .O(N__27897),
            .I(n3115_cascade_));
    InMux I__3893 (
            .O(N__27894),
            .I(N__27891));
    LocalMux I__3892 (
            .O(N__27891),
            .I(N__27888));
    Span4Mux_v I__3891 (
            .O(N__27888),
            .I(N__27885));
    Odrv4 I__3890 (
            .O(N__27885),
            .I(n14156));
    InMux I__3889 (
            .O(N__27882),
            .I(N__27878));
    InMux I__3888 (
            .O(N__27881),
            .I(N__27874));
    LocalMux I__3887 (
            .O(N__27878),
            .I(N__27871));
    InMux I__3886 (
            .O(N__27877),
            .I(N__27868));
    LocalMux I__3885 (
            .O(N__27874),
            .I(N__27863));
    Span4Mux_s3_h I__3884 (
            .O(N__27871),
            .I(N__27863));
    LocalMux I__3883 (
            .O(N__27868),
            .I(N__27860));
    Span4Mux_v I__3882 (
            .O(N__27863),
            .I(N__27857));
    Span12Mux_s2_v I__3881 (
            .O(N__27860),
            .I(N__27854));
    Odrv4 I__3880 (
            .O(N__27857),
            .I(n3113));
    Odrv12 I__3879 (
            .O(N__27854),
            .I(n3113));
    CascadeMux I__3878 (
            .O(N__27849),
            .I(n14162_cascade_));
    CascadeMux I__3877 (
            .O(N__27846),
            .I(n14168_cascade_));
    InMux I__3876 (
            .O(N__27843),
            .I(N__27839));
    InMux I__3875 (
            .O(N__27842),
            .I(N__27836));
    LocalMux I__3874 (
            .O(N__27839),
            .I(n3108));
    LocalMux I__3873 (
            .O(N__27836),
            .I(n3108));
    InMux I__3872 (
            .O(N__27831),
            .I(N__27828));
    LocalMux I__3871 (
            .O(N__27828),
            .I(n14174));
    CascadeMux I__3870 (
            .O(N__27825),
            .I(N__27822));
    InMux I__3869 (
            .O(N__27822),
            .I(N__27819));
    LocalMux I__3868 (
            .O(N__27819),
            .I(N__27816));
    Odrv4 I__3867 (
            .O(N__27816),
            .I(n3190));
    InMux I__3866 (
            .O(N__27813),
            .I(N__27810));
    LocalMux I__3865 (
            .O(N__27810),
            .I(N__27806));
    InMux I__3864 (
            .O(N__27809),
            .I(N__27803));
    Span4Mux_h I__3863 (
            .O(N__27806),
            .I(N__27799));
    LocalMux I__3862 (
            .O(N__27803),
            .I(N__27796));
    InMux I__3861 (
            .O(N__27802),
            .I(N__27793));
    Odrv4 I__3860 (
            .O(N__27799),
            .I(n3121));
    Odrv4 I__3859 (
            .O(N__27796),
            .I(n3121));
    LocalMux I__3858 (
            .O(N__27793),
            .I(n3121));
    InMux I__3857 (
            .O(N__27786),
            .I(N__27783));
    LocalMux I__3856 (
            .O(N__27783),
            .I(N__27780));
    Odrv12 I__3855 (
            .O(N__27780),
            .I(n3188));
    InMux I__3854 (
            .O(N__27777),
            .I(N__27774));
    LocalMux I__3853 (
            .O(N__27774),
            .I(N__27771));
    Odrv4 I__3852 (
            .O(N__27771),
            .I(n3192));
    CascadeMux I__3851 (
            .O(N__27768),
            .I(N__27765));
    InMux I__3850 (
            .O(N__27765),
            .I(N__27761));
    CascadeMux I__3849 (
            .O(N__27764),
            .I(N__27758));
    LocalMux I__3848 (
            .O(N__27761),
            .I(N__27755));
    InMux I__3847 (
            .O(N__27758),
            .I(N__27752));
    Span4Mux_h I__3846 (
            .O(N__27755),
            .I(N__27748));
    LocalMux I__3845 (
            .O(N__27752),
            .I(N__27745));
    InMux I__3844 (
            .O(N__27751),
            .I(N__27742));
    Odrv4 I__3843 (
            .O(N__27748),
            .I(n3125));
    Odrv4 I__3842 (
            .O(N__27745),
            .I(n3125));
    LocalMux I__3841 (
            .O(N__27742),
            .I(n3125));
    InMux I__3840 (
            .O(N__27735),
            .I(N__27730));
    InMux I__3839 (
            .O(N__27734),
            .I(N__27727));
    InMux I__3838 (
            .O(N__27733),
            .I(N__27724));
    LocalMux I__3837 (
            .O(N__27730),
            .I(N__27721));
    LocalMux I__3836 (
            .O(N__27727),
            .I(N__27718));
    LocalMux I__3835 (
            .O(N__27724),
            .I(N__27715));
    Span4Mux_s2_h I__3834 (
            .O(N__27721),
            .I(N__27712));
    Odrv4 I__3833 (
            .O(N__27718),
            .I(n3127));
    Odrv4 I__3832 (
            .O(N__27715),
            .I(n3127));
    Odrv4 I__3831 (
            .O(N__27712),
            .I(n3127));
    CascadeMux I__3830 (
            .O(N__27705),
            .I(N__27702));
    InMux I__3829 (
            .O(N__27702),
            .I(N__27699));
    LocalMux I__3828 (
            .O(N__27699),
            .I(N__27696));
    Span4Mux_h I__3827 (
            .O(N__27696),
            .I(N__27693));
    Odrv4 I__3826 (
            .O(N__27693),
            .I(n3194));
    CascadeMux I__3825 (
            .O(N__27690),
            .I(n3226_cascade_));
    InMux I__3824 (
            .O(N__27687),
            .I(N__27684));
    LocalMux I__3823 (
            .O(N__27684),
            .I(N__27680));
    InMux I__3822 (
            .O(N__27683),
            .I(N__27677));
    Span4Mux_h I__3821 (
            .O(N__27680),
            .I(N__27671));
    LocalMux I__3820 (
            .O(N__27677),
            .I(N__27671));
    InMux I__3819 (
            .O(N__27676),
            .I(N__27668));
    Odrv4 I__3818 (
            .O(N__27671),
            .I(n3119));
    LocalMux I__3817 (
            .O(N__27668),
            .I(n3119));
    CascadeMux I__3816 (
            .O(N__27663),
            .I(N__27660));
    InMux I__3815 (
            .O(N__27660),
            .I(N__27657));
    LocalMux I__3814 (
            .O(N__27657),
            .I(N__27654));
    Span4Mux_s2_v I__3813 (
            .O(N__27654),
            .I(N__27651));
    Odrv4 I__3812 (
            .O(N__27651),
            .I(n3186));
    CascadeMux I__3811 (
            .O(N__27648),
            .I(n3218_cascade_));
    CascadeMux I__3810 (
            .O(N__27645),
            .I(N__27642));
    InMux I__3809 (
            .O(N__27642),
            .I(N__27639));
    LocalMux I__3808 (
            .O(N__27639),
            .I(N__27636));
    Odrv4 I__3807 (
            .O(N__27636),
            .I(n3180));
    CascadeMux I__3806 (
            .O(N__27633),
            .I(N__27630));
    InMux I__3805 (
            .O(N__27630),
            .I(N__27627));
    LocalMux I__3804 (
            .O(N__27627),
            .I(n3098));
    CascadeMux I__3803 (
            .O(N__27624),
            .I(n3130_cascade_));
    InMux I__3802 (
            .O(N__27621),
            .I(N__27618));
    LocalMux I__3801 (
            .O(N__27618),
            .I(n3101));
    InMux I__3800 (
            .O(N__27615),
            .I(N__27612));
    LocalMux I__3799 (
            .O(N__27612),
            .I(n3097));
    InMux I__3798 (
            .O(N__27609),
            .I(N__27606));
    LocalMux I__3797 (
            .O(N__27606),
            .I(n3100));
    CascadeMux I__3796 (
            .O(N__27603),
            .I(n3132_cascade_));
    InMux I__3795 (
            .O(N__27600),
            .I(N__27597));
    LocalMux I__3794 (
            .O(N__27597),
            .I(n11945));
    InMux I__3793 (
            .O(N__27594),
            .I(N__27591));
    LocalMux I__3792 (
            .O(N__27591),
            .I(n3080));
    CascadeMux I__3791 (
            .O(N__27588),
            .I(N__27584));
    InMux I__3790 (
            .O(N__27587),
            .I(N__27581));
    InMux I__3789 (
            .O(N__27584),
            .I(N__27578));
    LocalMux I__3788 (
            .O(N__27581),
            .I(N__27575));
    LocalMux I__3787 (
            .O(N__27578),
            .I(N__27571));
    Span4Mux_v I__3786 (
            .O(N__27575),
            .I(N__27568));
    InMux I__3785 (
            .O(N__27574),
            .I(N__27565));
    Odrv4 I__3784 (
            .O(N__27571),
            .I(n3013));
    Odrv4 I__3783 (
            .O(N__27568),
            .I(n3013));
    LocalMux I__3782 (
            .O(N__27565),
            .I(n3013));
    CascadeMux I__3781 (
            .O(N__27558),
            .I(n23_adj_715_cascade_));
    InMux I__3780 (
            .O(N__27555),
            .I(N__27552));
    LocalMux I__3779 (
            .O(N__27552),
            .I(N__27548));
    CascadeMux I__3778 (
            .O(N__27551),
            .I(N__27545));
    Span4Mux_h I__3777 (
            .O(N__27548),
            .I(N__27541));
    InMux I__3776 (
            .O(N__27545),
            .I(N__27538));
    InMux I__3775 (
            .O(N__27544),
            .I(N__27535));
    Odrv4 I__3774 (
            .O(N__27541),
            .I(n3123));
    LocalMux I__3773 (
            .O(N__27538),
            .I(n3123));
    LocalMux I__3772 (
            .O(N__27535),
            .I(n3123));
    CascadeMux I__3771 (
            .O(N__27528),
            .I(N__27525));
    InMux I__3770 (
            .O(N__27525),
            .I(N__27522));
    LocalMux I__3769 (
            .O(N__27522),
            .I(N__27519));
    Span4Mux_h I__3768 (
            .O(N__27519),
            .I(N__27516));
    Odrv4 I__3767 (
            .O(N__27516),
            .I(n2995));
    CascadeMux I__3766 (
            .O(N__27513),
            .I(N__27510));
    InMux I__3765 (
            .O(N__27510),
            .I(N__27507));
    LocalMux I__3764 (
            .O(N__27507),
            .I(N__27504));
    Span4Mux_v I__3763 (
            .O(N__27504),
            .I(N__27501));
    Odrv4 I__3762 (
            .O(N__27501),
            .I(n3000));
    InMux I__3761 (
            .O(N__27498),
            .I(N__27495));
    LocalMux I__3760 (
            .O(N__27495),
            .I(N__27491));
    InMux I__3759 (
            .O(N__27494),
            .I(N__27488));
    Span4Mux_s2_v I__3758 (
            .O(N__27491),
            .I(N__27482));
    LocalMux I__3757 (
            .O(N__27488),
            .I(N__27482));
    InMux I__3756 (
            .O(N__27487),
            .I(N__27479));
    Odrv4 I__3755 (
            .O(N__27482),
            .I(n3015));
    LocalMux I__3754 (
            .O(N__27479),
            .I(n3015));
    InMux I__3753 (
            .O(N__27474),
            .I(N__27471));
    LocalMux I__3752 (
            .O(N__27471),
            .I(N__27468));
    Span4Mux_v I__3751 (
            .O(N__27468),
            .I(N__27465));
    Odrv4 I__3750 (
            .O(N__27465),
            .I(n14736));
    InMux I__3749 (
            .O(N__27462),
            .I(N__27458));
    CascadeMux I__3748 (
            .O(N__27461),
            .I(N__27454));
    LocalMux I__3747 (
            .O(N__27458),
            .I(N__27451));
    InMux I__3746 (
            .O(N__27457),
            .I(N__27448));
    InMux I__3745 (
            .O(N__27454),
            .I(N__27445));
    Span4Mux_s3_v I__3744 (
            .O(N__27451),
            .I(N__27440));
    LocalMux I__3743 (
            .O(N__27448),
            .I(N__27440));
    LocalMux I__3742 (
            .O(N__27445),
            .I(n3014));
    Odrv4 I__3741 (
            .O(N__27440),
            .I(n3014));
    CascadeMux I__3740 (
            .O(N__27435),
            .I(n14742_cascade_));
    InMux I__3739 (
            .O(N__27432),
            .I(N__27428));
    CascadeMux I__3738 (
            .O(N__27431),
            .I(N__27425));
    LocalMux I__3737 (
            .O(N__27428),
            .I(N__27422));
    InMux I__3736 (
            .O(N__27425),
            .I(N__27419));
    Span4Mux_s2_v I__3735 (
            .O(N__27422),
            .I(N__27413));
    LocalMux I__3734 (
            .O(N__27419),
            .I(N__27413));
    InMux I__3733 (
            .O(N__27418),
            .I(N__27410));
    Odrv4 I__3732 (
            .O(N__27413),
            .I(n3011));
    LocalMux I__3731 (
            .O(N__27410),
            .I(n3011));
    InMux I__3730 (
            .O(N__27405),
            .I(N__27401));
    InMux I__3729 (
            .O(N__27404),
            .I(N__27398));
    LocalMux I__3728 (
            .O(N__27401),
            .I(N__27395));
    LocalMux I__3727 (
            .O(N__27398),
            .I(N__27391));
    Span4Mux_h I__3726 (
            .O(N__27395),
            .I(N__27388));
    InMux I__3725 (
            .O(N__27394),
            .I(N__27385));
    Span4Mux_h I__3724 (
            .O(N__27391),
            .I(N__27382));
    Span4Mux_v I__3723 (
            .O(N__27388),
            .I(N__27377));
    LocalMux I__3722 (
            .O(N__27385),
            .I(N__27377));
    Odrv4 I__3721 (
            .O(N__27382),
            .I(n3009));
    Odrv4 I__3720 (
            .O(N__27377),
            .I(n3009));
    CascadeMux I__3719 (
            .O(N__27372),
            .I(n14748_cascade_));
    CascadeMux I__3718 (
            .O(N__27369),
            .I(N__27366));
    InMux I__3717 (
            .O(N__27366),
            .I(N__27362));
    InMux I__3716 (
            .O(N__27365),
            .I(N__27359));
    LocalMux I__3715 (
            .O(N__27362),
            .I(N__27356));
    LocalMux I__3714 (
            .O(N__27359),
            .I(N__27353));
    Odrv4 I__3713 (
            .O(N__27356),
            .I(n3006));
    Odrv4 I__3712 (
            .O(N__27353),
            .I(n3006));
    InMux I__3711 (
            .O(N__27348),
            .I(N__27342));
    InMux I__3710 (
            .O(N__27347),
            .I(N__27342));
    LocalMux I__3709 (
            .O(N__27342),
            .I(N__27338));
    InMux I__3708 (
            .O(N__27341),
            .I(N__27335));
    Sp12to4 I__3707 (
            .O(N__27338),
            .I(N__27330));
    LocalMux I__3706 (
            .O(N__27335),
            .I(N__27330));
    Odrv12 I__3705 (
            .O(N__27330),
            .I(n3008));
    CascadeMux I__3704 (
            .O(N__27327),
            .I(n14754_cascade_));
    InMux I__3703 (
            .O(N__27324),
            .I(N__27318));
    InMux I__3702 (
            .O(N__27323),
            .I(N__27318));
    LocalMux I__3701 (
            .O(N__27318),
            .I(N__27315));
    Span4Mux_s2_v I__3700 (
            .O(N__27315),
            .I(N__27312));
    IoSpan4Mux I__3699 (
            .O(N__27312),
            .I(N__27308));
    InMux I__3698 (
            .O(N__27311),
            .I(N__27305));
    IoSpan4Mux I__3697 (
            .O(N__27308),
            .I(N__27302));
    LocalMux I__3696 (
            .O(N__27305),
            .I(N__27299));
    Span4Mux_s0_h I__3695 (
            .O(N__27302),
            .I(N__27294));
    Span4Mux_v I__3694 (
            .O(N__27299),
            .I(N__27294));
    Odrv4 I__3693 (
            .O(N__27294),
            .I(n3007));
    InMux I__3692 (
            .O(N__27291),
            .I(N__27288));
    LocalMux I__3691 (
            .O(N__27288),
            .I(n3099));
    CascadeMux I__3690 (
            .O(N__27285),
            .I(n3039_cascade_));
    InMux I__3689 (
            .O(N__27282),
            .I(N__27279));
    LocalMux I__3688 (
            .O(N__27279),
            .I(N__27274));
    InMux I__3687 (
            .O(N__27278),
            .I(N__27271));
    InMux I__3686 (
            .O(N__27277),
            .I(N__27268));
    Span4Mux_h I__3685 (
            .O(N__27274),
            .I(N__27263));
    LocalMux I__3684 (
            .O(N__27271),
            .I(N__27263));
    LocalMux I__3683 (
            .O(N__27268),
            .I(N__27260));
    Span4Mux_v I__3682 (
            .O(N__27263),
            .I(N__27257));
    Odrv4 I__3681 (
            .O(N__27260),
            .I(n3018));
    Odrv4 I__3680 (
            .O(N__27257),
            .I(n3018));
    CascadeMux I__3679 (
            .O(N__27252),
            .I(N__27249));
    InMux I__3678 (
            .O(N__27249),
            .I(N__27246));
    LocalMux I__3677 (
            .O(N__27246),
            .I(n3085));
    InMux I__3676 (
            .O(N__27243),
            .I(N__27240));
    LocalMux I__3675 (
            .O(N__27240),
            .I(N__27236));
    InMux I__3674 (
            .O(N__27239),
            .I(N__27232));
    Span4Mux_h I__3673 (
            .O(N__27236),
            .I(N__27229));
    InMux I__3672 (
            .O(N__27235),
            .I(N__27226));
    LocalMux I__3671 (
            .O(N__27232),
            .I(N__27223));
    Odrv4 I__3670 (
            .O(N__27229),
            .I(n2817));
    LocalMux I__3669 (
            .O(N__27226),
            .I(n2817));
    Odrv4 I__3668 (
            .O(N__27223),
            .I(n2817));
    InMux I__3667 (
            .O(N__27216),
            .I(N__27213));
    LocalMux I__3666 (
            .O(N__27213),
            .I(N__27210));
    Span4Mux_h I__3665 (
            .O(N__27210),
            .I(N__27207));
    Odrv4 I__3664 (
            .O(N__27207),
            .I(n2884));
    InMux I__3663 (
            .O(N__27204),
            .I(N__27201));
    LocalMux I__3662 (
            .O(N__27201),
            .I(N__27197));
    InMux I__3661 (
            .O(N__27200),
            .I(N__27193));
    Span4Mux_s3_h I__3660 (
            .O(N__27197),
            .I(N__27190));
    InMux I__3659 (
            .O(N__27196),
            .I(N__27187));
    LocalMux I__3658 (
            .O(N__27193),
            .I(n2916));
    Odrv4 I__3657 (
            .O(N__27190),
            .I(n2916));
    LocalMux I__3656 (
            .O(N__27187),
            .I(n2916));
    CascadeMux I__3655 (
            .O(N__27180),
            .I(N__27177));
    InMux I__3654 (
            .O(N__27177),
            .I(N__27174));
    LocalMux I__3653 (
            .O(N__27174),
            .I(N__27171));
    Odrv4 I__3652 (
            .O(N__27171),
            .I(n2981));
    CascadeMux I__3651 (
            .O(N__27168),
            .I(N__27163));
    CascadeMux I__3650 (
            .O(N__27167),
            .I(N__27160));
    CascadeMux I__3649 (
            .O(N__27166),
            .I(N__27157));
    InMux I__3648 (
            .O(N__27163),
            .I(N__27154));
    InMux I__3647 (
            .O(N__27160),
            .I(N__27151));
    InMux I__3646 (
            .O(N__27157),
            .I(N__27148));
    LocalMux I__3645 (
            .O(N__27154),
            .I(N__27145));
    LocalMux I__3644 (
            .O(N__27151),
            .I(N__27142));
    LocalMux I__3643 (
            .O(N__27148),
            .I(N__27139));
    Span4Mux_v I__3642 (
            .O(N__27145),
            .I(N__27134));
    Span4Mux_s3_h I__3641 (
            .O(N__27142),
            .I(N__27134));
    Odrv12 I__3640 (
            .O(N__27139),
            .I(n2929));
    Odrv4 I__3639 (
            .O(N__27134),
            .I(n2929));
    InMux I__3638 (
            .O(N__27129),
            .I(N__27126));
    LocalMux I__3637 (
            .O(N__27126),
            .I(n14222));
    InMux I__3636 (
            .O(N__27123),
            .I(N__27120));
    LocalMux I__3635 (
            .O(N__27120),
            .I(N__27115));
    InMux I__3634 (
            .O(N__27119),
            .I(N__27112));
    InMux I__3633 (
            .O(N__27118),
            .I(N__27109));
    Span4Mux_v I__3632 (
            .O(N__27115),
            .I(N__27106));
    LocalMux I__3631 (
            .O(N__27112),
            .I(N__27103));
    LocalMux I__3630 (
            .O(N__27109),
            .I(n2915));
    Odrv4 I__3629 (
            .O(N__27106),
            .I(n2915));
    Odrv4 I__3628 (
            .O(N__27103),
            .I(n2915));
    CascadeMux I__3627 (
            .O(N__27096),
            .I(n14224_cascade_));
    InMux I__3626 (
            .O(N__27093),
            .I(N__27088));
    InMux I__3625 (
            .O(N__27092),
            .I(N__27083));
    InMux I__3624 (
            .O(N__27091),
            .I(N__27083));
    LocalMux I__3623 (
            .O(N__27088),
            .I(N__27078));
    LocalMux I__3622 (
            .O(N__27083),
            .I(N__27078));
    Span4Mux_h I__3621 (
            .O(N__27078),
            .I(N__27075));
    Odrv4 I__3620 (
            .O(N__27075),
            .I(n2914));
    InMux I__3619 (
            .O(N__27072),
            .I(N__27068));
    InMux I__3618 (
            .O(N__27071),
            .I(N__27065));
    LocalMux I__3617 (
            .O(N__27068),
            .I(N__27059));
    LocalMux I__3616 (
            .O(N__27065),
            .I(N__27059));
    InMux I__3615 (
            .O(N__27064),
            .I(N__27056));
    Span12Mux_s3_h I__3614 (
            .O(N__27059),
            .I(N__27053));
    LocalMux I__3613 (
            .O(N__27056),
            .I(N__27050));
    Odrv12 I__3612 (
            .O(N__27053),
            .I(n2910));
    Odrv4 I__3611 (
            .O(N__27050),
            .I(n2910));
    CascadeMux I__3610 (
            .O(N__27045),
            .I(n14230_cascade_));
    InMux I__3609 (
            .O(N__27042),
            .I(N__27038));
    InMux I__3608 (
            .O(N__27041),
            .I(N__27035));
    LocalMux I__3607 (
            .O(N__27038),
            .I(n2912));
    LocalMux I__3606 (
            .O(N__27035),
            .I(n2912));
    CascadeMux I__3605 (
            .O(N__27030),
            .I(N__27027));
    InMux I__3604 (
            .O(N__27027),
            .I(N__27023));
    InMux I__3603 (
            .O(N__27026),
            .I(N__27020));
    LocalMux I__3602 (
            .O(N__27023),
            .I(N__27017));
    LocalMux I__3601 (
            .O(N__27020),
            .I(N__27014));
    Span4Mux_h I__3600 (
            .O(N__27017),
            .I(N__27011));
    Span4Mux_h I__3599 (
            .O(N__27014),
            .I(N__27008));
    Odrv4 I__3598 (
            .O(N__27011),
            .I(n2908));
    Odrv4 I__3597 (
            .O(N__27008),
            .I(n2908));
    InMux I__3596 (
            .O(N__27003),
            .I(N__26999));
    InMux I__3595 (
            .O(N__27002),
            .I(N__26996));
    LocalMux I__3594 (
            .O(N__26999),
            .I(N__26993));
    LocalMux I__3593 (
            .O(N__26996),
            .I(N__26990));
    Span4Mux_v I__3592 (
            .O(N__26993),
            .I(N__26987));
    Odrv4 I__3591 (
            .O(N__26990),
            .I(n2907));
    Odrv4 I__3590 (
            .O(N__26987),
            .I(n2907));
    CascadeMux I__3589 (
            .O(N__26982),
            .I(n14236_cascade_));
    CascadeMux I__3588 (
            .O(N__26979),
            .I(N__26976));
    InMux I__3587 (
            .O(N__26976),
            .I(N__26973));
    LocalMux I__3586 (
            .O(N__26973),
            .I(N__26968));
    InMux I__3585 (
            .O(N__26972),
            .I(N__26965));
    InMux I__3584 (
            .O(N__26971),
            .I(N__26962));
    Span4Mux_s3_h I__3583 (
            .O(N__26968),
            .I(N__26957));
    LocalMux I__3582 (
            .O(N__26965),
            .I(N__26957));
    LocalMux I__3581 (
            .O(N__26962),
            .I(n2909));
    Odrv4 I__3580 (
            .O(N__26957),
            .I(n2909));
    CascadeMux I__3579 (
            .O(N__26952),
            .I(n2940_cascade_));
    InMux I__3578 (
            .O(N__26949),
            .I(N__26946));
    LocalMux I__3577 (
            .O(N__26946),
            .I(N__26943));
    Span4Mux_h I__3576 (
            .O(N__26943),
            .I(N__26940));
    Odrv4 I__3575 (
            .O(N__26940),
            .I(n2997));
    InMux I__3574 (
            .O(N__26937),
            .I(N__26932));
    InMux I__3573 (
            .O(N__26936),
            .I(N__26927));
    InMux I__3572 (
            .O(N__26935),
            .I(N__26927));
    LocalMux I__3571 (
            .O(N__26932),
            .I(n2911));
    LocalMux I__3570 (
            .O(N__26927),
            .I(n2911));
    InMux I__3569 (
            .O(N__26922),
            .I(N__26919));
    LocalMux I__3568 (
            .O(N__26919),
            .I(N__26916));
    Odrv4 I__3567 (
            .O(N__26916),
            .I(n2978));
    InMux I__3566 (
            .O(N__26913),
            .I(N__26910));
    LocalMux I__3565 (
            .O(N__26910),
            .I(N__26907));
    Span4Mux_v I__3564 (
            .O(N__26907),
            .I(N__26904));
    Odrv4 I__3563 (
            .O(N__26904),
            .I(n3081));
    InMux I__3562 (
            .O(N__26901),
            .I(N__26898));
    LocalMux I__3561 (
            .O(N__26898),
            .I(N__26895));
    Span4Mux_s2_h I__3560 (
            .O(N__26895),
            .I(N__26890));
    InMux I__3559 (
            .O(N__26894),
            .I(N__26885));
    InMux I__3558 (
            .O(N__26893),
            .I(N__26885));
    Odrv4 I__3557 (
            .O(N__26890),
            .I(n2810));
    LocalMux I__3556 (
            .O(N__26885),
            .I(n2810));
    InMux I__3555 (
            .O(N__26880),
            .I(N__26877));
    LocalMux I__3554 (
            .O(N__26877),
            .I(N__26874));
    Odrv12 I__3553 (
            .O(N__26874),
            .I(n2877));
    CascadeMux I__3552 (
            .O(N__26871),
            .I(N__26868));
    InMux I__3551 (
            .O(N__26868),
            .I(N__26865));
    LocalMux I__3550 (
            .O(N__26865),
            .I(N__26862));
    Span4Mux_v I__3549 (
            .O(N__26862),
            .I(N__26859));
    Odrv4 I__3548 (
            .O(N__26859),
            .I(n2976));
    InMux I__3547 (
            .O(N__26856),
            .I(N__26853));
    LocalMux I__3546 (
            .O(N__26853),
            .I(N__26850));
    Span4Mux_h I__3545 (
            .O(N__26850),
            .I(N__26847));
    Odrv4 I__3544 (
            .O(N__26847),
            .I(n2886));
    InMux I__3543 (
            .O(N__26844),
            .I(N__26840));
    CascadeMux I__3542 (
            .O(N__26843),
            .I(N__26837));
    LocalMux I__3541 (
            .O(N__26840),
            .I(N__26834));
    InMux I__3540 (
            .O(N__26837),
            .I(N__26830));
    Span4Mux_s2_h I__3539 (
            .O(N__26834),
            .I(N__26827));
    InMux I__3538 (
            .O(N__26833),
            .I(N__26824));
    LocalMux I__3537 (
            .O(N__26830),
            .I(n2819));
    Odrv4 I__3536 (
            .O(N__26827),
            .I(n2819));
    LocalMux I__3535 (
            .O(N__26824),
            .I(n2819));
    InMux I__3534 (
            .O(N__26817),
            .I(N__26814));
    LocalMux I__3533 (
            .O(N__26814),
            .I(N__26810));
    InMux I__3532 (
            .O(N__26813),
            .I(N__26807));
    IoSpan4Mux I__3531 (
            .O(N__26810),
            .I(N__26802));
    LocalMux I__3530 (
            .O(N__26807),
            .I(N__26802));
    Span4Mux_s3_h I__3529 (
            .O(N__26802),
            .I(N__26799));
    Odrv4 I__3528 (
            .O(N__26799),
            .I(n2918));
    InMux I__3527 (
            .O(N__26796),
            .I(N__26792));
    InMux I__3526 (
            .O(N__26795),
            .I(N__26789));
    LocalMux I__3525 (
            .O(N__26792),
            .I(N__26786));
    LocalMux I__3524 (
            .O(N__26789),
            .I(n2927));
    Odrv4 I__3523 (
            .O(N__26786),
            .I(n2927));
    InMux I__3522 (
            .O(N__26781),
            .I(N__26778));
    LocalMux I__3521 (
            .O(N__26778),
            .I(N__26775));
    Span4Mux_s2_h I__3520 (
            .O(N__26775),
            .I(N__26770));
    InMux I__3519 (
            .O(N__26774),
            .I(N__26767));
    InMux I__3518 (
            .O(N__26773),
            .I(N__26764));
    Odrv4 I__3517 (
            .O(N__26770),
            .I(n2926));
    LocalMux I__3516 (
            .O(N__26767),
            .I(n2926));
    LocalMux I__3515 (
            .O(N__26764),
            .I(n2926));
    CascadeMux I__3514 (
            .O(N__26757),
            .I(n2918_cascade_));
    InMux I__3513 (
            .O(N__26754),
            .I(N__26751));
    LocalMux I__3512 (
            .O(N__26751),
            .I(N__26747));
    CascadeMux I__3511 (
            .O(N__26750),
            .I(N__26744));
    Span4Mux_v I__3510 (
            .O(N__26747),
            .I(N__26741));
    InMux I__3509 (
            .O(N__26744),
            .I(N__26737));
    IoSpan4Mux I__3508 (
            .O(N__26741),
            .I(N__26734));
    InMux I__3507 (
            .O(N__26740),
            .I(N__26731));
    LocalMux I__3506 (
            .O(N__26737),
            .I(N__26728));
    Span4Mux_s1_h I__3505 (
            .O(N__26734),
            .I(N__26723));
    LocalMux I__3504 (
            .O(N__26731),
            .I(N__26723));
    Span4Mux_v I__3503 (
            .O(N__26728),
            .I(N__26720));
    Odrv4 I__3502 (
            .O(N__26723),
            .I(n2825));
    Odrv4 I__3501 (
            .O(N__26720),
            .I(n2825));
    CascadeMux I__3500 (
            .O(N__26715),
            .I(N__26712));
    InMux I__3499 (
            .O(N__26712),
            .I(N__26709));
    LocalMux I__3498 (
            .O(N__26709),
            .I(N__26706));
    Span4Mux_v I__3497 (
            .O(N__26706),
            .I(N__26703));
    Odrv4 I__3496 (
            .O(N__26703),
            .I(n2892));
    InMux I__3495 (
            .O(N__26700),
            .I(N__26695));
    InMux I__3494 (
            .O(N__26699),
            .I(N__26692));
    InMux I__3493 (
            .O(N__26698),
            .I(N__26689));
    LocalMux I__3492 (
            .O(N__26695),
            .I(n2921));
    LocalMux I__3491 (
            .O(N__26692),
            .I(n2921));
    LocalMux I__3490 (
            .O(N__26689),
            .I(n2921));
    InMux I__3489 (
            .O(N__26682),
            .I(N__26679));
    LocalMux I__3488 (
            .O(N__26679),
            .I(N__26676));
    Span4Mux_s2_h I__3487 (
            .O(N__26676),
            .I(N__26671));
    InMux I__3486 (
            .O(N__26675),
            .I(N__26668));
    InMux I__3485 (
            .O(N__26674),
            .I(N__26665));
    Odrv4 I__3484 (
            .O(N__26671),
            .I(n2922));
    LocalMux I__3483 (
            .O(N__26668),
            .I(n2922));
    LocalMux I__3482 (
            .O(N__26665),
            .I(n2922));
    CascadeMux I__3481 (
            .O(N__26658),
            .I(n2924_cascade_));
    InMux I__3480 (
            .O(N__26655),
            .I(N__26650));
    InMux I__3479 (
            .O(N__26654),
            .I(N__26647));
    InMux I__3478 (
            .O(N__26653),
            .I(N__26644));
    LocalMux I__3477 (
            .O(N__26650),
            .I(n2919));
    LocalMux I__3476 (
            .O(N__26647),
            .I(n2919));
    LocalMux I__3475 (
            .O(N__26644),
            .I(n2919));
    CascadeMux I__3474 (
            .O(N__26637),
            .I(n14212_cascade_));
    InMux I__3473 (
            .O(N__26634),
            .I(N__26631));
    LocalMux I__3472 (
            .O(N__26631),
            .I(n14216));
    CascadeMux I__3471 (
            .O(N__26628),
            .I(N__26625));
    InMux I__3470 (
            .O(N__26625),
            .I(N__26622));
    LocalMux I__3469 (
            .O(N__26622),
            .I(N__26619));
    Span4Mux_v I__3468 (
            .O(N__26619),
            .I(N__26615));
    InMux I__3467 (
            .O(N__26618),
            .I(N__26611));
    Span4Mux_s2_h I__3466 (
            .O(N__26615),
            .I(N__26608));
    InMux I__3465 (
            .O(N__26614),
            .I(N__26605));
    LocalMux I__3464 (
            .O(N__26611),
            .I(n2733));
    Odrv4 I__3463 (
            .O(N__26608),
            .I(n2733));
    LocalMux I__3462 (
            .O(N__26605),
            .I(n2733));
    CascadeMux I__3461 (
            .O(N__26598),
            .I(N__26595));
    InMux I__3460 (
            .O(N__26595),
            .I(N__26592));
    LocalMux I__3459 (
            .O(N__26592),
            .I(N__26589));
    Span4Mux_v I__3458 (
            .O(N__26589),
            .I(N__26586));
    Span4Mux_v I__3457 (
            .O(N__26586),
            .I(N__26583));
    Odrv4 I__3456 (
            .O(N__26583),
            .I(n2800));
    CascadeMux I__3455 (
            .O(N__26580),
            .I(n2832_cascade_));
    CascadeMux I__3454 (
            .O(N__26577),
            .I(N__26574));
    InMux I__3453 (
            .O(N__26574),
            .I(N__26569));
    InMux I__3452 (
            .O(N__26573),
            .I(N__26566));
    InMux I__3451 (
            .O(N__26572),
            .I(N__26563));
    LocalMux I__3450 (
            .O(N__26569),
            .I(N__26560));
    LocalMux I__3449 (
            .O(N__26566),
            .I(N__26557));
    LocalMux I__3448 (
            .O(N__26563),
            .I(N__26552));
    Span4Mux_s1_h I__3447 (
            .O(N__26560),
            .I(N__26552));
    Span4Mux_v I__3446 (
            .O(N__26557),
            .I(N__26549));
    Odrv4 I__3445 (
            .O(N__26552),
            .I(n2833));
    Odrv4 I__3444 (
            .O(N__26549),
            .I(n2833));
    CascadeMux I__3443 (
            .O(N__26544),
            .I(N__26541));
    InMux I__3442 (
            .O(N__26541),
            .I(N__26537));
    CascadeMux I__3441 (
            .O(N__26540),
            .I(N__26534));
    LocalMux I__3440 (
            .O(N__26537),
            .I(N__26530));
    InMux I__3439 (
            .O(N__26534),
            .I(N__26525));
    InMux I__3438 (
            .O(N__26533),
            .I(N__26525));
    Span4Mux_s2_h I__3437 (
            .O(N__26530),
            .I(N__26522));
    LocalMux I__3436 (
            .O(N__26525),
            .I(n2830));
    Odrv4 I__3435 (
            .O(N__26522),
            .I(n2830));
    CascadeMux I__3434 (
            .O(N__26517),
            .I(n11953_cascade_));
    InMux I__3433 (
            .O(N__26514),
            .I(N__26511));
    LocalMux I__3432 (
            .O(N__26511),
            .I(n13857));
    CascadeMux I__3431 (
            .O(N__26508),
            .I(N__26505));
    InMux I__3430 (
            .O(N__26505),
            .I(N__26501));
    CascadeMux I__3429 (
            .O(N__26504),
            .I(N__26497));
    LocalMux I__3428 (
            .O(N__26501),
            .I(N__26494));
    InMux I__3427 (
            .O(N__26500),
            .I(N__26491));
    InMux I__3426 (
            .O(N__26497),
            .I(N__26488));
    Span4Mux_h I__3425 (
            .O(N__26494),
            .I(N__26485));
    LocalMux I__3424 (
            .O(N__26491),
            .I(n2815));
    LocalMux I__3423 (
            .O(N__26488),
            .I(n2815));
    Odrv4 I__3422 (
            .O(N__26485),
            .I(n2815));
    InMux I__3421 (
            .O(N__26478),
            .I(N__26475));
    LocalMux I__3420 (
            .O(N__26475),
            .I(n14702));
    InMux I__3419 (
            .O(N__26472),
            .I(N__26468));
    InMux I__3418 (
            .O(N__26471),
            .I(N__26465));
    LocalMux I__3417 (
            .O(N__26468),
            .I(N__26461));
    LocalMux I__3416 (
            .O(N__26465),
            .I(N__26458));
    InMux I__3415 (
            .O(N__26464),
            .I(N__26455));
    Odrv4 I__3414 (
            .O(N__26461),
            .I(n2812));
    Odrv4 I__3413 (
            .O(N__26458),
            .I(n2812));
    LocalMux I__3412 (
            .O(N__26455),
            .I(n2812));
    CascadeMux I__3411 (
            .O(N__26448),
            .I(N__26444));
    InMux I__3410 (
            .O(N__26447),
            .I(N__26441));
    InMux I__3409 (
            .O(N__26444),
            .I(N__26438));
    LocalMux I__3408 (
            .O(N__26441),
            .I(N__26435));
    LocalMux I__3407 (
            .O(N__26438),
            .I(N__26429));
    Span4Mux_s2_h I__3406 (
            .O(N__26435),
            .I(N__26429));
    InMux I__3405 (
            .O(N__26434),
            .I(N__26426));
    Odrv4 I__3404 (
            .O(N__26429),
            .I(n2813));
    LocalMux I__3403 (
            .O(N__26426),
            .I(n2813));
    CascadeMux I__3402 (
            .O(N__26421),
            .I(n14708_cascade_));
    InMux I__3401 (
            .O(N__26418),
            .I(N__26415));
    LocalMux I__3400 (
            .O(N__26415),
            .I(N__26411));
    InMux I__3399 (
            .O(N__26414),
            .I(N__26408));
    Odrv4 I__3398 (
            .O(N__26411),
            .I(n2811));
    LocalMux I__3397 (
            .O(N__26408),
            .I(n2811));
    InMux I__3396 (
            .O(N__26403),
            .I(N__26399));
    InMux I__3395 (
            .O(N__26402),
            .I(N__26396));
    LocalMux I__3394 (
            .O(N__26399),
            .I(N__26392));
    LocalMux I__3393 (
            .O(N__26396),
            .I(N__26389));
    InMux I__3392 (
            .O(N__26395),
            .I(N__26386));
    Span4Mux_v I__3391 (
            .O(N__26392),
            .I(N__26383));
    Span4Mux_s2_h I__3390 (
            .O(N__26389),
            .I(N__26380));
    LocalMux I__3389 (
            .O(N__26386),
            .I(N__26377));
    Odrv4 I__3388 (
            .O(N__26383),
            .I(n2809));
    Odrv4 I__3387 (
            .O(N__26380),
            .I(n2809));
    Odrv4 I__3386 (
            .O(N__26377),
            .I(n2809));
    CascadeMux I__3385 (
            .O(N__26370),
            .I(n14714_cascade_));
    CascadeMux I__3384 (
            .O(N__26367),
            .I(N__26363));
    InMux I__3383 (
            .O(N__26366),
            .I(N__26360));
    InMux I__3382 (
            .O(N__26363),
            .I(N__26357));
    LocalMux I__3381 (
            .O(N__26360),
            .I(N__26354));
    LocalMux I__3380 (
            .O(N__26357),
            .I(N__26351));
    Span4Mux_v I__3379 (
            .O(N__26354),
            .I(N__26348));
    Span4Mux_v I__3378 (
            .O(N__26351),
            .I(N__26345));
    Span4Mux_v I__3377 (
            .O(N__26348),
            .I(N__26342));
    Odrv4 I__3376 (
            .O(N__26345),
            .I(n2808));
    Odrv4 I__3375 (
            .O(N__26342),
            .I(n2808));
    InMux I__3374 (
            .O(N__26337),
            .I(N__26334));
    LocalMux I__3373 (
            .O(N__26334),
            .I(N__26329));
    InMux I__3372 (
            .O(N__26333),
            .I(N__26324));
    InMux I__3371 (
            .O(N__26332),
            .I(N__26324));
    Odrv4 I__3370 (
            .O(N__26329),
            .I(n2816));
    LocalMux I__3369 (
            .O(N__26324),
            .I(n2816));
    CascadeMux I__3368 (
            .O(N__26319),
            .I(n2841_cascade_));
    InMux I__3367 (
            .O(N__26316),
            .I(N__26313));
    LocalMux I__3366 (
            .O(N__26313),
            .I(N__26310));
    Span4Mux_h I__3365 (
            .O(N__26310),
            .I(N__26307));
    Odrv4 I__3364 (
            .O(N__26307),
            .I(n2883));
    InMux I__3363 (
            .O(N__26304),
            .I(N__26301));
    LocalMux I__3362 (
            .O(N__26301),
            .I(N__26298));
    Span4Mux_h I__3361 (
            .O(N__26298),
            .I(N__26295));
    Odrv4 I__3360 (
            .O(N__26295),
            .I(n2885));
    InMux I__3359 (
            .O(N__26292),
            .I(N__26288));
    CascadeMux I__3358 (
            .O(N__26291),
            .I(N__26285));
    LocalMux I__3357 (
            .O(N__26288),
            .I(N__26282));
    InMux I__3356 (
            .O(N__26285),
            .I(N__26278));
    Span4Mux_s1_h I__3355 (
            .O(N__26282),
            .I(N__26275));
    InMux I__3354 (
            .O(N__26281),
            .I(N__26272));
    LocalMux I__3353 (
            .O(N__26278),
            .I(n2818));
    Odrv4 I__3352 (
            .O(N__26275),
            .I(n2818));
    LocalMux I__3351 (
            .O(N__26272),
            .I(n2818));
    InMux I__3350 (
            .O(N__26265),
            .I(N__26262));
    LocalMux I__3349 (
            .O(N__26262),
            .I(N__26258));
    InMux I__3348 (
            .O(N__26261),
            .I(N__26255));
    Span12Mux_s3_h I__3347 (
            .O(N__26258),
            .I(N__26252));
    LocalMux I__3346 (
            .O(N__26255),
            .I(n2633));
    Odrv12 I__3345 (
            .O(N__26252),
            .I(n2633));
    CascadeMux I__3344 (
            .O(N__26247),
            .I(n2633_cascade_));
    CascadeMux I__3343 (
            .O(N__26244),
            .I(N__26241));
    InMux I__3342 (
            .O(N__26241),
            .I(N__26238));
    LocalMux I__3341 (
            .O(N__26238),
            .I(n12059));
    InMux I__3340 (
            .O(N__26235),
            .I(N__26232));
    LocalMux I__3339 (
            .O(N__26232),
            .I(N__26227));
    CascadeMux I__3338 (
            .O(N__26231),
            .I(N__26224));
    InMux I__3337 (
            .O(N__26230),
            .I(N__26221));
    Span12Mux_s3_h I__3336 (
            .O(N__26227),
            .I(N__26218));
    InMux I__3335 (
            .O(N__26224),
            .I(N__26215));
    LocalMux I__3334 (
            .O(N__26221),
            .I(n2618));
    Odrv12 I__3333 (
            .O(N__26218),
            .I(n2618));
    LocalMux I__3332 (
            .O(N__26215),
            .I(n2618));
    InMux I__3331 (
            .O(N__26208),
            .I(N__26204));
    InMux I__3330 (
            .O(N__26207),
            .I(N__26201));
    LocalMux I__3329 (
            .O(N__26204),
            .I(N__26198));
    LocalMux I__3328 (
            .O(N__26201),
            .I(N__26195));
    Span4Mux_s3_h I__3327 (
            .O(N__26198),
            .I(N__26192));
    Span4Mux_s3_h I__3326 (
            .O(N__26195),
            .I(N__26188));
    Span4Mux_v I__3325 (
            .O(N__26192),
            .I(N__26185));
    InMux I__3324 (
            .O(N__26191),
            .I(N__26182));
    Odrv4 I__3323 (
            .O(N__26188),
            .I(n2614));
    Odrv4 I__3322 (
            .O(N__26185),
            .I(n2614));
    LocalMux I__3321 (
            .O(N__26182),
            .I(n2614));
    InMux I__3320 (
            .O(N__26175),
            .I(N__26172));
    LocalMux I__3319 (
            .O(N__26172),
            .I(N__26169));
    Span4Mux_s3_h I__3318 (
            .O(N__26169),
            .I(N__26165));
    InMux I__3317 (
            .O(N__26168),
            .I(N__26161));
    Sp12to4 I__3316 (
            .O(N__26165),
            .I(N__26158));
    InMux I__3315 (
            .O(N__26164),
            .I(N__26155));
    LocalMux I__3314 (
            .O(N__26161),
            .I(n2613));
    Odrv12 I__3313 (
            .O(N__26158),
            .I(n2613));
    LocalMux I__3312 (
            .O(N__26155),
            .I(n2613));
    CascadeMux I__3311 (
            .O(N__26148),
            .I(N__26145));
    InMux I__3310 (
            .O(N__26145),
            .I(N__26142));
    LocalMux I__3309 (
            .O(N__26142),
            .I(N__26139));
    Span4Mux_s3_h I__3308 (
            .O(N__26139),
            .I(N__26136));
    Span4Mux_v I__3307 (
            .O(N__26136),
            .I(N__26131));
    InMux I__3306 (
            .O(N__26135),
            .I(N__26126));
    InMux I__3305 (
            .O(N__26134),
            .I(N__26126));
    Span4Mux_v I__3304 (
            .O(N__26131),
            .I(N__26123));
    LocalMux I__3303 (
            .O(N__26126),
            .I(n2619));
    Odrv4 I__3302 (
            .O(N__26123),
            .I(n2619));
    InMux I__3301 (
            .O(N__26118),
            .I(N__26115));
    LocalMux I__3300 (
            .O(N__26115),
            .I(N__26112));
    Span4Mux_h I__3299 (
            .O(N__26112),
            .I(N__26109));
    Odrv4 I__3298 (
            .O(N__26109),
            .I(n2897));
    InMux I__3297 (
            .O(N__26106),
            .I(N__26103));
    LocalMux I__3296 (
            .O(N__26103),
            .I(N__26099));
    InMux I__3295 (
            .O(N__26102),
            .I(N__26095));
    Span12Mux_s2_h I__3294 (
            .O(N__26099),
            .I(N__26092));
    InMux I__3293 (
            .O(N__26098),
            .I(N__26089));
    LocalMux I__3292 (
            .O(N__26095),
            .I(n2712));
    Odrv12 I__3291 (
            .O(N__26092),
            .I(n2712));
    LocalMux I__3290 (
            .O(N__26089),
            .I(n2712));
    CascadeMux I__3289 (
            .O(N__26082),
            .I(N__26079));
    InMux I__3288 (
            .O(N__26079),
            .I(N__26076));
    LocalMux I__3287 (
            .O(N__26076),
            .I(N__26073));
    Span12Mux_v I__3286 (
            .O(N__26073),
            .I(N__26070));
    Odrv12 I__3285 (
            .O(N__26070),
            .I(n2779));
    InMux I__3284 (
            .O(N__26067),
            .I(N__26064));
    LocalMux I__3283 (
            .O(N__26064),
            .I(N__26061));
    Odrv12 I__3282 (
            .O(N__26061),
            .I(n2878));
    CascadeMux I__3281 (
            .O(N__26058),
            .I(n2811_cascade_));
    CascadeMux I__3280 (
            .O(N__26055),
            .I(n2524_cascade_));
    CascadeMux I__3279 (
            .O(N__26052),
            .I(n14574_cascade_));
    CascadeMux I__3278 (
            .O(N__26049),
            .I(n2523_cascade_));
    InMux I__3277 (
            .O(N__26046),
            .I(N__26043));
    LocalMux I__3276 (
            .O(N__26043),
            .I(n14576));
    CascadeMux I__3275 (
            .O(N__26040),
            .I(n2527_cascade_));
    CascadeMux I__3274 (
            .O(N__26037),
            .I(N__26034));
    InMux I__3273 (
            .O(N__26034),
            .I(N__26030));
    CascadeMux I__3272 (
            .O(N__26033),
            .I(N__26027));
    LocalMux I__3271 (
            .O(N__26030),
            .I(N__26024));
    InMux I__3270 (
            .O(N__26027),
            .I(N__26021));
    Span4Mux_s2_h I__3269 (
            .O(N__26024),
            .I(N__26018));
    LocalMux I__3268 (
            .O(N__26021),
            .I(N__26014));
    Span4Mux_v I__3267 (
            .O(N__26018),
            .I(N__26011));
    InMux I__3266 (
            .O(N__26017),
            .I(N__26008));
    Span4Mux_s2_h I__3265 (
            .O(N__26014),
            .I(N__26003));
    Span4Mux_v I__3264 (
            .O(N__26011),
            .I(N__26003));
    LocalMux I__3263 (
            .O(N__26008),
            .I(n2626));
    Odrv4 I__3262 (
            .O(N__26003),
            .I(n2626));
    CascadeMux I__3261 (
            .O(N__25998),
            .I(N__25994));
    InMux I__3260 (
            .O(N__25997),
            .I(N__25991));
    InMux I__3259 (
            .O(N__25994),
            .I(N__25988));
    LocalMux I__3258 (
            .O(N__25991),
            .I(N__25985));
    LocalMux I__3257 (
            .O(N__25988),
            .I(N__25982));
    Span4Mux_s3_h I__3256 (
            .O(N__25985),
            .I(N__25979));
    Span4Mux_s3_h I__3255 (
            .O(N__25982),
            .I(N__25974));
    Span4Mux_v I__3254 (
            .O(N__25979),
            .I(N__25974));
    Odrv4 I__3253 (
            .O(N__25974),
            .I(n2617));
    CascadeMux I__3252 (
            .O(N__25971),
            .I(N__25968));
    InMux I__3251 (
            .O(N__25968),
            .I(N__25965));
    LocalMux I__3250 (
            .O(N__25965),
            .I(N__25960));
    CascadeMux I__3249 (
            .O(N__25964),
            .I(N__25957));
    InMux I__3248 (
            .O(N__25963),
            .I(N__25954));
    Span4Mux_s3_h I__3247 (
            .O(N__25960),
            .I(N__25951));
    InMux I__3246 (
            .O(N__25957),
            .I(N__25948));
    LocalMux I__3245 (
            .O(N__25954),
            .I(N__25945));
    Span4Mux_v I__3244 (
            .O(N__25951),
            .I(N__25942));
    LocalMux I__3243 (
            .O(N__25948),
            .I(n2625));
    Odrv4 I__3242 (
            .O(N__25945),
            .I(n2625));
    Odrv4 I__3241 (
            .O(N__25942),
            .I(n2625));
    CascadeMux I__3240 (
            .O(N__25935),
            .I(n2617_cascade_));
    InMux I__3239 (
            .O(N__25932),
            .I(N__25929));
    LocalMux I__3238 (
            .O(N__25929),
            .I(n14812));
    InMux I__3237 (
            .O(N__25926),
            .I(N__25923));
    LocalMux I__3236 (
            .O(N__25923),
            .I(N__25920));
    Odrv4 I__3235 (
            .O(N__25920),
            .I(n2382));
    InMux I__3234 (
            .O(N__25917),
            .I(N__25914));
    LocalMux I__3233 (
            .O(N__25914),
            .I(N__25911));
    Span4Mux_h I__3232 (
            .O(N__25911),
            .I(N__25908));
    Odrv4 I__3231 (
            .O(N__25908),
            .I(n2396));
    CascadeMux I__3230 (
            .O(N__25905),
            .I(N__25901));
    CascadeMux I__3229 (
            .O(N__25904),
            .I(N__25898));
    InMux I__3228 (
            .O(N__25901),
            .I(N__25895));
    InMux I__3227 (
            .O(N__25898),
            .I(N__25891));
    LocalMux I__3226 (
            .O(N__25895),
            .I(N__25888));
    InMux I__3225 (
            .O(N__25894),
            .I(N__25885));
    LocalMux I__3224 (
            .O(N__25891),
            .I(N__25882));
    Odrv4 I__3223 (
            .O(N__25888),
            .I(n2329));
    LocalMux I__3222 (
            .O(N__25885),
            .I(n2329));
    Odrv4 I__3221 (
            .O(N__25882),
            .I(n2329));
    CascadeMux I__3220 (
            .O(N__25875),
            .I(N__25871));
    InMux I__3219 (
            .O(N__25874),
            .I(N__25868));
    InMux I__3218 (
            .O(N__25871),
            .I(N__25865));
    LocalMux I__3217 (
            .O(N__25868),
            .I(N__25861));
    LocalMux I__3216 (
            .O(N__25865),
            .I(N__25858));
    InMux I__3215 (
            .O(N__25864),
            .I(N__25855));
    Odrv4 I__3214 (
            .O(N__25861),
            .I(n2328));
    Odrv4 I__3213 (
            .O(N__25858),
            .I(n2328));
    LocalMux I__3212 (
            .O(N__25855),
            .I(n2328));
    InMux I__3211 (
            .O(N__25848),
            .I(N__25845));
    LocalMux I__3210 (
            .O(N__25845),
            .I(N__25842));
    Span4Mux_h I__3209 (
            .O(N__25842),
            .I(N__25839));
    Odrv4 I__3208 (
            .O(N__25839),
            .I(n2395));
    CascadeMux I__3207 (
            .O(N__25836),
            .I(n2427_cascade_));
    CascadeMux I__3206 (
            .O(N__25833),
            .I(n14620_cascade_));
    CascadeMux I__3205 (
            .O(N__25830),
            .I(n2526_cascade_));
    InMux I__3204 (
            .O(N__25827),
            .I(N__25824));
    LocalMux I__3203 (
            .O(N__25824),
            .I(N__25821));
    Odrv4 I__3202 (
            .O(N__25821),
            .I(n14816));
    InMux I__3201 (
            .O(N__25818),
            .I(N__25815));
    LocalMux I__3200 (
            .O(N__25815),
            .I(n14392));
    CascadeMux I__3199 (
            .O(N__25812),
            .I(N__25809));
    InMux I__3198 (
            .O(N__25809),
            .I(N__25806));
    LocalMux I__3197 (
            .O(N__25806),
            .I(N__25802));
    InMux I__3196 (
            .O(N__25805),
            .I(N__25799));
    Span4Mux_v I__3195 (
            .O(N__25802),
            .I(N__25796));
    LocalMux I__3194 (
            .O(N__25799),
            .I(N__25793));
    Span4Mux_v I__3193 (
            .O(N__25796),
            .I(N__25788));
    Span4Mux_v I__3192 (
            .O(N__25793),
            .I(N__25788));
    Odrv4 I__3191 (
            .O(N__25788),
            .I(n2313));
    CascadeMux I__3190 (
            .O(N__25785),
            .I(n14398_cascade_));
    CascadeMux I__3189 (
            .O(N__25782),
            .I(N__25779));
    InMux I__3188 (
            .O(N__25779),
            .I(N__25775));
    InMux I__3187 (
            .O(N__25778),
            .I(N__25771));
    LocalMux I__3186 (
            .O(N__25775),
            .I(N__25768));
    InMux I__3185 (
            .O(N__25774),
            .I(N__25765));
    LocalMux I__3184 (
            .O(N__25771),
            .I(n2327));
    Odrv4 I__3183 (
            .O(N__25768),
            .I(n2327));
    LocalMux I__3182 (
            .O(N__25765),
            .I(n2327));
    CascadeMux I__3181 (
            .O(N__25758),
            .I(n2346_cascade_));
    InMux I__3180 (
            .O(N__25755),
            .I(N__25752));
    LocalMux I__3179 (
            .O(N__25752),
            .I(N__25749));
    Span4Mux_h I__3178 (
            .O(N__25749),
            .I(N__25746));
    Odrv4 I__3177 (
            .O(N__25746),
            .I(n2394));
    InMux I__3176 (
            .O(N__25743),
            .I(N__25740));
    LocalMux I__3175 (
            .O(N__25740),
            .I(N__25737));
    Span4Mux_v I__3174 (
            .O(N__25737),
            .I(N__25734));
    Odrv4 I__3173 (
            .O(N__25734),
            .I(n2284));
    InMux I__3172 (
            .O(N__25731),
            .I(N__25728));
    LocalMux I__3171 (
            .O(N__25728),
            .I(N__25724));
    InMux I__3170 (
            .O(N__25727),
            .I(N__25720));
    Span4Mux_h I__3169 (
            .O(N__25724),
            .I(N__25717));
    InMux I__3168 (
            .O(N__25723),
            .I(N__25714));
    LocalMux I__3167 (
            .O(N__25720),
            .I(n2316));
    Odrv4 I__3166 (
            .O(N__25717),
            .I(n2316));
    LocalMux I__3165 (
            .O(N__25714),
            .I(n2316));
    InMux I__3164 (
            .O(N__25707),
            .I(N__25704));
    LocalMux I__3163 (
            .O(N__25704),
            .I(N__25701));
    Span4Mux_v I__3162 (
            .O(N__25701),
            .I(N__25698));
    Odrv4 I__3161 (
            .O(N__25698),
            .I(n2282));
    InMux I__3160 (
            .O(N__25695),
            .I(N__25692));
    LocalMux I__3159 (
            .O(N__25692),
            .I(N__25689));
    Span4Mux_v I__3158 (
            .O(N__25689),
            .I(N__25685));
    InMux I__3157 (
            .O(N__25688),
            .I(N__25682));
    Odrv4 I__3156 (
            .O(N__25685),
            .I(n2314));
    LocalMux I__3155 (
            .O(N__25682),
            .I(n2314));
    CascadeMux I__3154 (
            .O(N__25677),
            .I(n2314_cascade_));
    InMux I__3153 (
            .O(N__25674),
            .I(N__25671));
    LocalMux I__3152 (
            .O(N__25671),
            .I(N__25668));
    Span4Mux_h I__3151 (
            .O(N__25668),
            .I(N__25665));
    Odrv4 I__3150 (
            .O(N__25665),
            .I(n2381));
    InMux I__3149 (
            .O(N__25662),
            .I(N__25659));
    LocalMux I__3148 (
            .O(N__25659),
            .I(N__25656));
    Odrv4 I__3147 (
            .O(N__25656),
            .I(n2392));
    CascadeMux I__3146 (
            .O(N__25653),
            .I(N__25649));
    CascadeMux I__3145 (
            .O(N__25652),
            .I(N__25646));
    InMux I__3144 (
            .O(N__25649),
            .I(N__25643));
    InMux I__3143 (
            .O(N__25646),
            .I(N__25640));
    LocalMux I__3142 (
            .O(N__25643),
            .I(N__25637));
    LocalMux I__3141 (
            .O(N__25640),
            .I(N__25631));
    Span4Mux_s3_h I__3140 (
            .O(N__25637),
            .I(N__25631));
    InMux I__3139 (
            .O(N__25636),
            .I(N__25628));
    Odrv4 I__3138 (
            .O(N__25631),
            .I(n2325));
    LocalMux I__3137 (
            .O(N__25628),
            .I(n2325));
    InMux I__3136 (
            .O(N__25623),
            .I(N__25619));
    InMux I__3135 (
            .O(N__25622),
            .I(N__25615));
    LocalMux I__3134 (
            .O(N__25619),
            .I(N__25612));
    InMux I__3133 (
            .O(N__25618),
            .I(N__25609));
    LocalMux I__3132 (
            .O(N__25615),
            .I(n2320));
    Odrv4 I__3131 (
            .O(N__25612),
            .I(n2320));
    LocalMux I__3130 (
            .O(N__25609),
            .I(n2320));
    InMux I__3129 (
            .O(N__25602),
            .I(N__25599));
    LocalMux I__3128 (
            .O(N__25599),
            .I(N__25596));
    Odrv12 I__3127 (
            .O(N__25596),
            .I(n2387));
    InMux I__3126 (
            .O(N__25593),
            .I(n12671));
    InMux I__3125 (
            .O(N__25590),
            .I(bfn_4_19_0_));
    InMux I__3124 (
            .O(N__25587),
            .I(n12673));
    InMux I__3123 (
            .O(N__25584),
            .I(n12674));
    InMux I__3122 (
            .O(N__25581),
            .I(n12675));
    InMux I__3121 (
            .O(N__25578),
            .I(N__25575));
    LocalMux I__3120 (
            .O(N__25575),
            .I(N__25571));
    InMux I__3119 (
            .O(N__25574),
            .I(N__25568));
    Odrv4 I__3118 (
            .O(N__25571),
            .I(n2214));
    LocalMux I__3117 (
            .O(N__25568),
            .I(n2214));
    CascadeMux I__3116 (
            .O(N__25563),
            .I(N__25560));
    InMux I__3115 (
            .O(N__25560),
            .I(N__25557));
    LocalMux I__3114 (
            .O(N__25557),
            .I(N__25554));
    Span4Mux_v I__3113 (
            .O(N__25554),
            .I(N__25551));
    Odrv4 I__3112 (
            .O(N__25551),
            .I(n2294));
    CascadeMux I__3111 (
            .O(N__25548),
            .I(N__25545));
    InMux I__3110 (
            .O(N__25545),
            .I(N__25542));
    LocalMux I__3109 (
            .O(N__25542),
            .I(n2186));
    CascadeMux I__3108 (
            .O(N__25539),
            .I(N__25536));
    InMux I__3107 (
            .O(N__25536),
            .I(N__25533));
    LocalMux I__3106 (
            .O(N__25533),
            .I(N__25530));
    Span4Mux_v I__3105 (
            .O(N__25530),
            .I(N__25526));
    InMux I__3104 (
            .O(N__25529),
            .I(N__25523));
    Odrv4 I__3103 (
            .O(N__25526),
            .I(n2218));
    LocalMux I__3102 (
            .O(N__25523),
            .I(n2218));
    InMux I__3101 (
            .O(N__25518),
            .I(N__25515));
    LocalMux I__3100 (
            .O(N__25515),
            .I(N__25512));
    Span4Mux_v I__3099 (
            .O(N__25512),
            .I(N__25509));
    Odrv4 I__3098 (
            .O(N__25509),
            .I(n2285));
    CascadeMux I__3097 (
            .O(N__25506),
            .I(n2218_cascade_));
    CascadeMux I__3096 (
            .O(N__25503),
            .I(N__25500));
    InMux I__3095 (
            .O(N__25500),
            .I(N__25497));
    LocalMux I__3094 (
            .O(N__25497),
            .I(n2188));
    InMux I__3093 (
            .O(N__25494),
            .I(N__25491));
    LocalMux I__3092 (
            .O(N__25491),
            .I(N__25487));
    InMux I__3091 (
            .O(N__25490),
            .I(N__25483));
    Span4Mux_v I__3090 (
            .O(N__25487),
            .I(N__25480));
    InMux I__3089 (
            .O(N__25486),
            .I(N__25477));
    LocalMux I__3088 (
            .O(N__25483),
            .I(n2220));
    Odrv4 I__3087 (
            .O(N__25480),
            .I(n2220));
    LocalMux I__3086 (
            .O(N__25477),
            .I(n2220));
    InMux I__3085 (
            .O(N__25470),
            .I(n12662));
    InMux I__3084 (
            .O(N__25467),
            .I(N__25464));
    LocalMux I__3083 (
            .O(N__25464),
            .I(n2194));
    InMux I__3082 (
            .O(N__25461),
            .I(n12663));
    InMux I__3081 (
            .O(N__25458),
            .I(N__25455));
    LocalMux I__3080 (
            .O(N__25455),
            .I(N__25452));
    Odrv4 I__3079 (
            .O(N__25452),
            .I(n2193));
    InMux I__3078 (
            .O(N__25449),
            .I(bfn_4_18_0_));
    InMux I__3077 (
            .O(N__25446),
            .I(n12665));
    InMux I__3076 (
            .O(N__25443),
            .I(n12666));
    InMux I__3075 (
            .O(N__25440),
            .I(N__25437));
    LocalMux I__3074 (
            .O(N__25437),
            .I(n2190));
    InMux I__3073 (
            .O(N__25434),
            .I(n12667));
    InMux I__3072 (
            .O(N__25431),
            .I(N__25428));
    LocalMux I__3071 (
            .O(N__25428),
            .I(N__25425));
    Odrv4 I__3070 (
            .O(N__25425),
            .I(n2189));
    InMux I__3069 (
            .O(N__25422),
            .I(n12668));
    InMux I__3068 (
            .O(N__25419),
            .I(n12669));
    InMux I__3067 (
            .O(N__25416),
            .I(N__25413));
    LocalMux I__3066 (
            .O(N__25413),
            .I(n2187));
    InMux I__3065 (
            .O(N__25410),
            .I(n12670));
    CascadeMux I__3064 (
            .O(N__25407),
            .I(n2129_cascade_));
    CascadeMux I__3063 (
            .O(N__25404),
            .I(N__25401));
    InMux I__3062 (
            .O(N__25401),
            .I(N__25397));
    CascadeMux I__3061 (
            .O(N__25400),
            .I(N__25394));
    LocalMux I__3060 (
            .O(N__25397),
            .I(N__25391));
    InMux I__3059 (
            .O(N__25394),
            .I(N__25388));
    Span4Mux_s3_h I__3058 (
            .O(N__25391),
            .I(N__25385));
    LocalMux I__3057 (
            .O(N__25388),
            .I(N__25382));
    Odrv4 I__3056 (
            .O(N__25385),
            .I(n2228));
    Odrv4 I__3055 (
            .O(N__25382),
            .I(n2228));
    InMux I__3054 (
            .O(N__25377),
            .I(N__25373));
    CascadeMux I__3053 (
            .O(N__25376),
            .I(N__25370));
    LocalMux I__3052 (
            .O(N__25373),
            .I(N__25366));
    InMux I__3051 (
            .O(N__25370),
            .I(N__25363));
    InMux I__3050 (
            .O(N__25369),
            .I(N__25360));
    Odrv4 I__3049 (
            .O(N__25366),
            .I(n2226));
    LocalMux I__3048 (
            .O(N__25363),
            .I(n2226));
    LocalMux I__3047 (
            .O(N__25360),
            .I(n2226));
    InMux I__3046 (
            .O(N__25353),
            .I(N__25350));
    LocalMux I__3045 (
            .O(N__25350),
            .I(N__25346));
    CascadeMux I__3044 (
            .O(N__25349),
            .I(N__25343));
    Span4Mux_v I__3043 (
            .O(N__25346),
            .I(N__25339));
    InMux I__3042 (
            .O(N__25343),
            .I(N__25336));
    InMux I__3041 (
            .O(N__25342),
            .I(N__25333));
    Odrv4 I__3040 (
            .O(N__25339),
            .I(n2225));
    LocalMux I__3039 (
            .O(N__25336),
            .I(n2225));
    LocalMux I__3038 (
            .O(N__25333),
            .I(n2225));
    CascadeMux I__3037 (
            .O(N__25326),
            .I(n2228_cascade_));
    InMux I__3036 (
            .O(N__25323),
            .I(N__25320));
    LocalMux I__3035 (
            .O(N__25320),
            .I(n14588));
    InMux I__3034 (
            .O(N__25317),
            .I(N__25314));
    LocalMux I__3033 (
            .O(N__25314),
            .I(n2201));
    InMux I__3032 (
            .O(N__25311),
            .I(bfn_4_17_0_));
    InMux I__3031 (
            .O(N__25308),
            .I(N__25305));
    LocalMux I__3030 (
            .O(N__25305),
            .I(N__25302));
    Odrv4 I__3029 (
            .O(N__25302),
            .I(n2200));
    InMux I__3028 (
            .O(N__25299),
            .I(n12657));
    InMux I__3027 (
            .O(N__25296),
            .I(N__25293));
    LocalMux I__3026 (
            .O(N__25293),
            .I(N__25290));
    Odrv4 I__3025 (
            .O(N__25290),
            .I(n2199));
    InMux I__3024 (
            .O(N__25287),
            .I(n12658));
    InMux I__3023 (
            .O(N__25284),
            .I(n12659));
    InMux I__3022 (
            .O(N__25281),
            .I(N__25278));
    LocalMux I__3021 (
            .O(N__25278),
            .I(n2197));
    InMux I__3020 (
            .O(N__25275),
            .I(n12660));
    CascadeMux I__3019 (
            .O(N__25272),
            .I(N__25268));
    CascadeMux I__3018 (
            .O(N__25271),
            .I(N__25265));
    InMux I__3017 (
            .O(N__25268),
            .I(N__25262));
    InMux I__3016 (
            .O(N__25265),
            .I(N__25259));
    LocalMux I__3015 (
            .O(N__25262),
            .I(n2129));
    LocalMux I__3014 (
            .O(N__25259),
            .I(n2129));
    InMux I__3013 (
            .O(N__25254),
            .I(N__25251));
    LocalMux I__3012 (
            .O(N__25251),
            .I(n2196));
    InMux I__3011 (
            .O(N__25248),
            .I(n12661));
    InMux I__3010 (
            .O(N__25245),
            .I(N__25242));
    LocalMux I__3009 (
            .O(N__25242),
            .I(n3175));
    CascadeMux I__3008 (
            .O(N__25239),
            .I(n3108_cascade_));
    InMux I__3007 (
            .O(N__25236),
            .I(N__25232));
    CascadeMux I__3006 (
            .O(N__25235),
            .I(N__25228));
    LocalMux I__3005 (
            .O(N__25232),
            .I(N__25225));
    InMux I__3004 (
            .O(N__25231),
            .I(N__25222));
    InMux I__3003 (
            .O(N__25228),
            .I(N__25219));
    Odrv4 I__3002 (
            .O(N__25225),
            .I(n2232));
    LocalMux I__3001 (
            .O(N__25222),
            .I(n2232));
    LocalMux I__3000 (
            .O(N__25219),
            .I(n2232));
    InMux I__2999 (
            .O(N__25212),
            .I(N__25209));
    LocalMux I__2998 (
            .O(N__25209),
            .I(N__25205));
    CascadeMux I__2997 (
            .O(N__25208),
            .I(N__25202));
    Span4Mux_v I__2996 (
            .O(N__25205),
            .I(N__25198));
    InMux I__2995 (
            .O(N__25202),
            .I(N__25195));
    InMux I__2994 (
            .O(N__25201),
            .I(N__25192));
    Odrv4 I__2993 (
            .O(N__25198),
            .I(n2231));
    LocalMux I__2992 (
            .O(N__25195),
            .I(n2231));
    LocalMux I__2991 (
            .O(N__25192),
            .I(n2231));
    CascadeMux I__2990 (
            .O(N__25185),
            .I(N__25182));
    InMux I__2989 (
            .O(N__25182),
            .I(N__25179));
    LocalMux I__2988 (
            .O(N__25179),
            .I(N__25174));
    CascadeMux I__2987 (
            .O(N__25178),
            .I(N__25171));
    CascadeMux I__2986 (
            .O(N__25177),
            .I(N__25168));
    Span4Mux_v I__2985 (
            .O(N__25174),
            .I(N__25165));
    InMux I__2984 (
            .O(N__25171),
            .I(N__25162));
    InMux I__2983 (
            .O(N__25168),
            .I(N__25159));
    Odrv4 I__2982 (
            .O(N__25165),
            .I(n2221));
    LocalMux I__2981 (
            .O(N__25162),
            .I(n2221));
    LocalMux I__2980 (
            .O(N__25159),
            .I(n2221));
    CascadeMux I__2979 (
            .O(N__25152),
            .I(N__25147));
    InMux I__2978 (
            .O(N__25151),
            .I(N__25142));
    InMux I__2977 (
            .O(N__25150),
            .I(N__25142));
    InMux I__2976 (
            .O(N__25147),
            .I(N__25139));
    LocalMux I__2975 (
            .O(N__25142),
            .I(N__25136));
    LocalMux I__2974 (
            .O(N__25139),
            .I(N__25133));
    Odrv4 I__2973 (
            .O(N__25136),
            .I(n2229));
    Odrv4 I__2972 (
            .O(N__25133),
            .I(n2229));
    InMux I__2971 (
            .O(N__25128),
            .I(n12891));
    CascadeMux I__2970 (
            .O(N__25125),
            .I(N__25122));
    InMux I__2969 (
            .O(N__25122),
            .I(N__25119));
    LocalMux I__2968 (
            .O(N__25119),
            .I(n3075));
    InMux I__2967 (
            .O(N__25116),
            .I(N__25113));
    LocalMux I__2966 (
            .O(N__25113),
            .I(n3082));
    CascadeMux I__2965 (
            .O(N__25110),
            .I(N__25107));
    InMux I__2964 (
            .O(N__25107),
            .I(N__25104));
    LocalMux I__2963 (
            .O(N__25104),
            .I(n3074));
    InMux I__2962 (
            .O(N__25101),
            .I(N__25098));
    LocalMux I__2961 (
            .O(N__25098),
            .I(n3173));
    InMux I__2960 (
            .O(N__25095),
            .I(N__25092));
    LocalMux I__2959 (
            .O(N__25092),
            .I(n3174));
    InMux I__2958 (
            .O(N__25089),
            .I(N__25086));
    LocalMux I__2957 (
            .O(N__25086),
            .I(N__25083));
    Odrv4 I__2956 (
            .O(N__25083),
            .I(n3079));
    CascadeMux I__2955 (
            .O(N__25080),
            .I(N__25077));
    InMux I__2954 (
            .O(N__25077),
            .I(N__25074));
    LocalMux I__2953 (
            .O(N__25074),
            .I(N__25071));
    Odrv4 I__2952 (
            .O(N__25071),
            .I(n3078));
    InMux I__2951 (
            .O(N__25068),
            .I(N__25065));
    LocalMux I__2950 (
            .O(N__25065),
            .I(n3076));
    InMux I__2949 (
            .O(N__25062),
            .I(n12882));
    InMux I__2948 (
            .O(N__25059),
            .I(n12883));
    InMux I__2947 (
            .O(N__25056),
            .I(n12884));
    InMux I__2946 (
            .O(N__25053),
            .I(n12885));
    InMux I__2945 (
            .O(N__25050),
            .I(n12886));
    InMux I__2944 (
            .O(N__25047),
            .I(bfn_3_31_0_));
    InMux I__2943 (
            .O(N__25044),
            .I(n12888));
    InMux I__2942 (
            .O(N__25041),
            .I(n12889));
    InMux I__2941 (
            .O(N__25038),
            .I(n12890));
    CascadeMux I__2940 (
            .O(N__25035),
            .I(N__25032));
    InMux I__2939 (
            .O(N__25032),
            .I(N__25029));
    LocalMux I__2938 (
            .O(N__25029),
            .I(N__25026));
    Span4Mux_s2_h I__2937 (
            .O(N__25026),
            .I(N__25023));
    Odrv4 I__2936 (
            .O(N__25023),
            .I(n3090));
    InMux I__2935 (
            .O(N__25020),
            .I(n12874));
    CascadeMux I__2934 (
            .O(N__25017),
            .I(N__25014));
    InMux I__2933 (
            .O(N__25014),
            .I(N__25011));
    LocalMux I__2932 (
            .O(N__25011),
            .I(N__25007));
    InMux I__2931 (
            .O(N__25010),
            .I(N__25003));
    Span4Mux_h I__2930 (
            .O(N__25007),
            .I(N__25000));
    InMux I__2929 (
            .O(N__25006),
            .I(N__24997));
    LocalMux I__2928 (
            .O(N__25003),
            .I(n3022));
    Odrv4 I__2927 (
            .O(N__25000),
            .I(n3022));
    LocalMux I__2926 (
            .O(N__24997),
            .I(n3022));
    CascadeMux I__2925 (
            .O(N__24990),
            .I(N__24987));
    InMux I__2924 (
            .O(N__24987),
            .I(N__24984));
    LocalMux I__2923 (
            .O(N__24984),
            .I(n3089));
    InMux I__2922 (
            .O(N__24981),
            .I(n12875));
    CascadeMux I__2921 (
            .O(N__24978),
            .I(N__24974));
    CascadeMux I__2920 (
            .O(N__24977),
            .I(N__24971));
    InMux I__2919 (
            .O(N__24974),
            .I(N__24968));
    InMux I__2918 (
            .O(N__24971),
            .I(N__24965));
    LocalMux I__2917 (
            .O(N__24968),
            .I(N__24962));
    LocalMux I__2916 (
            .O(N__24965),
            .I(N__24959));
    Span4Mux_s1_h I__2915 (
            .O(N__24962),
            .I(N__24954));
    Span4Mux_h I__2914 (
            .O(N__24959),
            .I(N__24954));
    Odrv4 I__2913 (
            .O(N__24954),
            .I(n3021));
    InMux I__2912 (
            .O(N__24951),
            .I(N__24948));
    LocalMux I__2911 (
            .O(N__24948),
            .I(N__24945));
    Odrv4 I__2910 (
            .O(N__24945),
            .I(n3088));
    InMux I__2909 (
            .O(N__24942),
            .I(n12876));
    CascadeMux I__2908 (
            .O(N__24939),
            .I(N__24936));
    InMux I__2907 (
            .O(N__24936),
            .I(N__24931));
    InMux I__2906 (
            .O(N__24935),
            .I(N__24928));
    InMux I__2905 (
            .O(N__24934),
            .I(N__24925));
    LocalMux I__2904 (
            .O(N__24931),
            .I(N__24922));
    LocalMux I__2903 (
            .O(N__24928),
            .I(N__24919));
    LocalMux I__2902 (
            .O(N__24925),
            .I(n3020));
    Odrv4 I__2901 (
            .O(N__24922),
            .I(n3020));
    Odrv12 I__2900 (
            .O(N__24919),
            .I(n3020));
    InMux I__2899 (
            .O(N__24912),
            .I(N__24909));
    LocalMux I__2898 (
            .O(N__24909),
            .I(n3087));
    InMux I__2897 (
            .O(N__24906),
            .I(n12877));
    InMux I__2896 (
            .O(N__24903),
            .I(N__24900));
    LocalMux I__2895 (
            .O(N__24900),
            .I(N__24897));
    Odrv4 I__2894 (
            .O(N__24897),
            .I(n3086));
    InMux I__2893 (
            .O(N__24894),
            .I(n12878));
    InMux I__2892 (
            .O(N__24891),
            .I(bfn_3_30_0_));
    InMux I__2891 (
            .O(N__24888),
            .I(N__24885));
    LocalMux I__2890 (
            .O(N__24885),
            .I(N__24881));
    InMux I__2889 (
            .O(N__24884),
            .I(N__24877));
    Span4Mux_h I__2888 (
            .O(N__24881),
            .I(N__24874));
    InMux I__2887 (
            .O(N__24880),
            .I(N__24871));
    LocalMux I__2886 (
            .O(N__24877),
            .I(n3017));
    Odrv4 I__2885 (
            .O(N__24874),
            .I(n3017));
    LocalMux I__2884 (
            .O(N__24871),
            .I(n3017));
    InMux I__2883 (
            .O(N__24864),
            .I(N__24861));
    LocalMux I__2882 (
            .O(N__24861),
            .I(N__24858));
    Odrv4 I__2881 (
            .O(N__24858),
            .I(n3084));
    InMux I__2880 (
            .O(N__24855),
            .I(n12880));
    InMux I__2879 (
            .O(N__24852),
            .I(n12881));
    InMux I__2878 (
            .O(N__24849),
            .I(n12866));
    InMux I__2877 (
            .O(N__24846),
            .I(n12867));
    InMux I__2876 (
            .O(N__24843),
            .I(N__24840));
    LocalMux I__2875 (
            .O(N__24840),
            .I(N__24837));
    Odrv12 I__2874 (
            .O(N__24837),
            .I(n3096));
    InMux I__2873 (
            .O(N__24834),
            .I(n12868));
    CascadeMux I__2872 (
            .O(N__24831),
            .I(N__24827));
    InMux I__2871 (
            .O(N__24830),
            .I(N__24824));
    InMux I__2870 (
            .O(N__24827),
            .I(N__24821));
    LocalMux I__2869 (
            .O(N__24824),
            .I(N__24818));
    LocalMux I__2868 (
            .O(N__24821),
            .I(n3028));
    Odrv12 I__2867 (
            .O(N__24818),
            .I(n3028));
    InMux I__2866 (
            .O(N__24813),
            .I(N__24810));
    LocalMux I__2865 (
            .O(N__24810),
            .I(n3095));
    InMux I__2864 (
            .O(N__24807),
            .I(n12869));
    InMux I__2863 (
            .O(N__24804),
            .I(N__24801));
    LocalMux I__2862 (
            .O(N__24801),
            .I(N__24798));
    Odrv12 I__2861 (
            .O(N__24798),
            .I(n3094));
    InMux I__2860 (
            .O(N__24795),
            .I(n12870));
    CascadeMux I__2859 (
            .O(N__24792),
            .I(N__24789));
    InMux I__2858 (
            .O(N__24789),
            .I(N__24785));
    InMux I__2857 (
            .O(N__24788),
            .I(N__24782));
    LocalMux I__2856 (
            .O(N__24785),
            .I(N__24779));
    LocalMux I__2855 (
            .O(N__24782),
            .I(N__24775));
    Span4Mux_h I__2854 (
            .O(N__24779),
            .I(N__24772));
    InMux I__2853 (
            .O(N__24778),
            .I(N__24769));
    Odrv4 I__2852 (
            .O(N__24775),
            .I(n3026));
    Odrv4 I__2851 (
            .O(N__24772),
            .I(n3026));
    LocalMux I__2850 (
            .O(N__24769),
            .I(n3026));
    CascadeMux I__2849 (
            .O(N__24762),
            .I(N__24759));
    InMux I__2848 (
            .O(N__24759),
            .I(N__24756));
    LocalMux I__2847 (
            .O(N__24756),
            .I(n3093));
    InMux I__2846 (
            .O(N__24753),
            .I(bfn_3_29_0_));
    CascadeMux I__2845 (
            .O(N__24750),
            .I(N__24747));
    InMux I__2844 (
            .O(N__24747),
            .I(N__24743));
    InMux I__2843 (
            .O(N__24746),
            .I(N__24740));
    LocalMux I__2842 (
            .O(N__24743),
            .I(N__24737));
    LocalMux I__2841 (
            .O(N__24740),
            .I(N__24731));
    Span4Mux_h I__2840 (
            .O(N__24737),
            .I(N__24731));
    InMux I__2839 (
            .O(N__24736),
            .I(N__24728));
    Odrv4 I__2838 (
            .O(N__24731),
            .I(n3025));
    LocalMux I__2837 (
            .O(N__24728),
            .I(n3025));
    InMux I__2836 (
            .O(N__24723),
            .I(N__24720));
    LocalMux I__2835 (
            .O(N__24720),
            .I(N__24717));
    Odrv4 I__2834 (
            .O(N__24717),
            .I(n3092));
    InMux I__2833 (
            .O(N__24714),
            .I(n12872));
    CascadeMux I__2832 (
            .O(N__24711),
            .I(N__24708));
    InMux I__2831 (
            .O(N__24708),
            .I(N__24704));
    InMux I__2830 (
            .O(N__24707),
            .I(N__24701));
    LocalMux I__2829 (
            .O(N__24704),
            .I(N__24698));
    LocalMux I__2828 (
            .O(N__24701),
            .I(N__24695));
    Span4Mux_v I__2827 (
            .O(N__24698),
            .I(N__24692));
    Odrv12 I__2826 (
            .O(N__24695),
            .I(n3024));
    Odrv4 I__2825 (
            .O(N__24692),
            .I(n3024));
    CascadeMux I__2824 (
            .O(N__24687),
            .I(N__24684));
    InMux I__2823 (
            .O(N__24684),
            .I(N__24681));
    LocalMux I__2822 (
            .O(N__24681),
            .I(N__24678));
    Odrv4 I__2821 (
            .O(N__24678),
            .I(n3091));
    InMux I__2820 (
            .O(N__24675),
            .I(n12873));
    CascadeMux I__2819 (
            .O(N__24672),
            .I(n3028_cascade_));
    CascadeMux I__2818 (
            .O(N__24669),
            .I(N__24666));
    InMux I__2817 (
            .O(N__24666),
            .I(N__24663));
    LocalMux I__2816 (
            .O(N__24663),
            .I(n2988));
    InMux I__2815 (
            .O(N__24660),
            .I(N__24657));
    LocalMux I__2814 (
            .O(N__24657),
            .I(N__24654));
    Span4Mux_v I__2813 (
            .O(N__24654),
            .I(N__24651));
    Odrv4 I__2812 (
            .O(N__24651),
            .I(n2880));
    InMux I__2811 (
            .O(N__24648),
            .I(N__24645));
    LocalMux I__2810 (
            .O(N__24645),
            .I(n2979));
    CascadeMux I__2809 (
            .O(N__24642),
            .I(n2912_cascade_));
    CascadeMux I__2808 (
            .O(N__24639),
            .I(N__24636));
    InMux I__2807 (
            .O(N__24636),
            .I(N__24633));
    LocalMux I__2806 (
            .O(N__24633),
            .I(n2983));
    InMux I__2805 (
            .O(N__24630),
            .I(bfn_3_28_0_));
    InMux I__2804 (
            .O(N__24627),
            .I(n12864));
    InMux I__2803 (
            .O(N__24624),
            .I(n12865));
    CascadeMux I__2802 (
            .O(N__24621),
            .I(N__24618));
    InMux I__2801 (
            .O(N__24618),
            .I(N__24613));
    InMux I__2800 (
            .O(N__24617),
            .I(N__24608));
    InMux I__2799 (
            .O(N__24616),
            .I(N__24608));
    LocalMux I__2798 (
            .O(N__24613),
            .I(n2823));
    LocalMux I__2797 (
            .O(N__24608),
            .I(n2823));
    CascadeMux I__2796 (
            .O(N__24603),
            .I(N__24600));
    InMux I__2795 (
            .O(N__24600),
            .I(N__24597));
    LocalMux I__2794 (
            .O(N__24597),
            .I(N__24594));
    Span4Mux_v I__2793 (
            .O(N__24594),
            .I(N__24591));
    Odrv4 I__2792 (
            .O(N__24591),
            .I(n2890));
    InMux I__2791 (
            .O(N__24588),
            .I(N__24585));
    LocalMux I__2790 (
            .O(N__24585),
            .I(N__24581));
    CascadeMux I__2789 (
            .O(N__24584),
            .I(N__24578));
    Span4Mux_v I__2788 (
            .O(N__24581),
            .I(N__24574));
    InMux I__2787 (
            .O(N__24578),
            .I(N__24571));
    InMux I__2786 (
            .O(N__24577),
            .I(N__24568));
    Odrv4 I__2785 (
            .O(N__24574),
            .I(n2827));
    LocalMux I__2784 (
            .O(N__24571),
            .I(n2827));
    LocalMux I__2783 (
            .O(N__24568),
            .I(n2827));
    CascadeMux I__2782 (
            .O(N__24561),
            .I(N__24558));
    InMux I__2781 (
            .O(N__24558),
            .I(N__24555));
    LocalMux I__2780 (
            .O(N__24555),
            .I(N__24552));
    Span4Mux_v I__2779 (
            .O(N__24552),
            .I(N__24549));
    Odrv4 I__2778 (
            .O(N__24549),
            .I(n2894));
    InMux I__2777 (
            .O(N__24546),
            .I(N__24543));
    LocalMux I__2776 (
            .O(N__24543),
            .I(N__24539));
    CascadeMux I__2775 (
            .O(N__24542),
            .I(N__24536));
    Span4Mux_v I__2774 (
            .O(N__24539),
            .I(N__24532));
    InMux I__2773 (
            .O(N__24536),
            .I(N__24529));
    InMux I__2772 (
            .O(N__24535),
            .I(N__24526));
    Odrv4 I__2771 (
            .O(N__24532),
            .I(n2822));
    LocalMux I__2770 (
            .O(N__24529),
            .I(n2822));
    LocalMux I__2769 (
            .O(N__24526),
            .I(n2822));
    CascadeMux I__2768 (
            .O(N__24519),
            .I(N__24516));
    InMux I__2767 (
            .O(N__24516),
            .I(N__24513));
    LocalMux I__2766 (
            .O(N__24513),
            .I(N__24510));
    Span4Mux_h I__2765 (
            .O(N__24510),
            .I(N__24507));
    Odrv4 I__2764 (
            .O(N__24507),
            .I(n2889));
    CascadeMux I__2763 (
            .O(N__24504),
            .I(N__24501));
    InMux I__2762 (
            .O(N__24501),
            .I(N__24498));
    LocalMux I__2761 (
            .O(N__24498),
            .I(n2982));
    CascadeMux I__2760 (
            .O(N__24495),
            .I(N__24492));
    InMux I__2759 (
            .O(N__24492),
            .I(N__24489));
    LocalMux I__2758 (
            .O(N__24489),
            .I(n2986));
    InMux I__2757 (
            .O(N__24486),
            .I(N__24483));
    LocalMux I__2756 (
            .O(N__24483),
            .I(N__24480));
    Span4Mux_h I__2755 (
            .O(N__24480),
            .I(N__24477));
    Span4Mux_s0_h I__2754 (
            .O(N__24477),
            .I(N__24474));
    Odrv4 I__2753 (
            .O(N__24474),
            .I(n2879));
    InMux I__2752 (
            .O(N__24471),
            .I(N__24468));
    LocalMux I__2751 (
            .O(N__24468),
            .I(N__24464));
    InMux I__2750 (
            .O(N__24467),
            .I(N__24460));
    Span4Mux_v I__2749 (
            .O(N__24464),
            .I(N__24457));
    InMux I__2748 (
            .O(N__24463),
            .I(N__24454));
    LocalMux I__2747 (
            .O(N__24460),
            .I(N__24451));
    Odrv4 I__2746 (
            .O(N__24457),
            .I(n2710));
    LocalMux I__2745 (
            .O(N__24454),
            .I(n2710));
    Odrv12 I__2744 (
            .O(N__24451),
            .I(n2710));
    CascadeMux I__2743 (
            .O(N__24444),
            .I(N__24441));
    InMux I__2742 (
            .O(N__24441),
            .I(N__24438));
    LocalMux I__2741 (
            .O(N__24438),
            .I(N__24435));
    Span4Mux_v I__2740 (
            .O(N__24435),
            .I(N__24432));
    Span4Mux_v I__2739 (
            .O(N__24432),
            .I(N__24429));
    Odrv4 I__2738 (
            .O(N__24429),
            .I(n2777));
    InMux I__2737 (
            .O(N__24426),
            .I(N__24423));
    LocalMux I__2736 (
            .O(N__24423),
            .I(N__24420));
    Odrv4 I__2735 (
            .O(N__24420),
            .I(n2996));
    InMux I__2734 (
            .O(N__24417),
            .I(N__24412));
    InMux I__2733 (
            .O(N__24416),
            .I(N__24409));
    InMux I__2732 (
            .O(N__24415),
            .I(N__24406));
    LocalMux I__2731 (
            .O(N__24412),
            .I(N__24403));
    LocalMux I__2730 (
            .O(N__24409),
            .I(N__24398));
    LocalMux I__2729 (
            .O(N__24406),
            .I(N__24398));
    Odrv4 I__2728 (
            .O(N__24403),
            .I(n2713));
    Odrv4 I__2727 (
            .O(N__24398),
            .I(n2713));
    InMux I__2726 (
            .O(N__24393),
            .I(N__24390));
    LocalMux I__2725 (
            .O(N__24390),
            .I(N__24387));
    Span4Mux_v I__2724 (
            .O(N__24387),
            .I(N__24384));
    Odrv4 I__2723 (
            .O(N__24384),
            .I(n2780));
    InMux I__2722 (
            .O(N__24381),
            .I(N__24378));
    LocalMux I__2721 (
            .O(N__24378),
            .I(N__24375));
    Span4Mux_v I__2720 (
            .O(N__24375),
            .I(N__24372));
    Odrv4 I__2719 (
            .O(N__24372),
            .I(n2798));
    CascadeMux I__2718 (
            .O(N__24369),
            .I(N__24365));
    CascadeMux I__2717 (
            .O(N__24368),
            .I(N__24362));
    InMux I__2716 (
            .O(N__24365),
            .I(N__24359));
    InMux I__2715 (
            .O(N__24362),
            .I(N__24356));
    LocalMux I__2714 (
            .O(N__24359),
            .I(N__24353));
    LocalMux I__2713 (
            .O(N__24356),
            .I(N__24349));
    Span12Mux_s2_h I__2712 (
            .O(N__24353),
            .I(N__24346));
    InMux I__2711 (
            .O(N__24352),
            .I(N__24343));
    Odrv4 I__2710 (
            .O(N__24349),
            .I(n2731));
    Odrv12 I__2709 (
            .O(N__24346),
            .I(n2731));
    LocalMux I__2708 (
            .O(N__24343),
            .I(n2731));
    InMux I__2707 (
            .O(N__24336),
            .I(N__24333));
    LocalMux I__2706 (
            .O(N__24333),
            .I(N__24330));
    Span4Mux_v I__2705 (
            .O(N__24330),
            .I(N__24327));
    Span4Mux_v I__2704 (
            .O(N__24327),
            .I(N__24324));
    Odrv4 I__2703 (
            .O(N__24324),
            .I(n2680));
    InMux I__2702 (
            .O(N__24321),
            .I(N__24318));
    LocalMux I__2701 (
            .O(N__24318),
            .I(N__24315));
    Span4Mux_h I__2700 (
            .O(N__24315),
            .I(N__24312));
    Odrv4 I__2699 (
            .O(N__24312),
            .I(n2887));
    InMux I__2698 (
            .O(N__24309),
            .I(N__24304));
    InMux I__2697 (
            .O(N__24308),
            .I(N__24299));
    InMux I__2696 (
            .O(N__24307),
            .I(N__24299));
    LocalMux I__2695 (
            .O(N__24304),
            .I(n2820));
    LocalMux I__2694 (
            .O(N__24299),
            .I(n2820));
    CascadeMux I__2693 (
            .O(N__24294),
            .I(n14690_cascade_));
    InMux I__2692 (
            .O(N__24291),
            .I(N__24288));
    LocalMux I__2691 (
            .O(N__24288),
            .I(N__24285));
    Odrv4 I__2690 (
            .O(N__24285),
            .I(n14688));
    CascadeMux I__2689 (
            .O(N__24282),
            .I(n14696_cascade_));
    InMux I__2688 (
            .O(N__24279),
            .I(N__24274));
    InMux I__2687 (
            .O(N__24278),
            .I(N__24271));
    InMux I__2686 (
            .O(N__24277),
            .I(N__24268));
    LocalMux I__2685 (
            .O(N__24274),
            .I(N__24265));
    LocalMux I__2684 (
            .O(N__24271),
            .I(N__24262));
    LocalMux I__2683 (
            .O(N__24268),
            .I(N__24259));
    Span4Mux_v I__2682 (
            .O(N__24265),
            .I(N__24256));
    Span4Mux_h I__2681 (
            .O(N__24262),
            .I(N__24253));
    Odrv4 I__2680 (
            .O(N__24259),
            .I(n2714));
    Odrv4 I__2679 (
            .O(N__24256),
            .I(n2714));
    Odrv4 I__2678 (
            .O(N__24253),
            .I(n2714));
    CascadeMux I__2677 (
            .O(N__24246),
            .I(N__24243));
    InMux I__2676 (
            .O(N__24243),
            .I(N__24240));
    LocalMux I__2675 (
            .O(N__24240),
            .I(N__24237));
    Span4Mux_v I__2674 (
            .O(N__24237),
            .I(N__24234));
    Odrv4 I__2673 (
            .O(N__24234),
            .I(n2781));
    InMux I__2672 (
            .O(N__24231),
            .I(N__24228));
    LocalMux I__2671 (
            .O(N__24228),
            .I(N__24224));
    InMux I__2670 (
            .O(N__24227),
            .I(N__24221));
    Span4Mux_v I__2669 (
            .O(N__24224),
            .I(N__24217));
    LocalMux I__2668 (
            .O(N__24221),
            .I(N__24214));
    InMux I__2667 (
            .O(N__24220),
            .I(N__24211));
    Odrv4 I__2666 (
            .O(N__24217),
            .I(n2720));
    Odrv4 I__2665 (
            .O(N__24214),
            .I(n2720));
    LocalMux I__2664 (
            .O(N__24211),
            .I(n2720));
    CascadeMux I__2663 (
            .O(N__24204),
            .I(N__24201));
    InMux I__2662 (
            .O(N__24201),
            .I(N__24198));
    LocalMux I__2661 (
            .O(N__24198),
            .I(N__24195));
    Span4Mux_v I__2660 (
            .O(N__24195),
            .I(N__24192));
    Odrv4 I__2659 (
            .O(N__24192),
            .I(n2787));
    CascadeMux I__2658 (
            .O(N__24189),
            .I(n14660_cascade_));
    InMux I__2657 (
            .O(N__24186),
            .I(N__24183));
    LocalMux I__2656 (
            .O(N__24183),
            .I(n14674));
    CascadeMux I__2655 (
            .O(N__24180),
            .I(n2643_cascade_));
    InMux I__2654 (
            .O(N__24177),
            .I(N__24174));
    LocalMux I__2653 (
            .O(N__24174),
            .I(N__24171));
    Span12Mux_v I__2652 (
            .O(N__24171),
            .I(N__24168));
    Odrv12 I__2651 (
            .O(N__24168),
            .I(n2686));
    InMux I__2650 (
            .O(N__24165),
            .I(N__24162));
    LocalMux I__2649 (
            .O(N__24162),
            .I(N__24159));
    Span4Mux_v I__2648 (
            .O(N__24159),
            .I(N__24154));
    InMux I__2647 (
            .O(N__24158),
            .I(N__24149));
    InMux I__2646 (
            .O(N__24157),
            .I(N__24149));
    Odrv4 I__2645 (
            .O(N__24154),
            .I(n2718));
    LocalMux I__2644 (
            .O(N__24149),
            .I(n2718));
    InMux I__2643 (
            .O(N__24144),
            .I(N__24141));
    LocalMux I__2642 (
            .O(N__24141),
            .I(N__24138));
    Span4Mux_v I__2641 (
            .O(N__24138),
            .I(N__24135));
    Span4Mux_v I__2640 (
            .O(N__24135),
            .I(N__24132));
    Odrv4 I__2639 (
            .O(N__24132),
            .I(n2690));
    CascadeMux I__2638 (
            .O(N__24129),
            .I(N__24125));
    InMux I__2637 (
            .O(N__24128),
            .I(N__24121));
    InMux I__2636 (
            .O(N__24125),
            .I(N__24116));
    InMux I__2635 (
            .O(N__24124),
            .I(N__24116));
    LocalMux I__2634 (
            .O(N__24121),
            .I(N__24113));
    LocalMux I__2633 (
            .O(N__24116),
            .I(N__24110));
    Span4Mux_v I__2632 (
            .O(N__24113),
            .I(N__24107));
    Odrv4 I__2631 (
            .O(N__24110),
            .I(n2623));
    Odrv4 I__2630 (
            .O(N__24107),
            .I(n2623));
    CascadeMux I__2629 (
            .O(N__24102),
            .I(N__24099));
    InMux I__2628 (
            .O(N__24099),
            .I(N__24096));
    LocalMux I__2627 (
            .O(N__24096),
            .I(N__24093));
    Span12Mux_s2_h I__2626 (
            .O(N__24093),
            .I(N__24088));
    InMux I__2625 (
            .O(N__24092),
            .I(N__24083));
    InMux I__2624 (
            .O(N__24091),
            .I(N__24083));
    Odrv12 I__2623 (
            .O(N__24088),
            .I(n2722));
    LocalMux I__2622 (
            .O(N__24083),
            .I(n2722));
    CascadeMux I__2621 (
            .O(N__24078),
            .I(N__24075));
    InMux I__2620 (
            .O(N__24075),
            .I(N__24071));
    InMux I__2619 (
            .O(N__24074),
            .I(N__24068));
    LocalMux I__2618 (
            .O(N__24071),
            .I(N__24065));
    LocalMux I__2617 (
            .O(N__24068),
            .I(N__24062));
    Span4Mux_v I__2616 (
            .O(N__24065),
            .I(N__24059));
    Odrv4 I__2615 (
            .O(N__24062),
            .I(n2732));
    Odrv4 I__2614 (
            .O(N__24059),
            .I(n2732));
    CascadeMux I__2613 (
            .O(N__24054),
            .I(N__24051));
    InMux I__2612 (
            .O(N__24051),
            .I(N__24048));
    LocalMux I__2611 (
            .O(N__24048),
            .I(N__24045));
    Span4Mux_v I__2610 (
            .O(N__24045),
            .I(N__24042));
    Odrv4 I__2609 (
            .O(N__24042),
            .I(n2799));
    InMux I__2608 (
            .O(N__24039),
            .I(N__24036));
    LocalMux I__2607 (
            .O(N__24036),
            .I(N__24032));
    InMux I__2606 (
            .O(N__24035),
            .I(N__24029));
    Span4Mux_v I__2605 (
            .O(N__24032),
            .I(N__24026));
    LocalMux I__2604 (
            .O(N__24029),
            .I(n2711));
    Odrv4 I__2603 (
            .O(N__24026),
            .I(n2711));
    InMux I__2602 (
            .O(N__24021),
            .I(N__24018));
    LocalMux I__2601 (
            .O(N__24018),
            .I(N__24015));
    Span4Mux_h I__2600 (
            .O(N__24015),
            .I(N__24012));
    Span4Mux_s1_h I__2599 (
            .O(N__24012),
            .I(N__24009));
    Span4Mux_v I__2598 (
            .O(N__24009),
            .I(N__24006));
    Odrv4 I__2597 (
            .O(N__24006),
            .I(n2778));
    InMux I__2596 (
            .O(N__24003),
            .I(N__24000));
    LocalMux I__2595 (
            .O(N__24000),
            .I(N__23997));
    Span4Mux_v I__2594 (
            .O(N__23997),
            .I(N__23994));
    Odrv4 I__2593 (
            .O(N__23994),
            .I(n2786));
    CascadeMux I__2592 (
            .O(N__23991),
            .I(N__23987));
    InMux I__2591 (
            .O(N__23990),
            .I(N__23984));
    InMux I__2590 (
            .O(N__23987),
            .I(N__23980));
    LocalMux I__2589 (
            .O(N__23984),
            .I(N__23977));
    InMux I__2588 (
            .O(N__23983),
            .I(N__23974));
    LocalMux I__2587 (
            .O(N__23980),
            .I(n2719));
    Odrv12 I__2586 (
            .O(N__23977),
            .I(n2719));
    LocalMux I__2585 (
            .O(N__23974),
            .I(n2719));
    InMux I__2584 (
            .O(N__23967),
            .I(N__23964));
    LocalMux I__2583 (
            .O(N__23964),
            .I(N__23961));
    Span4Mux_v I__2582 (
            .O(N__23961),
            .I(N__23958));
    Span4Mux_v I__2581 (
            .O(N__23958),
            .I(N__23955));
    Odrv4 I__2580 (
            .O(N__23955),
            .I(n2685));
    InMux I__2579 (
            .O(N__23952),
            .I(N__23949));
    LocalMux I__2578 (
            .O(N__23949),
            .I(N__23946));
    Span4Mux_v I__2577 (
            .O(N__23946),
            .I(N__23942));
    InMux I__2576 (
            .O(N__23945),
            .I(N__23939));
    Odrv4 I__2575 (
            .O(N__23942),
            .I(n2717));
    LocalMux I__2574 (
            .O(N__23939),
            .I(n2717));
    InMux I__2573 (
            .O(N__23934),
            .I(N__23931));
    LocalMux I__2572 (
            .O(N__23931),
            .I(N__23928));
    Span4Mux_v I__2571 (
            .O(N__23928),
            .I(N__23925));
    Odrv4 I__2570 (
            .O(N__23925),
            .I(n2784));
    CascadeMux I__2569 (
            .O(N__23922),
            .I(n2717_cascade_));
    CascadeMux I__2568 (
            .O(N__23919),
            .I(n2732_cascade_));
    InMux I__2567 (
            .O(N__23916),
            .I(N__23912));
    InMux I__2566 (
            .O(N__23915),
            .I(N__23909));
    LocalMux I__2565 (
            .O(N__23912),
            .I(N__23906));
    LocalMux I__2564 (
            .O(N__23909),
            .I(N__23902));
    Span4Mux_v I__2563 (
            .O(N__23906),
            .I(N__23899));
    InMux I__2562 (
            .O(N__23905),
            .I(N__23896));
    Odrv4 I__2561 (
            .O(N__23902),
            .I(n2729));
    Odrv4 I__2560 (
            .O(N__23899),
            .I(n2729));
    LocalMux I__2559 (
            .O(N__23896),
            .I(n2729));
    CascadeMux I__2558 (
            .O(N__23889),
            .I(n11957_cascade_));
    InMux I__2557 (
            .O(N__23886),
            .I(N__23883));
    LocalMux I__2556 (
            .O(N__23883),
            .I(n13808));
    CascadeMux I__2555 (
            .O(N__23880),
            .I(N__23877));
    InMux I__2554 (
            .O(N__23877),
            .I(N__23874));
    LocalMux I__2553 (
            .O(N__23874),
            .I(N__23871));
    Span4Mux_v I__2552 (
            .O(N__23871),
            .I(N__23867));
    InMux I__2551 (
            .O(N__23870),
            .I(N__23864));
    Odrv4 I__2550 (
            .O(N__23867),
            .I(n2621));
    LocalMux I__2549 (
            .O(N__23864),
            .I(n2621));
    InMux I__2548 (
            .O(N__23859),
            .I(N__23856));
    LocalMux I__2547 (
            .O(N__23856),
            .I(n14668));
    InMux I__2546 (
            .O(N__23853),
            .I(N__23850));
    LocalMux I__2545 (
            .O(N__23850),
            .I(N__23847));
    Span4Mux_v I__2544 (
            .O(N__23847),
            .I(N__23844));
    Span4Mux_v I__2543 (
            .O(N__23844),
            .I(N__23841));
    Odrv4 I__2542 (
            .O(N__23841),
            .I(n2698));
    CascadeMux I__2541 (
            .O(N__23838),
            .I(N__23835));
    InMux I__2540 (
            .O(N__23835),
            .I(N__23832));
    LocalMux I__2539 (
            .O(N__23832),
            .I(N__23828));
    InMux I__2538 (
            .O(N__23831),
            .I(N__23824));
    Span4Mux_v I__2537 (
            .O(N__23828),
            .I(N__23821));
    InMux I__2536 (
            .O(N__23827),
            .I(N__23818));
    LocalMux I__2535 (
            .O(N__23824),
            .I(n2730));
    Odrv4 I__2534 (
            .O(N__23821),
            .I(n2730));
    LocalMux I__2533 (
            .O(N__23818),
            .I(n2730));
    InMux I__2532 (
            .O(N__23811),
            .I(N__23808));
    LocalMux I__2531 (
            .O(N__23808),
            .I(N__23805));
    Span4Mux_v I__2530 (
            .O(N__23805),
            .I(N__23802));
    Span4Mux_v I__2529 (
            .O(N__23802),
            .I(N__23799));
    Odrv4 I__2528 (
            .O(N__23799),
            .I(n2699));
    InMux I__2527 (
            .O(N__23796),
            .I(N__23793));
    LocalMux I__2526 (
            .O(N__23793),
            .I(N__23790));
    Span4Mux_h I__2525 (
            .O(N__23790),
            .I(N__23787));
    Span4Mux_v I__2524 (
            .O(N__23787),
            .I(N__23784));
    Span4Mux_v I__2523 (
            .O(N__23784),
            .I(N__23781));
    Odrv4 I__2522 (
            .O(N__23781),
            .I(n2701));
    CascadeMux I__2521 (
            .O(N__23778),
            .I(n14650_cascade_));
    CascadeMux I__2520 (
            .O(N__23775),
            .I(n14654_cascade_));
    InMux I__2519 (
            .O(N__23772),
            .I(N__23769));
    LocalMux I__2518 (
            .O(N__23769),
            .I(N__23766));
    Span4Mux_v I__2517 (
            .O(N__23766),
            .I(N__23763));
    Odrv4 I__2516 (
            .O(N__23763),
            .I(n2689));
    CascadeMux I__2515 (
            .O(N__23760),
            .I(n2622_cascade_));
    InMux I__2514 (
            .O(N__23757),
            .I(N__23753));
    CascadeMux I__2513 (
            .O(N__23756),
            .I(N__23750));
    LocalMux I__2512 (
            .O(N__23753),
            .I(N__23747));
    InMux I__2511 (
            .O(N__23750),
            .I(N__23744));
    Span4Mux_v I__2510 (
            .O(N__23747),
            .I(N__23741));
    LocalMux I__2509 (
            .O(N__23744),
            .I(N__23738));
    Odrv4 I__2508 (
            .O(N__23741),
            .I(n2721));
    Odrv4 I__2507 (
            .O(N__23738),
            .I(n2721));
    CascadeMux I__2506 (
            .O(N__23733),
            .I(N__23730));
    InMux I__2505 (
            .O(N__23730),
            .I(N__23727));
    LocalMux I__2504 (
            .O(N__23727),
            .I(N__23723));
    InMux I__2503 (
            .O(N__23726),
            .I(N__23720));
    Odrv12 I__2502 (
            .O(N__23723),
            .I(n2728));
    LocalMux I__2501 (
            .O(N__23720),
            .I(n2728));
    CascadeMux I__2500 (
            .O(N__23715),
            .I(N__23712));
    InMux I__2499 (
            .O(N__23712),
            .I(N__23709));
    LocalMux I__2498 (
            .O(N__23709),
            .I(N__23705));
    InMux I__2497 (
            .O(N__23708),
            .I(N__23702));
    Odrv4 I__2496 (
            .O(N__23705),
            .I(n2726));
    LocalMux I__2495 (
            .O(N__23702),
            .I(n2726));
    CascadeMux I__2494 (
            .O(N__23697),
            .I(n2721_cascade_));
    InMux I__2493 (
            .O(N__23694),
            .I(N__23691));
    LocalMux I__2492 (
            .O(N__23691),
            .I(N__23688));
    Odrv4 I__2491 (
            .O(N__23688),
            .I(n14348));
    InMux I__2490 (
            .O(N__23685),
            .I(N__23682));
    LocalMux I__2489 (
            .O(N__23682),
            .I(N__23679));
    Odrv4 I__2488 (
            .O(N__23679),
            .I(n2383));
    CascadeMux I__2487 (
            .O(N__23676),
            .I(N__23673));
    InMux I__2486 (
            .O(N__23673),
            .I(N__23670));
    LocalMux I__2485 (
            .O(N__23670),
            .I(N__23667));
    Span4Mux_v I__2484 (
            .O(N__23667),
            .I(N__23663));
    InMux I__2483 (
            .O(N__23666),
            .I(N__23660));
    Odrv4 I__2482 (
            .O(N__23663),
            .I(n2622));
    LocalMux I__2481 (
            .O(N__23660),
            .I(n2622));
    CascadeMux I__2480 (
            .O(N__23655),
            .I(n2628_cascade_));
    InMux I__2479 (
            .O(N__23652),
            .I(N__23649));
    LocalMux I__2478 (
            .O(N__23649),
            .I(N__23646));
    Span4Mux_v I__2477 (
            .O(N__23646),
            .I(N__23643));
    Span4Mux_v I__2476 (
            .O(N__23643),
            .I(N__23640));
    Odrv4 I__2475 (
            .O(N__23640),
            .I(n2692));
    CascadeMux I__2474 (
            .O(N__23637),
            .I(N__23633));
    CascadeMux I__2473 (
            .O(N__23636),
            .I(N__23630));
    InMux I__2472 (
            .O(N__23633),
            .I(N__23627));
    InMux I__2471 (
            .O(N__23630),
            .I(N__23624));
    LocalMux I__2470 (
            .O(N__23627),
            .I(N__23621));
    LocalMux I__2469 (
            .O(N__23624),
            .I(N__23617));
    Span4Mux_s3_h I__2468 (
            .O(N__23621),
            .I(N__23614));
    InMux I__2467 (
            .O(N__23620),
            .I(N__23611));
    Odrv4 I__2466 (
            .O(N__23617),
            .I(n2724));
    Odrv4 I__2465 (
            .O(N__23614),
            .I(n2724));
    LocalMux I__2464 (
            .O(N__23611),
            .I(n2724));
    InMux I__2463 (
            .O(N__23604),
            .I(N__23601));
    LocalMux I__2462 (
            .O(N__23601),
            .I(N__23598));
    Span4Mux_v I__2461 (
            .O(N__23598),
            .I(N__23595));
    Span4Mux_v I__2460 (
            .O(N__23595),
            .I(N__23592));
    Odrv4 I__2459 (
            .O(N__23592),
            .I(n2695));
    CascadeMux I__2458 (
            .O(N__23589),
            .I(N__23586));
    InMux I__2457 (
            .O(N__23586),
            .I(N__23583));
    LocalMux I__2456 (
            .O(N__23583),
            .I(N__23579));
    CascadeMux I__2455 (
            .O(N__23582),
            .I(N__23576));
    Span4Mux_s3_h I__2454 (
            .O(N__23579),
            .I(N__23573));
    InMux I__2453 (
            .O(N__23576),
            .I(N__23570));
    Span4Mux_v I__2452 (
            .O(N__23573),
            .I(N__23567));
    LocalMux I__2451 (
            .O(N__23570),
            .I(n2628));
    Odrv4 I__2450 (
            .O(N__23567),
            .I(n2628));
    CascadeMux I__2449 (
            .O(N__23562),
            .I(N__23559));
    InMux I__2448 (
            .O(N__23559),
            .I(N__23556));
    LocalMux I__2447 (
            .O(N__23556),
            .I(N__23553));
    Span4Mux_v I__2446 (
            .O(N__23553),
            .I(N__23548));
    InMux I__2445 (
            .O(N__23552),
            .I(N__23543));
    InMux I__2444 (
            .O(N__23551),
            .I(N__23543));
    Odrv4 I__2443 (
            .O(N__23548),
            .I(n2727));
    LocalMux I__2442 (
            .O(N__23543),
            .I(n2727));
    InMux I__2441 (
            .O(N__23538),
            .I(N__23535));
    LocalMux I__2440 (
            .O(N__23535),
            .I(N__23532));
    Span4Mux_v I__2439 (
            .O(N__23532),
            .I(N__23529));
    Span4Mux_v I__2438 (
            .O(N__23529),
            .I(N__23526));
    Odrv4 I__2437 (
            .O(N__23526),
            .I(n2700));
    InMux I__2436 (
            .O(N__23523),
            .I(N__23520));
    LocalMux I__2435 (
            .O(N__23520),
            .I(N__23517));
    Odrv12 I__2434 (
            .O(N__23517),
            .I(n2288));
    InMux I__2433 (
            .O(N__23514),
            .I(N__23511));
    LocalMux I__2432 (
            .O(N__23511),
            .I(N__23508));
    Odrv4 I__2431 (
            .O(N__23508),
            .I(n2391));
    InMux I__2430 (
            .O(N__23505),
            .I(N__23502));
    LocalMux I__2429 (
            .O(N__23502),
            .I(N__23499));
    Odrv12 I__2428 (
            .O(N__23499),
            .I(n2287));
    InMux I__2427 (
            .O(N__23496),
            .I(N__23493));
    LocalMux I__2426 (
            .O(N__23493),
            .I(N__23490));
    Odrv4 I__2425 (
            .O(N__23490),
            .I(n2386));
    CascadeMux I__2424 (
            .O(N__23487),
            .I(n2319_cascade_));
    InMux I__2423 (
            .O(N__23484),
            .I(N__23481));
    LocalMux I__2422 (
            .O(N__23481),
            .I(N__23478));
    Odrv4 I__2421 (
            .O(N__23478),
            .I(n11971));
    InMux I__2420 (
            .O(N__23475),
            .I(N__23472));
    LocalMux I__2419 (
            .O(N__23472),
            .I(N__23469));
    Span4Mux_v I__2418 (
            .O(N__23469),
            .I(N__23466));
    Odrv4 I__2417 (
            .O(N__23466),
            .I(n2292));
    CascadeMux I__2416 (
            .O(N__23463),
            .I(N__23459));
    CascadeMux I__2415 (
            .O(N__23462),
            .I(N__23456));
    InMux I__2414 (
            .O(N__23459),
            .I(N__23453));
    InMux I__2413 (
            .O(N__23456),
            .I(N__23450));
    LocalMux I__2412 (
            .O(N__23453),
            .I(N__23447));
    LocalMux I__2411 (
            .O(N__23450),
            .I(n2324));
    Odrv4 I__2410 (
            .O(N__23447),
            .I(n2324));
    CascadeMux I__2409 (
            .O(N__23442),
            .I(n2324_cascade_));
    InMux I__2408 (
            .O(N__23439),
            .I(N__23436));
    LocalMux I__2407 (
            .O(N__23436),
            .I(N__23432));
    InMux I__2406 (
            .O(N__23435),
            .I(N__23429));
    Odrv4 I__2405 (
            .O(N__23432),
            .I(n2319));
    LocalMux I__2404 (
            .O(N__23429),
            .I(n2319));
    CascadeMux I__2403 (
            .O(N__23424),
            .I(n14384_cascade_));
    InMux I__2402 (
            .O(N__23421),
            .I(N__23418));
    LocalMux I__2401 (
            .O(N__23418),
            .I(N__23415));
    Odrv4 I__2400 (
            .O(N__23415),
            .I(n14382));
    InMux I__2399 (
            .O(N__23412),
            .I(N__23409));
    LocalMux I__2398 (
            .O(N__23409),
            .I(n14390));
    InMux I__2397 (
            .O(N__23406),
            .I(N__23403));
    LocalMux I__2396 (
            .O(N__23403),
            .I(N__23400));
    Odrv12 I__2395 (
            .O(N__23400),
            .I(n2293));
    InMux I__2394 (
            .O(N__23397),
            .I(N__23394));
    LocalMux I__2393 (
            .O(N__23394),
            .I(N__23391));
    Odrv12 I__2392 (
            .O(N__23391),
            .I(n2298));
    InMux I__2391 (
            .O(N__23388),
            .I(N__23385));
    LocalMux I__2390 (
            .O(N__23385),
            .I(N__23382));
    Odrv12 I__2389 (
            .O(N__23382),
            .I(n2295));
    InMux I__2388 (
            .O(N__23379),
            .I(N__23376));
    LocalMux I__2387 (
            .O(N__23376),
            .I(N__23373));
    Odrv12 I__2386 (
            .O(N__23373),
            .I(n2296));
    InMux I__2385 (
            .O(N__23370),
            .I(N__23367));
    LocalMux I__2384 (
            .O(N__23367),
            .I(N__23364));
    Odrv4 I__2383 (
            .O(N__23364),
            .I(n11977));
    CascadeMux I__2382 (
            .O(N__23361),
            .I(n14808_cascade_));
    InMux I__2381 (
            .O(N__23358),
            .I(N__23355));
    LocalMux I__2380 (
            .O(N__23355),
            .I(N__23352));
    Odrv4 I__2379 (
            .O(N__23352),
            .I(n14594));
    CascadeMux I__2378 (
            .O(N__23349),
            .I(N__23346));
    InMux I__2377 (
            .O(N__23346),
            .I(N__23343));
    LocalMux I__2376 (
            .O(N__23343),
            .I(N__23339));
    InMux I__2375 (
            .O(N__23342),
            .I(N__23336));
    Odrv4 I__2374 (
            .O(N__23339),
            .I(n2219));
    LocalMux I__2373 (
            .O(N__23336),
            .I(n2219));
    CascadeMux I__2372 (
            .O(N__23331),
            .I(n14598_cascade_));
    CascadeMux I__2371 (
            .O(N__23328),
            .I(n14604_cascade_));
    CascadeMux I__2370 (
            .O(N__23325),
            .I(n2247_cascade_));
    InMux I__2369 (
            .O(N__23322),
            .I(N__23319));
    LocalMux I__2368 (
            .O(N__23319),
            .I(N__23316));
    Span4Mux_v I__2367 (
            .O(N__23316),
            .I(N__23313));
    Odrv4 I__2366 (
            .O(N__23313),
            .I(n2297));
    CascadeMux I__2365 (
            .O(N__23310),
            .I(N__23307));
    InMux I__2364 (
            .O(N__23307),
            .I(N__23304));
    LocalMux I__2363 (
            .O(N__23304),
            .I(N__23300));
    InMux I__2362 (
            .O(N__23303),
            .I(N__23297));
    Odrv4 I__2361 (
            .O(N__23300),
            .I(n2222));
    LocalMux I__2360 (
            .O(N__23297),
            .I(n2222));
    CascadeMux I__2359 (
            .O(N__23292),
            .I(n2222_cascade_));
    InMux I__2358 (
            .O(N__23289),
            .I(N__23286));
    LocalMux I__2357 (
            .O(N__23286),
            .I(N__23283));
    Odrv4 I__2356 (
            .O(N__23283),
            .I(n2289));
    InMux I__2355 (
            .O(N__23280),
            .I(N__23277));
    LocalMux I__2354 (
            .O(N__23277),
            .I(N__23274));
    Odrv4 I__2353 (
            .O(N__23274),
            .I(n2291));
    CascadeMux I__2352 (
            .O(N__23271),
            .I(n2323_cascade_));
    CascadeMux I__2351 (
            .O(N__23268),
            .I(n2219_cascade_));
    InMux I__2350 (
            .O(N__23265),
            .I(N__23262));
    LocalMux I__2349 (
            .O(N__23262),
            .I(N__23259));
    Odrv12 I__2348 (
            .O(N__23259),
            .I(n2286));
    InMux I__2347 (
            .O(N__23256),
            .I(N__23253));
    LocalMux I__2346 (
            .O(N__23253),
            .I(N__23250));
    Odrv4 I__2345 (
            .O(N__23250),
            .I(n2290));
    InMux I__2344 (
            .O(N__23247),
            .I(n12693));
    InMux I__2343 (
            .O(N__23244),
            .I(n12694));
    InMux I__2342 (
            .O(N__23241),
            .I(n12695));
    CascadeMux I__2341 (
            .O(N__23238),
            .I(N__23235));
    InMux I__2340 (
            .O(N__23235),
            .I(N__23231));
    CascadeMux I__2339 (
            .O(N__23234),
            .I(N__23228));
    LocalMux I__2338 (
            .O(N__23231),
            .I(N__23225));
    InMux I__2337 (
            .O(N__23228),
            .I(N__23222));
    Odrv4 I__2336 (
            .O(N__23225),
            .I(n2233));
    LocalMux I__2335 (
            .O(N__23222),
            .I(n2233));
    InMux I__2334 (
            .O(N__23217),
            .I(N__23214));
    LocalMux I__2333 (
            .O(N__23214),
            .I(N__23211));
    Odrv12 I__2332 (
            .O(N__23211),
            .I(n2300));
    CascadeMux I__2331 (
            .O(N__23208),
            .I(n2233_cascade_));
    InMux I__2330 (
            .O(N__23205),
            .I(N__23202));
    LocalMux I__2329 (
            .O(N__23202),
            .I(N__23199));
    Odrv4 I__2328 (
            .O(N__23199),
            .I(n2299));
    CascadeMux I__2327 (
            .O(N__23196),
            .I(n2331_cascade_));
    InMux I__2326 (
            .O(N__23193),
            .I(N__23190));
    LocalMux I__2325 (
            .O(N__23190),
            .I(N__23187));
    Odrv12 I__2324 (
            .O(N__23187),
            .I(n2301));
    InMux I__2323 (
            .O(N__23184),
            .I(n12684));
    InMux I__2322 (
            .O(N__23181),
            .I(n12685));
    InMux I__2321 (
            .O(N__23178),
            .I(n12686));
    InMux I__2320 (
            .O(N__23175),
            .I(n12687));
    InMux I__2319 (
            .O(N__23172),
            .I(n12688));
    InMux I__2318 (
            .O(N__23169),
            .I(n12689));
    InMux I__2317 (
            .O(N__23166),
            .I(n12690));
    InMux I__2316 (
            .O(N__23163),
            .I(bfn_3_16_0_));
    InMux I__2315 (
            .O(N__23160),
            .I(n12692));
    InMux I__2314 (
            .O(N__23157),
            .I(bfn_3_14_0_));
    InMux I__2313 (
            .O(N__23154),
            .I(n12676));
    InMux I__2312 (
            .O(N__23151),
            .I(n12677));
    InMux I__2311 (
            .O(N__23148),
            .I(n12678));
    InMux I__2310 (
            .O(N__23145),
            .I(n12679));
    InMux I__2309 (
            .O(N__23142),
            .I(n12680));
    InMux I__2308 (
            .O(N__23139),
            .I(n12681));
    InMux I__2307 (
            .O(N__23136),
            .I(n12682));
    InMux I__2306 (
            .O(N__23133),
            .I(bfn_3_15_0_));
    InMux I__2305 (
            .O(N__23130),
            .I(n12912));
    InMux I__2304 (
            .O(N__23127),
            .I(n12913));
    InMux I__2303 (
            .O(N__23124),
            .I(n12914));
    InMux I__2302 (
            .O(N__23121),
            .I(bfn_2_32_0_));
    InMux I__2301 (
            .O(N__23118),
            .I(n12916));
    InMux I__2300 (
            .O(N__23115),
            .I(n12917));
    InMux I__2299 (
            .O(N__23112),
            .I(n12918));
    InMux I__2298 (
            .O(N__23109),
            .I(n12919));
    InMux I__2297 (
            .O(N__23106),
            .I(n12920));
    InMux I__2296 (
            .O(N__23103),
            .I(n12903));
    InMux I__2295 (
            .O(N__23100),
            .I(n12904));
    InMux I__2294 (
            .O(N__23097),
            .I(N__23093));
    InMux I__2293 (
            .O(N__23096),
            .I(N__23090));
    LocalMux I__2292 (
            .O(N__23093),
            .I(n3120));
    LocalMux I__2291 (
            .O(N__23090),
            .I(n3120));
    InMux I__2290 (
            .O(N__23085),
            .I(N__23082));
    LocalMux I__2289 (
            .O(N__23082),
            .I(n3187));
    InMux I__2288 (
            .O(N__23079),
            .I(n12905));
    InMux I__2287 (
            .O(N__23076),
            .I(n12906));
    InMux I__2286 (
            .O(N__23073),
            .I(bfn_2_31_0_));
    InMux I__2285 (
            .O(N__23070),
            .I(n12908));
    InMux I__2284 (
            .O(N__23067),
            .I(n12909));
    InMux I__2283 (
            .O(N__23064),
            .I(n12910));
    InMux I__2282 (
            .O(N__23061),
            .I(n12911));
    InMux I__2281 (
            .O(N__23058),
            .I(n12894));
    InMux I__2280 (
            .O(N__23055),
            .I(n12895));
    InMux I__2279 (
            .O(N__23052),
            .I(n12896));
    InMux I__2278 (
            .O(N__23049),
            .I(n12897));
    InMux I__2277 (
            .O(N__23046),
            .I(n12898));
    InMux I__2276 (
            .O(N__23043),
            .I(bfn_2_30_0_));
    InMux I__2275 (
            .O(N__23040),
            .I(n12900));
    InMux I__2274 (
            .O(N__23037),
            .I(n12901));
    InMux I__2273 (
            .O(N__23034),
            .I(n12902));
    InMux I__2272 (
            .O(N__23031),
            .I(n12861));
    InMux I__2271 (
            .O(N__23028),
            .I(N__23025));
    LocalMux I__2270 (
            .O(N__23025),
            .I(N__23022));
    Odrv4 I__2269 (
            .O(N__23022),
            .I(n2975));
    InMux I__2268 (
            .O(N__23019),
            .I(n12862));
    InMux I__2267 (
            .O(N__23016),
            .I(n12863));
    InMux I__2266 (
            .O(N__23013),
            .I(bfn_2_29_0_));
    InMux I__2265 (
            .O(N__23010),
            .I(n12892));
    InMux I__2264 (
            .O(N__23007),
            .I(n12893));
    InMux I__2263 (
            .O(N__23004),
            .I(N__23001));
    LocalMux I__2262 (
            .O(N__23001),
            .I(n2985));
    InMux I__2261 (
            .O(N__22998),
            .I(bfn_2_27_0_));
    InMux I__2260 (
            .O(N__22995),
            .I(n12853));
    InMux I__2259 (
            .O(N__22992),
            .I(n12854));
    InMux I__2258 (
            .O(N__22989),
            .I(n12855));
    InMux I__2257 (
            .O(N__22986),
            .I(n12856));
    InMux I__2256 (
            .O(N__22983),
            .I(n12857));
    InMux I__2255 (
            .O(N__22980),
            .I(n12858));
    InMux I__2254 (
            .O(N__22977),
            .I(n12859));
    CascadeMux I__2253 (
            .O(N__22974),
            .I(N__22971));
    InMux I__2252 (
            .O(N__22971),
            .I(N__22968));
    LocalMux I__2251 (
            .O(N__22968),
            .I(n2977));
    InMux I__2250 (
            .O(N__22965),
            .I(bfn_2_28_0_));
    InMux I__2249 (
            .O(N__22962),
            .I(N__22959));
    LocalMux I__2248 (
            .O(N__22959),
            .I(n2993));
    InMux I__2247 (
            .O(N__22956),
            .I(bfn_2_26_0_));
    InMux I__2246 (
            .O(N__22953),
            .I(N__22950));
    LocalMux I__2245 (
            .O(N__22950),
            .I(n2992));
    InMux I__2244 (
            .O(N__22947),
            .I(n12845));
    InMux I__2243 (
            .O(N__22944),
            .I(n12846));
    CascadeMux I__2242 (
            .O(N__22941),
            .I(N__22938));
    InMux I__2241 (
            .O(N__22938),
            .I(N__22935));
    LocalMux I__2240 (
            .O(N__22935),
            .I(n2990));
    InMux I__2239 (
            .O(N__22932),
            .I(n12847));
    InMux I__2238 (
            .O(N__22929),
            .I(N__22926));
    LocalMux I__2237 (
            .O(N__22926),
            .I(n2989));
    InMux I__2236 (
            .O(N__22923),
            .I(n12848));
    InMux I__2235 (
            .O(N__22920),
            .I(n12849));
    InMux I__2234 (
            .O(N__22917),
            .I(n12850));
    InMux I__2233 (
            .O(N__22914),
            .I(n12851));
    InMux I__2232 (
            .O(N__22911),
            .I(N__22908));
    LocalMux I__2231 (
            .O(N__22908),
            .I(N__22905));
    Odrv12 I__2230 (
            .O(N__22905),
            .I(n2791));
    InMux I__2229 (
            .O(N__22902),
            .I(bfn_2_25_0_));
    InMux I__2228 (
            .O(N__22899),
            .I(n12837));
    InMux I__2227 (
            .O(N__22896),
            .I(n12838));
    InMux I__2226 (
            .O(N__22893),
            .I(n12839));
    InMux I__2225 (
            .O(N__22890),
            .I(n12840));
    InMux I__2224 (
            .O(N__22887),
            .I(n12841));
    InMux I__2223 (
            .O(N__22884),
            .I(n12842));
    InMux I__2222 (
            .O(N__22881),
            .I(N__22878));
    LocalMux I__2221 (
            .O(N__22878),
            .I(n2994));
    InMux I__2220 (
            .O(N__22875),
            .I(n12843));
    InMux I__2219 (
            .O(N__22872),
            .I(N__22869));
    LocalMux I__2218 (
            .O(N__22869),
            .I(N__22866));
    Span4Mux_v I__2217 (
            .O(N__22866),
            .I(N__22863));
    Odrv4 I__2216 (
            .O(N__22863),
            .I(n2785));
    InMux I__2215 (
            .O(N__22860),
            .I(N__22857));
    LocalMux I__2214 (
            .O(N__22857),
            .I(N__22854));
    Span4Mux_v I__2213 (
            .O(N__22854),
            .I(N__22851));
    Span4Mux_v I__2212 (
            .O(N__22851),
            .I(N__22848));
    Odrv4 I__2211 (
            .O(N__22848),
            .I(n2684));
    InMux I__2210 (
            .O(N__22845),
            .I(N__22840));
    InMux I__2209 (
            .O(N__22844),
            .I(N__22837));
    CascadeMux I__2208 (
            .O(N__22843),
            .I(N__22834));
    LocalMux I__2207 (
            .O(N__22840),
            .I(N__22831));
    LocalMux I__2206 (
            .O(N__22837),
            .I(N__22828));
    InMux I__2205 (
            .O(N__22834),
            .I(N__22825));
    Odrv4 I__2204 (
            .O(N__22831),
            .I(n2716));
    Odrv12 I__2203 (
            .O(N__22828),
            .I(n2716));
    LocalMux I__2202 (
            .O(N__22825),
            .I(n2716));
    CascadeMux I__2201 (
            .O(N__22818),
            .I(N__22815));
    InMux I__2200 (
            .O(N__22815),
            .I(N__22812));
    LocalMux I__2199 (
            .O(N__22812),
            .I(N__22809));
    Span4Mux_v I__2198 (
            .O(N__22809),
            .I(N__22806));
    Span4Mux_v I__2197 (
            .O(N__22806),
            .I(N__22803));
    Odrv4 I__2196 (
            .O(N__22803),
            .I(n2679));
    InMux I__2195 (
            .O(N__22800),
            .I(N__22796));
    InMux I__2194 (
            .O(N__22799),
            .I(N__22793));
    LocalMux I__2193 (
            .O(N__22796),
            .I(N__22790));
    LocalMux I__2192 (
            .O(N__22793),
            .I(n2709));
    Odrv12 I__2191 (
            .O(N__22790),
            .I(n2709));
    CascadeMux I__2190 (
            .O(N__22785),
            .I(n2711_cascade_));
    InMux I__2189 (
            .O(N__22782),
            .I(N__22779));
    LocalMux I__2188 (
            .O(N__22779),
            .I(n14368));
    InMux I__2187 (
            .O(N__22776),
            .I(N__22773));
    LocalMux I__2186 (
            .O(N__22773),
            .I(N__22770));
    Span4Mux_v I__2185 (
            .O(N__22770),
            .I(N__22767));
    Odrv4 I__2184 (
            .O(N__22767),
            .I(n2796));
    CascadeMux I__2183 (
            .O(N__22764),
            .I(n2742_cascade_));
    CascadeMux I__2182 (
            .O(N__22761),
            .I(N__22758));
    InMux I__2181 (
            .O(N__22758),
            .I(N__22753));
    InMux I__2180 (
            .O(N__22757),
            .I(N__22750));
    InMux I__2179 (
            .O(N__22756),
            .I(N__22747));
    LocalMux I__2178 (
            .O(N__22753),
            .I(N__22744));
    LocalMux I__2177 (
            .O(N__22750),
            .I(N__22741));
    LocalMux I__2176 (
            .O(N__22747),
            .I(N__22738));
    Odrv4 I__2175 (
            .O(N__22744),
            .I(n2828));
    Odrv4 I__2174 (
            .O(N__22741),
            .I(n2828));
    Odrv4 I__2173 (
            .O(N__22738),
            .I(n2828));
    InMux I__2172 (
            .O(N__22731),
            .I(N__22728));
    LocalMux I__2171 (
            .O(N__22728),
            .I(N__22725));
    Span4Mux_v I__2170 (
            .O(N__22725),
            .I(N__22722));
    Odrv4 I__2169 (
            .O(N__22722),
            .I(n2788));
    InMux I__2168 (
            .O(N__22719),
            .I(N__22716));
    LocalMux I__2167 (
            .O(N__22716),
            .I(N__22713));
    Span12Mux_v I__2166 (
            .O(N__22713),
            .I(N__22710));
    Odrv12 I__2165 (
            .O(N__22710),
            .I(n2687));
    InMux I__2164 (
            .O(N__22707),
            .I(N__22704));
    LocalMux I__2163 (
            .O(N__22704),
            .I(N__22701));
    Odrv12 I__2162 (
            .O(N__22701),
            .I(n2792));
    CascadeMux I__2161 (
            .O(N__22698),
            .I(N__22695));
    InMux I__2160 (
            .O(N__22695),
            .I(N__22691));
    InMux I__2159 (
            .O(N__22694),
            .I(N__22687));
    LocalMux I__2158 (
            .O(N__22691),
            .I(N__22684));
    CascadeMux I__2157 (
            .O(N__22690),
            .I(N__22681));
    LocalMux I__2156 (
            .O(N__22687),
            .I(N__22678));
    Span4Mux_s2_h I__2155 (
            .O(N__22684),
            .I(N__22675));
    InMux I__2154 (
            .O(N__22681),
            .I(N__22672));
    Odrv4 I__2153 (
            .O(N__22678),
            .I(n2725));
    Odrv4 I__2152 (
            .O(N__22675),
            .I(n2725));
    LocalMux I__2151 (
            .O(N__22672),
            .I(n2725));
    CascadeMux I__2150 (
            .O(N__22665),
            .I(N__22662));
    InMux I__2149 (
            .O(N__22662),
            .I(N__22659));
    LocalMux I__2148 (
            .O(N__22659),
            .I(N__22656));
    Span4Mux_v I__2147 (
            .O(N__22656),
            .I(N__22653));
    Odrv4 I__2146 (
            .O(N__22653),
            .I(n2681));
    CascadeMux I__2145 (
            .O(N__22650),
            .I(N__22647));
    InMux I__2144 (
            .O(N__22647),
            .I(N__22644));
    LocalMux I__2143 (
            .O(N__22644),
            .I(N__22641));
    Span4Mux_v I__2142 (
            .O(N__22641),
            .I(N__22638));
    Odrv4 I__2141 (
            .O(N__22638),
            .I(n2794));
    CascadeMux I__2140 (
            .O(N__22635),
            .I(n2826_cascade_));
    CascadeMux I__2139 (
            .O(N__22632),
            .I(n14362_cascade_));
    InMux I__2138 (
            .O(N__22629),
            .I(N__22626));
    LocalMux I__2137 (
            .O(N__22626),
            .I(N__22623));
    Span4Mux_v I__2136 (
            .O(N__22623),
            .I(N__22620));
    Odrv4 I__2135 (
            .O(N__22620),
            .I(n2789));
    CascadeMux I__2134 (
            .O(N__22617),
            .I(N__22614));
    InMux I__2133 (
            .O(N__22614),
            .I(N__22611));
    LocalMux I__2132 (
            .O(N__22611),
            .I(n14346));
    CascadeMux I__2131 (
            .O(N__22608),
            .I(n14350_cascade_));
    InMux I__2130 (
            .O(N__22605),
            .I(N__22602));
    LocalMux I__2129 (
            .O(N__22602),
            .I(n14356));
    InMux I__2128 (
            .O(N__22599),
            .I(N__22596));
    LocalMux I__2127 (
            .O(N__22596),
            .I(N__22593));
    Span4Mux_v I__2126 (
            .O(N__22593),
            .I(N__22590));
    Odrv4 I__2125 (
            .O(N__22590),
            .I(n2782));
    CascadeMux I__2124 (
            .O(N__22587),
            .I(N__22584));
    InMux I__2123 (
            .O(N__22584),
            .I(N__22577));
    InMux I__2122 (
            .O(N__22583),
            .I(N__22577));
    InMux I__2121 (
            .O(N__22582),
            .I(N__22574));
    LocalMux I__2120 (
            .O(N__22577),
            .I(N__22571));
    LocalMux I__2119 (
            .O(N__22574),
            .I(n2715));
    Odrv4 I__2118 (
            .O(N__22571),
            .I(n2715));
    CascadeMux I__2117 (
            .O(N__22566),
            .I(n2621_cascade_));
    InMux I__2116 (
            .O(N__22563),
            .I(N__22560));
    LocalMux I__2115 (
            .O(N__22560),
            .I(N__22557));
    Span4Mux_v I__2114 (
            .O(N__22557),
            .I(N__22554));
    Odrv4 I__2113 (
            .O(N__22554),
            .I(n2688));
    InMux I__2112 (
            .O(N__22551),
            .I(N__22548));
    LocalMux I__2111 (
            .O(N__22548),
            .I(N__22545));
    Span4Mux_v I__2110 (
            .O(N__22545),
            .I(N__22542));
    Span4Mux_v I__2109 (
            .O(N__22542),
            .I(N__22539));
    Odrv4 I__2108 (
            .O(N__22539),
            .I(n2696));
    InMux I__2107 (
            .O(N__22536),
            .I(N__22533));
    LocalMux I__2106 (
            .O(N__22533),
            .I(N__22530));
    Odrv12 I__2105 (
            .O(N__22530),
            .I(n2795));
    CascadeMux I__2104 (
            .O(N__22527),
            .I(n2728_cascade_));
    CascadeMux I__2103 (
            .O(N__22524),
            .I(N__22521));
    InMux I__2102 (
            .O(N__22521),
            .I(N__22518));
    LocalMux I__2101 (
            .O(N__22518),
            .I(N__22515));
    Odrv12 I__2100 (
            .O(N__22515),
            .I(n2691));
    CascadeMux I__2099 (
            .O(N__22512),
            .I(N__22509));
    InMux I__2098 (
            .O(N__22509),
            .I(N__22506));
    LocalMux I__2097 (
            .O(N__22506),
            .I(N__22503));
    Span4Mux_s2_h I__2096 (
            .O(N__22503),
            .I(N__22499));
    InMux I__2095 (
            .O(N__22502),
            .I(N__22496));
    Odrv4 I__2094 (
            .O(N__22499),
            .I(n2723));
    LocalMux I__2093 (
            .O(N__22496),
            .I(n2723));
    InMux I__2092 (
            .O(N__22491),
            .I(N__22488));
    LocalMux I__2091 (
            .O(N__22488),
            .I(N__22485));
    Span4Mux_v I__2090 (
            .O(N__22485),
            .I(N__22482));
    Odrv4 I__2089 (
            .O(N__22482),
            .I(n2790));
    CascadeMux I__2088 (
            .O(N__22479),
            .I(n2723_cascade_));
    InMux I__2087 (
            .O(N__22476),
            .I(N__22473));
    LocalMux I__2086 (
            .O(N__22473),
            .I(N__22470));
    Odrv12 I__2085 (
            .O(N__22470),
            .I(n2693));
    InMux I__2084 (
            .O(N__22467),
            .I(N__22464));
    LocalMux I__2083 (
            .O(N__22464),
            .I(N__22461));
    Span4Mux_v I__2082 (
            .O(N__22461),
            .I(N__22458));
    Span4Mux_v I__2081 (
            .O(N__22458),
            .I(N__22455));
    Odrv4 I__2080 (
            .O(N__22455),
            .I(n2697));
    InMux I__2079 (
            .O(N__22452),
            .I(bfn_2_20_0_));
    InMux I__2078 (
            .O(N__22449),
            .I(n12810));
    InMux I__2077 (
            .O(N__22446),
            .I(N__22443));
    LocalMux I__2076 (
            .O(N__22443),
            .I(N__22440));
    Odrv12 I__2075 (
            .O(N__22440),
            .I(n2683));
    CascadeMux I__2074 (
            .O(N__22437),
            .I(N__22434));
    InMux I__2073 (
            .O(N__22434),
            .I(N__22431));
    LocalMux I__2072 (
            .O(N__22431),
            .I(N__22428));
    Span4Mux_v I__2071 (
            .O(N__22428),
            .I(N__22425));
    Odrv4 I__2070 (
            .O(N__22425),
            .I(n2677));
    InMux I__2069 (
            .O(N__22422),
            .I(N__22419));
    LocalMux I__2068 (
            .O(N__22419),
            .I(N__22416));
    Odrv12 I__2067 (
            .O(N__22416),
            .I(n2678));
    InMux I__2066 (
            .O(N__22413),
            .I(N__22410));
    LocalMux I__2065 (
            .O(N__22410),
            .I(N__22407));
    Odrv12 I__2064 (
            .O(N__22407),
            .I(n2797));
    CascadeMux I__2063 (
            .O(N__22404),
            .I(N__22401));
    InMux I__2062 (
            .O(N__22401),
            .I(N__22398));
    LocalMux I__2061 (
            .O(N__22398),
            .I(N__22395));
    Sp12to4 I__2060 (
            .O(N__22395),
            .I(N__22392));
    Odrv12 I__2059 (
            .O(N__22392),
            .I(n2694));
    InMux I__2058 (
            .O(N__22389),
            .I(N__22386));
    LocalMux I__2057 (
            .O(N__22386),
            .I(N__22383));
    Span4Mux_v I__2056 (
            .O(N__22383),
            .I(N__22380));
    Odrv4 I__2055 (
            .O(N__22380),
            .I(n2793));
    CascadeMux I__2054 (
            .O(N__22377),
            .I(n2726_cascade_));
    InMux I__2053 (
            .O(N__22374),
            .I(n12800));
    InMux I__2052 (
            .O(N__22371),
            .I(bfn_2_19_0_));
    InMux I__2051 (
            .O(N__22368),
            .I(n12802));
    CascadeMux I__2050 (
            .O(N__22365),
            .I(N__22362));
    InMux I__2049 (
            .O(N__22362),
            .I(N__22359));
    LocalMux I__2048 (
            .O(N__22359),
            .I(N__22356));
    Sp12to4 I__2047 (
            .O(N__22356),
            .I(N__22353));
    Odrv12 I__2046 (
            .O(N__22353),
            .I(n2783));
    InMux I__2045 (
            .O(N__22350),
            .I(n12803));
    InMux I__2044 (
            .O(N__22347),
            .I(n12804));
    InMux I__2043 (
            .O(N__22344),
            .I(n12805));
    InMux I__2042 (
            .O(N__22341),
            .I(n12806));
    InMux I__2041 (
            .O(N__22338),
            .I(n12807));
    InMux I__2040 (
            .O(N__22335),
            .I(n12808));
    InMux I__2039 (
            .O(N__22332),
            .I(n12791));
    InMux I__2038 (
            .O(N__22329),
            .I(n12792));
    InMux I__2037 (
            .O(N__22326),
            .I(bfn_2_18_0_));
    InMux I__2036 (
            .O(N__22323),
            .I(n12794));
    InMux I__2035 (
            .O(N__22320),
            .I(n12795));
    InMux I__2034 (
            .O(N__22317),
            .I(n12796));
    InMux I__2033 (
            .O(N__22314),
            .I(n12797));
    InMux I__2032 (
            .O(N__22311),
            .I(n12798));
    InMux I__2031 (
            .O(N__22308),
            .I(n12799));
    InMux I__2030 (
            .O(N__22305),
            .I(n12783));
    InMux I__2029 (
            .O(N__22302),
            .I(n12784));
    InMux I__2028 (
            .O(N__22299),
            .I(bfn_2_16_0_));
    InMux I__2027 (
            .O(N__22296),
            .I(N__22293));
    LocalMux I__2026 (
            .O(N__22293),
            .I(N__22290));
    Span4Mux_v I__2025 (
            .O(N__22290),
            .I(N__22287));
    Span4Mux_v I__2024 (
            .O(N__22287),
            .I(N__22284));
    Odrv4 I__2023 (
            .O(N__22284),
            .I(n2801));
    InMux I__2022 (
            .O(N__22281),
            .I(bfn_2_17_0_));
    InMux I__2021 (
            .O(N__22278),
            .I(n12786));
    InMux I__2020 (
            .O(N__22275),
            .I(n12787));
    InMux I__2019 (
            .O(N__22272),
            .I(n12788));
    InMux I__2018 (
            .O(N__22269),
            .I(n12789));
    InMux I__2017 (
            .O(N__22266),
            .I(n12790));
    InMux I__2016 (
            .O(N__22263),
            .I(n12774));
    InMux I__2015 (
            .O(N__22260),
            .I(n12775));
    InMux I__2014 (
            .O(N__22257),
            .I(n12776));
    InMux I__2013 (
            .O(N__22254),
            .I(bfn_2_15_0_));
    InMux I__2012 (
            .O(N__22251),
            .I(n12778));
    InMux I__2011 (
            .O(N__22248),
            .I(n12779));
    InMux I__2010 (
            .O(N__22245),
            .I(N__22242));
    LocalMux I__2009 (
            .O(N__22242),
            .I(N__22239));
    Sp12to4 I__2008 (
            .O(N__22239),
            .I(N__22236));
    Odrv12 I__2007 (
            .O(N__22236),
            .I(n2682));
    InMux I__2006 (
            .O(N__22233),
            .I(n12780));
    InMux I__2005 (
            .O(N__22230),
            .I(n12781));
    InMux I__2004 (
            .O(N__22227),
            .I(n12782));
    InMux I__2003 (
            .O(N__22224),
            .I(n12764));
    InMux I__2002 (
            .O(N__22221),
            .I(n12765));
    InMux I__2001 (
            .O(N__22218),
            .I(n12766));
    InMux I__2000 (
            .O(N__22215),
            .I(n12767));
    InMux I__1999 (
            .O(N__22212),
            .I(n12768));
    InMux I__1998 (
            .O(N__22209),
            .I(bfn_2_14_0_));
    InMux I__1997 (
            .O(N__22206),
            .I(n12770));
    InMux I__1996 (
            .O(N__22203),
            .I(n12771));
    InMux I__1995 (
            .O(N__22200),
            .I(n12772));
    InMux I__1994 (
            .O(N__22197),
            .I(n12773));
    InMux I__1993 (
            .O(N__22194),
            .I(N__22190));
    InMux I__1992 (
            .O(N__22193),
            .I(N__22187));
    LocalMux I__1991 (
            .O(N__22190),
            .I(\debounce.cnt_reg_5 ));
    LocalMux I__1990 (
            .O(N__22187),
            .I(\debounce.cnt_reg_5 ));
    InMux I__1989 (
            .O(N__22182),
            .I(\debounce.n13017 ));
    InMux I__1988 (
            .O(N__22179),
            .I(N__22175));
    InMux I__1987 (
            .O(N__22178),
            .I(N__22172));
    LocalMux I__1986 (
            .O(N__22175),
            .I(\debounce.cnt_reg_6 ));
    LocalMux I__1985 (
            .O(N__22172),
            .I(\debounce.cnt_reg_6 ));
    InMux I__1984 (
            .O(N__22167),
            .I(\debounce.n13018 ));
    InMux I__1983 (
            .O(N__22164),
            .I(N__22160));
    InMux I__1982 (
            .O(N__22163),
            .I(N__22157));
    LocalMux I__1981 (
            .O(N__22160),
            .I(\debounce.cnt_reg_7 ));
    LocalMux I__1980 (
            .O(N__22157),
            .I(\debounce.cnt_reg_7 ));
    InMux I__1979 (
            .O(N__22152),
            .I(\debounce.n13019 ));
    InMux I__1978 (
            .O(N__22149),
            .I(N__22145));
    InMux I__1977 (
            .O(N__22148),
            .I(N__22142));
    LocalMux I__1976 (
            .O(N__22145),
            .I(N__22139));
    LocalMux I__1975 (
            .O(N__22142),
            .I(\debounce.cnt_reg_8 ));
    Odrv4 I__1974 (
            .O(N__22139),
            .I(\debounce.cnt_reg_8 ));
    InMux I__1973 (
            .O(N__22134),
            .I(bfn_1_32_0_));
    InMux I__1972 (
            .O(N__22131),
            .I(\debounce.n13021 ));
    CascadeMux I__1971 (
            .O(N__22128),
            .I(N__22125));
    InMux I__1970 (
            .O(N__22125),
            .I(N__22121));
    InMux I__1969 (
            .O(N__22124),
            .I(N__22118));
    LocalMux I__1968 (
            .O(N__22121),
            .I(N__22115));
    LocalMux I__1967 (
            .O(N__22118),
            .I(\debounce.cnt_reg_9 ));
    Odrv4 I__1966 (
            .O(N__22115),
            .I(\debounce.cnt_reg_9 ));
    SRMux I__1965 (
            .O(N__22110),
            .I(N__22107));
    LocalMux I__1964 (
            .O(N__22107),
            .I(N__22103));
    SRMux I__1963 (
            .O(N__22106),
            .I(N__22100));
    Span4Mux_s1_v I__1962 (
            .O(N__22103),
            .I(N__22097));
    LocalMux I__1961 (
            .O(N__22100),
            .I(N__22094));
    Odrv4 I__1960 (
            .O(N__22097),
            .I(\debounce.cnt_next_9__N_424 ));
    Odrv12 I__1959 (
            .O(N__22094),
            .I(\debounce.cnt_next_9__N_424 ));
    InMux I__1958 (
            .O(N__22089),
            .I(bfn_2_13_0_));
    InMux I__1957 (
            .O(N__22086),
            .I(n12762));
    InMux I__1956 (
            .O(N__22083),
            .I(n12763));
    CascadeMux I__1955 (
            .O(N__22080),
            .I(\debounce.n16_cascade_ ));
    InMux I__1954 (
            .O(N__22077),
            .I(N__22074));
    LocalMux I__1953 (
            .O(N__22074),
            .I(\debounce.n17 ));
    InMux I__1952 (
            .O(N__22071),
            .I(N__22065));
    InMux I__1951 (
            .O(N__22070),
            .I(N__22065));
    LocalMux I__1950 (
            .O(N__22065),
            .I(reg_B_2));
    CascadeMux I__1949 (
            .O(N__22062),
            .I(n14129_cascade_));
    InMux I__1948 (
            .O(N__22059),
            .I(N__22055));
    InMux I__1947 (
            .O(N__22058),
            .I(N__22052));
    LocalMux I__1946 (
            .O(N__22055),
            .I(\debounce.cnt_reg_0 ));
    LocalMux I__1945 (
            .O(N__22052),
            .I(\debounce.cnt_reg_0 ));
    InMux I__1944 (
            .O(N__22047),
            .I(bfn_1_31_0_));
    InMux I__1943 (
            .O(N__22044),
            .I(N__22040));
    InMux I__1942 (
            .O(N__22043),
            .I(N__22037));
    LocalMux I__1941 (
            .O(N__22040),
            .I(\debounce.cnt_reg_1 ));
    LocalMux I__1940 (
            .O(N__22037),
            .I(\debounce.cnt_reg_1 ));
    InMux I__1939 (
            .O(N__22032),
            .I(\debounce.n13013 ));
    CascadeMux I__1938 (
            .O(N__22029),
            .I(N__22025));
    InMux I__1937 (
            .O(N__22028),
            .I(N__22022));
    InMux I__1936 (
            .O(N__22025),
            .I(N__22019));
    LocalMux I__1935 (
            .O(N__22022),
            .I(\debounce.cnt_reg_2 ));
    LocalMux I__1934 (
            .O(N__22019),
            .I(\debounce.cnt_reg_2 ));
    InMux I__1933 (
            .O(N__22014),
            .I(\debounce.n13014 ));
    InMux I__1932 (
            .O(N__22011),
            .I(N__22007));
    InMux I__1931 (
            .O(N__22010),
            .I(N__22004));
    LocalMux I__1930 (
            .O(N__22007),
            .I(\debounce.cnt_reg_3 ));
    LocalMux I__1929 (
            .O(N__22004),
            .I(\debounce.cnt_reg_3 ));
    InMux I__1928 (
            .O(N__21999),
            .I(\debounce.n13015 ));
    InMux I__1927 (
            .O(N__21996),
            .I(N__21992));
    InMux I__1926 (
            .O(N__21995),
            .I(N__21989));
    LocalMux I__1925 (
            .O(N__21992),
            .I(\debounce.cnt_reg_4 ));
    LocalMux I__1924 (
            .O(N__21989),
            .I(\debounce.cnt_reg_4 ));
    InMux I__1923 (
            .O(N__21984),
            .I(\debounce.n13016 ));
    CascadeMux I__1922 (
            .O(N__21981),
            .I(n3120_cascade_));
    CascadeMux I__1921 (
            .O(N__21978),
            .I(n3122_cascade_));
    InMux I__1920 (
            .O(N__21975),
            .I(N__21972));
    LocalMux I__1919 (
            .O(N__21972),
            .I(n14146));
    InMux I__1918 (
            .O(N__21969),
            .I(N__21963));
    InMux I__1917 (
            .O(N__21968),
            .I(N__21963));
    LocalMux I__1916 (
            .O(N__21963),
            .I(\debounce.reg_A_2 ));
    CascadeMux I__1915 (
            .O(N__21960),
            .I(N__21956));
    InMux I__1914 (
            .O(N__21959),
            .I(N__21951));
    InMux I__1913 (
            .O(N__21956),
            .I(N__21951));
    LocalMux I__1912 (
            .O(N__21951),
            .I(N__21948));
    IoSpan4Mux I__1911 (
            .O(N__21948),
            .I(N__21945));
    Odrv4 I__1910 (
            .O(N__21945),
            .I(\debounce.reg_A_1 ));
    InMux I__1909 (
            .O(N__21942),
            .I(N__21938));
    InMux I__1908 (
            .O(N__21941),
            .I(N__21935));
    LocalMux I__1907 (
            .O(N__21938),
            .I(N__21932));
    LocalMux I__1906 (
            .O(N__21935),
            .I(N__21929));
    Span4Mux_h I__1905 (
            .O(N__21932),
            .I(N__21924));
    Span4Mux_v I__1904 (
            .O(N__21929),
            .I(N__21924));
    Odrv4 I__1903 (
            .O(N__21924),
            .I(\debounce.reg_A_0 ));
    InMux I__1902 (
            .O(N__21921),
            .I(N__21917));
    InMux I__1901 (
            .O(N__21920),
            .I(N__21914));
    LocalMux I__1900 (
            .O(N__21917),
            .I(N__21911));
    LocalMux I__1899 (
            .O(N__21914),
            .I(N__21908));
    Odrv4 I__1898 (
            .O(N__21911),
            .I(reg_B_0));
    Odrv12 I__1897 (
            .O(N__21908),
            .I(reg_B_0));
    CascadeMux I__1896 (
            .O(N__21903),
            .I(\debounce.n6_cascade_ ));
    CascadeMux I__1895 (
            .O(N__21900),
            .I(n3021_cascade_));
    InMux I__1894 (
            .O(N__21897),
            .I(N__21894));
    LocalMux I__1893 (
            .O(N__21894),
            .I(n14728));
    CascadeMux I__1892 (
            .O(N__21891),
            .I(n14150_cascade_));
    CascadeMux I__1891 (
            .O(N__21888),
            .I(n3128_cascade_));
    InMux I__1890 (
            .O(N__21885),
            .I(N__21882));
    LocalMux I__1889 (
            .O(N__21882),
            .I(n14148));
    InMux I__1888 (
            .O(N__21879),
            .I(N__21876));
    LocalMux I__1887 (
            .O(N__21876),
            .I(N__21873));
    Span4Mux_v I__1886 (
            .O(N__21873),
            .I(N__21870));
    Odrv4 I__1885 (
            .O(N__21870),
            .I(n2895));
    CascadeMux I__1884 (
            .O(N__21867),
            .I(n2927_cascade_));
    CascadeMux I__1883 (
            .O(N__21864),
            .I(n3024_cascade_));
    CascadeMux I__1882 (
            .O(N__21861),
            .I(n14730_cascade_));
    InMux I__1881 (
            .O(N__21858),
            .I(n12835));
    InMux I__1880 (
            .O(N__21855),
            .I(n12836));
    InMux I__1879 (
            .O(N__21852),
            .I(N__21849));
    LocalMux I__1878 (
            .O(N__21849),
            .I(n2882));
    CascadeMux I__1877 (
            .O(N__21846),
            .I(N__21843));
    InMux I__1876 (
            .O(N__21843),
            .I(N__21840));
    LocalMux I__1875 (
            .O(N__21840),
            .I(N__21837));
    Odrv12 I__1874 (
            .O(N__21837),
            .I(n2900));
    InMux I__1873 (
            .O(N__21834),
            .I(N__21831));
    LocalMux I__1872 (
            .O(N__21831),
            .I(n2876));
    CascadeMux I__1871 (
            .O(N__21828),
            .I(n2908_cascade_));
    InMux I__1870 (
            .O(N__21825),
            .I(bfn_1_24_0_));
    InMux I__1869 (
            .O(N__21822),
            .I(n12827));
    InMux I__1868 (
            .O(N__21819),
            .I(n12828));
    InMux I__1867 (
            .O(N__21816),
            .I(n12829));
    InMux I__1866 (
            .O(N__21813),
            .I(n12830));
    InMux I__1865 (
            .O(N__21810),
            .I(n12831));
    InMux I__1864 (
            .O(N__21807),
            .I(n12832));
    InMux I__1863 (
            .O(N__21804),
            .I(n12833));
    InMux I__1862 (
            .O(N__21801),
            .I(bfn_1_25_0_));
    InMux I__1861 (
            .O(N__21798),
            .I(n12817));
    InMux I__1860 (
            .O(N__21795),
            .I(bfn_1_23_0_));
    InMux I__1859 (
            .O(N__21792),
            .I(n12819));
    InMux I__1858 (
            .O(N__21789),
            .I(n12820));
    InMux I__1857 (
            .O(N__21786),
            .I(n12821));
    InMux I__1856 (
            .O(N__21783),
            .I(n12822));
    InMux I__1855 (
            .O(N__21780),
            .I(n12823));
    InMux I__1854 (
            .O(N__21777),
            .I(n12824));
    InMux I__1853 (
            .O(N__21774),
            .I(n12825));
    InMux I__1852 (
            .O(N__21771),
            .I(n12715));
    InMux I__1851 (
            .O(N__21768),
            .I(n12716));
    InMux I__1850 (
            .O(N__21765),
            .I(bfn_1_22_0_));
    InMux I__1849 (
            .O(N__21762),
            .I(n12811));
    InMux I__1848 (
            .O(N__21759),
            .I(n12812));
    InMux I__1847 (
            .O(N__21756),
            .I(n12813));
    InMux I__1846 (
            .O(N__21753),
            .I(n12814));
    InMux I__1845 (
            .O(N__21750),
            .I(n12815));
    InMux I__1844 (
            .O(N__21747),
            .I(n12816));
    InMux I__1843 (
            .O(N__21744),
            .I(n12706));
    InMux I__1842 (
            .O(N__21741),
            .I(n12707));
    InMux I__1841 (
            .O(N__21738),
            .I(n12708));
    InMux I__1840 (
            .O(N__21735),
            .I(n12709));
    InMux I__1839 (
            .O(N__21732),
            .I(n12710));
    InMux I__1838 (
            .O(N__21729),
            .I(bfn_1_21_0_));
    InMux I__1837 (
            .O(N__21726),
            .I(n12712));
    InMux I__1836 (
            .O(N__21723),
            .I(n12713));
    InMux I__1835 (
            .O(N__21720),
            .I(n12714));
    InMux I__1834 (
            .O(N__21717),
            .I(n12697));
    InMux I__1833 (
            .O(N__21714),
            .I(n12698));
    InMux I__1832 (
            .O(N__21711),
            .I(n12699));
    InMux I__1831 (
            .O(N__21708),
            .I(n12700));
    InMux I__1830 (
            .O(N__21705),
            .I(n12701));
    InMux I__1829 (
            .O(N__21702),
            .I(n12702));
    InMux I__1828 (
            .O(N__21699),
            .I(bfn_1_20_0_));
    InMux I__1827 (
            .O(N__21696),
            .I(n12704));
    InMux I__1826 (
            .O(N__21693),
            .I(n12705));
    InMux I__1825 (
            .O(N__21690),
            .I(bfn_1_19_0_));
    InMux I__1824 (
            .O(N__21687),
            .I(n12696));
    IoInMux I__1823 (
            .O(N__21684),
            .I(N__21681));
    LocalMux I__1822 (
            .O(N__21681),
            .I(N__21678));
    IoSpan4Mux I__1821 (
            .O(N__21678),
            .I(N__21675));
    IoSpan4Mux I__1820 (
            .O(N__21675),
            .I(N__21672));
    IoSpan4Mux I__1819 (
            .O(N__21672),
            .I(N__21669));
    Odrv4 I__1818 (
            .O(N__21669),
            .I(CLK_pad_gb_input));
    defparam IN_MUX_bfv_7_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_29_0_));
    defparam IN_MUX_bfv_7_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_30_0_ (
            .carryinitin(n12928),
            .carryinitout(bfn_7_30_0_));
    defparam IN_MUX_bfv_7_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_31_0_ (
            .carryinitin(n12936),
            .carryinitout(bfn_7_31_0_));
    defparam IN_MUX_bfv_7_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_32_0_ (
            .carryinitin(n12944),
            .carryinitout(bfn_7_32_0_));
    defparam IN_MUX_bfv_15_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_25_0_));
    defparam IN_MUX_bfv_15_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_26_0_ (
            .carryinitin(n12456),
            .carryinitout(bfn_15_26_0_));
    defparam IN_MUX_bfv_15_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_27_0_ (
            .carryinitin(n12464),
            .carryinitout(bfn_15_27_0_));
    defparam IN_MUX_bfv_15_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_28_0_ (
            .carryinitin(n12472),
            .carryinitout(bfn_15_28_0_));
    defparam IN_MUX_bfv_11_26_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_26_0_));
    defparam IN_MUX_bfv_11_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_27_0_ (
            .carryinitin(n12433),
            .carryinitout(bfn_11_27_0_));
    defparam IN_MUX_bfv_11_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_28_0_ (
            .carryinitin(n12441),
            .carryinitout(bfn_11_28_0_));
    defparam IN_MUX_bfv_16_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_25_0_));
    defparam IN_MUX_bfv_16_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_26_0_ (
            .carryinitin(n13060),
            .carryinitout(bfn_16_26_0_));
    defparam IN_MUX_bfv_16_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_27_0_ (
            .carryinitin(n13068),
            .carryinitout(bfn_16_27_0_));
    defparam IN_MUX_bfv_10_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_18_0_));
    defparam IN_MUX_bfv_10_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_19_0_ (
            .carryinitin(\quad_counter0.n13102 ),
            .carryinitout(bfn_10_19_0_));
    defparam IN_MUX_bfv_10_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_20_0_ (
            .carryinitin(\quad_counter0.n13110 ),
            .carryinitout(bfn_10_20_0_));
    defparam IN_MUX_bfv_10_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_21_0_ (
            .carryinitin(\quad_counter0.n13118 ),
            .carryinitout(bfn_10_21_0_));
    defparam IN_MUX_bfv_12_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_25_0_));
    defparam IN_MUX_bfv_12_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_26_0_ (
            .carryinitin(n12480),
            .carryinitout(bfn_12_26_0_));
    defparam IN_MUX_bfv_12_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_27_0_ (
            .carryinitin(n12488),
            .carryinitout(bfn_12_27_0_));
    defparam IN_MUX_bfv_9_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_22_0_));
    defparam IN_MUX_bfv_9_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_23_0_ (
            .carryinitin(n12982),
            .carryinitout(bfn_9_23_0_));
    defparam IN_MUX_bfv_9_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_24_0_ (
            .carryinitin(n12990),
            .carryinitout(bfn_9_24_0_));
    defparam IN_MUX_bfv_9_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_25_0_ (
            .carryinitin(n12998),
            .carryinitout(bfn_9_25_0_));
    defparam IN_MUX_bfv_16_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_17_0_));
    defparam IN_MUX_bfv_16_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_18_0_ (
            .carryinitin(n12559),
            .carryinitout(bfn_16_18_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(n12548),
            .carryinitout(bfn_14_21_0_));
    defparam IN_MUX_bfv_16_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_21_0_));
    defparam IN_MUX_bfv_16_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_22_0_ (
            .carryinitin(n12538),
            .carryinitout(bfn_16_22_0_));
    defparam IN_MUX_bfv_14_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_23_0_));
    defparam IN_MUX_bfv_14_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_24_0_ (
            .carryinitin(n12529),
            .carryinitout(bfn_14_24_0_));
    defparam IN_MUX_bfv_16_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_23_0_));
    defparam IN_MUX_bfv_16_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_24_0_ (
            .carryinitin(n12521),
            .carryinitout(bfn_16_24_0_));
    defparam IN_MUX_bfv_13_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_24_0_));
    defparam IN_MUX_bfv_11_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_24_0_));
    defparam IN_MUX_bfv_2_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_29_0_));
    defparam IN_MUX_bfv_2_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_30_0_ (
            .carryinitin(n12899),
            .carryinitout(bfn_2_30_0_));
    defparam IN_MUX_bfv_2_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_31_0_ (
            .carryinitin(n12907),
            .carryinitout(bfn_2_31_0_));
    defparam IN_MUX_bfv_2_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_32_0_ (
            .carryinitin(n12915),
            .carryinitout(bfn_2_32_0_));
    defparam IN_MUX_bfv_3_28_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_28_0_));
    defparam IN_MUX_bfv_3_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_29_0_ (
            .carryinitin(n12871),
            .carryinitout(bfn_3_29_0_));
    defparam IN_MUX_bfv_3_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_30_0_ (
            .carryinitin(n12879),
            .carryinitout(bfn_3_30_0_));
    defparam IN_MUX_bfv_3_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_31_0_ (
            .carryinitin(n12887),
            .carryinitout(bfn_3_31_0_));
    defparam IN_MUX_bfv_2_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_25_0_));
    defparam IN_MUX_bfv_2_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_26_0_ (
            .carryinitin(n12844),
            .carryinitout(bfn_2_26_0_));
    defparam IN_MUX_bfv_2_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_27_0_ (
            .carryinitin(n12852),
            .carryinitout(bfn_2_27_0_));
    defparam IN_MUX_bfv_2_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_28_0_ (
            .carryinitin(n12860),
            .carryinitout(bfn_2_28_0_));
    defparam IN_MUX_bfv_1_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_22_0_));
    defparam IN_MUX_bfv_1_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_23_0_ (
            .carryinitin(n12818),
            .carryinitout(bfn_1_23_0_));
    defparam IN_MUX_bfv_1_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_24_0_ (
            .carryinitin(n12826),
            .carryinitout(bfn_1_24_0_));
    defparam IN_MUX_bfv_1_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_25_0_ (
            .carryinitin(n12834),
            .carryinitout(bfn_1_25_0_));
    defparam IN_MUX_bfv_2_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_17_0_));
    defparam IN_MUX_bfv_2_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_18_0_ (
            .carryinitin(n12793),
            .carryinitout(bfn_2_18_0_));
    defparam IN_MUX_bfv_2_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_19_0_ (
            .carryinitin(n12801),
            .carryinitout(bfn_2_19_0_));
    defparam IN_MUX_bfv_2_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_20_0_ (
            .carryinitin(n12809),
            .carryinitout(bfn_2_20_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(n12769),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(n12777),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_2_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_16_0_ (
            .carryinitin(n12785),
            .carryinitout(bfn_2_16_0_));
    defparam IN_MUX_bfv_6_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_24_0_));
    defparam IN_MUX_bfv_6_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_25_0_ (
            .carryinitin(n12746),
            .carryinitout(bfn_6_25_0_));
    defparam IN_MUX_bfv_6_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_26_0_ (
            .carryinitin(n12754),
            .carryinitout(bfn_6_26_0_));
    defparam IN_MUX_bfv_6_21_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_21_0_));
    defparam IN_MUX_bfv_6_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_22_0_ (
            .carryinitin(n12724),
            .carryinitout(bfn_6_22_0_));
    defparam IN_MUX_bfv_6_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_23_0_ (
            .carryinitin(n12732),
            .carryinitout(bfn_6_23_0_));
    defparam IN_MUX_bfv_1_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_19_0_));
    defparam IN_MUX_bfv_1_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_20_0_ (
            .carryinitin(n12703),
            .carryinitout(bfn_1_20_0_));
    defparam IN_MUX_bfv_1_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_21_0_ (
            .carryinitin(n12711),
            .carryinitout(bfn_1_21_0_));
    defparam IN_MUX_bfv_3_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_14_0_));
    defparam IN_MUX_bfv_3_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_15_0_ (
            .carryinitin(n12683),
            .carryinitout(bfn_3_15_0_));
    defparam IN_MUX_bfv_3_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_16_0_ (
            .carryinitin(n12691),
            .carryinitout(bfn_3_16_0_));
    defparam IN_MUX_bfv_4_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_17_0_));
    defparam IN_MUX_bfv_4_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_18_0_ (
            .carryinitin(n12664),
            .carryinitout(bfn_4_18_0_));
    defparam IN_MUX_bfv_4_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_19_0_ (
            .carryinitin(n12672),
            .carryinitout(bfn_4_19_0_));
    defparam IN_MUX_bfv_6_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_17_0_));
    defparam IN_MUX_bfv_6_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_18_0_ (
            .carryinitin(n12646),
            .carryinitout(bfn_6_18_0_));
    defparam IN_MUX_bfv_6_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_19_0_ (
            .carryinitin(n12654),
            .carryinitout(bfn_6_19_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(n12629),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(n12637),
            .carryinitout(bfn_9_18_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(n12613),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(n12621),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_12_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_21_0_ (
            .carryinitin(n12598),
            .carryinitout(bfn_12_21_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(n12584),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_16_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_19_0_));
    defparam IN_MUX_bfv_16_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_20_0_ (
            .carryinitin(n12571),
            .carryinitout(bfn_16_20_0_));
    defparam IN_MUX_bfv_9_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_29_0_));
    defparam IN_MUX_bfv_1_31_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_31_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_31_0_));
    defparam IN_MUX_bfv_1_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_32_0_ (
            .carryinitin(\debounce.n13020 ),
            .carryinitout(bfn_1_32_0_));
    defparam IN_MUX_bfv_10_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_29_0_));
    defparam IN_MUX_bfv_10_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_30_0_ (
            .carryinitin(n13077),
            .carryinitout(bfn_10_30_0_));
    defparam IN_MUX_bfv_10_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_31_0_ (
            .carryinitin(n13085),
            .carryinitout(bfn_10_31_0_));
    defparam IN_MUX_bfv_10_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_32_0_ (
            .carryinitin(n13093),
            .carryinitout(bfn_10_32_0_));
    defparam IN_MUX_bfv_7_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_25_0_));
    defparam IN_MUX_bfv_7_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_26_0_ (
            .carryinitin(n12959),
            .carryinitout(bfn_7_26_0_));
    defparam IN_MUX_bfv_7_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_27_0_ (
            .carryinitin(n12967),
            .carryinitout(bfn_7_27_0_));
    defparam IN_MUX_bfv_10_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_22_0_));
    defparam IN_MUX_bfv_14_28_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_28_0_));
    defparam IN_MUX_bfv_14_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_29_0_ (
            .carryinitin(\PWM.n13029 ),
            .carryinitout(bfn_14_29_0_));
    defparam IN_MUX_bfv_14_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_30_0_ (
            .carryinitin(\PWM.n13037 ),
            .carryinitout(bfn_14_30_0_));
    defparam IN_MUX_bfv_14_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_31_0_ (
            .carryinitin(\PWM.n13045 ),
            .carryinitout(bfn_14_31_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__21684),
            .GLOBALBUFFEROUTPUT(CLK_N));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam i13072_1_lut_LC_1_18_1.C_ON=1'b0;
    defparam i13072_1_lut_LC_1_18_1.SEQ_MODE=4'b0000;
    defparam i13072_1_lut_LC_1_18_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 i13072_1_lut_LC_1_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35913),
            .lcout(n15802),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_2_lut_LC_1_19_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_2_lut_LC_1_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_2_lut_LC_1_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_2_lut_LC_1_19_0 (
            .in0(_gnd_net_),
            .in1(N__38349),
            .in2(_gnd_net_),
            .in3(N__21690),
            .lcout(n2401),
            .ltout(),
            .carryin(bfn_1_19_0_),
            .carryout(n12696),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_3_lut_LC_1_19_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_3_lut_LC_1_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_3_lut_LC_1_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_3_lut_LC_1_19_1 (
            .in0(_gnd_net_),
            .in1(N__55031),
            .in2(N__29123),
            .in3(N__21687),
            .lcout(n2400),
            .ltout(),
            .carryin(n12696),
            .carryout(n12697),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_4_lut_LC_1_19_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_4_lut_LC_1_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_4_lut_LC_1_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_4_lut_LC_1_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28737),
            .in3(N__21717),
            .lcout(n2399),
            .ltout(),
            .carryin(n12697),
            .carryout(n12698),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_5_lut_LC_1_19_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_5_lut_LC_1_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_5_lut_LC_1_19_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_5_lut_LC_1_19_3 (
            .in0(_gnd_net_),
            .in1(N__55032),
            .in2(N__28637),
            .in3(N__21714),
            .lcout(n2398),
            .ltout(),
            .carryin(n12698),
            .carryout(n12699),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_6_lut_LC_1_19_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_6_lut_LC_1_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_6_lut_LC_1_19_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_6_lut_LC_1_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28832),
            .in3(N__21711),
            .lcout(n2397),
            .ltout(),
            .carryin(n12699),
            .carryout(n12700),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_7_lut_LC_1_19_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_7_lut_LC_1_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_7_lut_LC_1_19_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_7_lut_LC_1_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25904),
            .in3(N__21708),
            .lcout(n2396),
            .ltout(),
            .carryin(n12700),
            .carryout(n12701),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_8_lut_LC_1_19_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_8_lut_LC_1_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_8_lut_LC_1_19_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_8_lut_LC_1_19_6 (
            .in0(_gnd_net_),
            .in1(N__55418),
            .in2(N__25875),
            .in3(N__21705),
            .lcout(n2395),
            .ltout(),
            .carryin(n12701),
            .carryout(n12702),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_9_lut_LC_1_19_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_9_lut_LC_1_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_9_lut_LC_1_19_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_9_lut_LC_1_19_7 (
            .in0(_gnd_net_),
            .in1(N__55033),
            .in2(N__25782),
            .in3(N__21702),
            .lcout(n2394),
            .ltout(),
            .carryin(n12702),
            .carryout(n12703),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_10_lut_LC_1_20_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_10_lut_LC_1_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_10_lut_LC_1_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_10_lut_LC_1_20_0 (
            .in0(_gnd_net_),
            .in1(N__55476),
            .in2(N__28863),
            .in3(N__21699),
            .lcout(n2393),
            .ltout(),
            .carryin(bfn_1_20_0_),
            .carryout(n12704),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_11_lut_LC_1_20_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_11_lut_LC_1_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_11_lut_LC_1_20_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_11_lut_LC_1_20_1 (
            .in0(_gnd_net_),
            .in1(N__55485),
            .in2(N__25653),
            .in3(N__21696),
            .lcout(n2392),
            .ltout(),
            .carryin(n12704),
            .carryout(n12705),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_12_lut_LC_1_20_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_12_lut_LC_1_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_12_lut_LC_1_20_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_12_lut_LC_1_20_2 (
            .in0(_gnd_net_),
            .in1(N__55477),
            .in2(N__23463),
            .in3(N__21693),
            .lcout(n2391),
            .ltout(),
            .carryin(n12705),
            .carryout(n12706),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_13_lut_LC_1_20_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_13_lut_LC_1_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_13_lut_LC_1_20_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_13_lut_LC_1_20_3 (
            .in0(_gnd_net_),
            .in1(N__55486),
            .in2(N__28922),
            .in3(N__21744),
            .lcout(n2390),
            .ltout(),
            .carryin(n12706),
            .carryout(n12707),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_14_lut_LC_1_20_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_14_lut_LC_1_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_14_lut_LC_1_20_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_14_lut_LC_1_20_4 (
            .in0(_gnd_net_),
            .in1(N__55478),
            .in2(N__28791),
            .in3(N__21741),
            .lcout(n2389),
            .ltout(),
            .carryin(n12707),
            .carryout(n12708),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_15_lut_LC_1_20_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_15_lut_LC_1_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_15_lut_LC_1_20_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_15_lut_LC_1_20_5 (
            .in0(_gnd_net_),
            .in1(N__28688),
            .in2(N__55548),
            .in3(N__21738),
            .lcout(n2388),
            .ltout(),
            .carryin(n12708),
            .carryout(n12709),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_16_lut_LC_1_20_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_16_lut_LC_1_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_16_lut_LC_1_20_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_16_lut_LC_1_20_6 (
            .in0(_gnd_net_),
            .in1(N__25623),
            .in2(N__55550),
            .in3(N__21735),
            .lcout(n2387),
            .ltout(),
            .carryin(n12709),
            .carryout(n12710),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_17_lut_LC_1_20_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_17_lut_LC_1_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_17_lut_LC_1_20_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_17_lut_LC_1_20_7 (
            .in0(_gnd_net_),
            .in1(N__23439),
            .in2(N__55549),
            .in3(N__21732),
            .lcout(n2386),
            .ltout(),
            .carryin(n12710),
            .carryout(n12711),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_18_lut_LC_1_21_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_18_lut_LC_1_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_18_lut_LC_1_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_18_lut_LC_1_21_0 (
            .in0(_gnd_net_),
            .in1(N__28979),
            .in2(N__54721),
            .in3(N__21729),
            .lcout(n2385),
            .ltout(),
            .carryin(bfn_1_21_0_),
            .carryout(n12712),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_19_lut_LC_1_21_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_19_lut_LC_1_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_19_lut_LC_1_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_19_lut_LC_1_21_1 (
            .in0(_gnd_net_),
            .in1(N__29024),
            .in2(N__54724),
            .in3(N__21726),
            .lcout(n2384),
            .ltout(),
            .carryin(n12712),
            .carryout(n12713),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_20_lut_LC_1_21_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_20_lut_LC_1_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_20_lut_LC_1_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_20_lut_LC_1_21_2 (
            .in0(_gnd_net_),
            .in1(N__25731),
            .in2(N__54722),
            .in3(N__21723),
            .lcout(n2383),
            .ltout(),
            .carryin(n12713),
            .carryout(n12714),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_21_lut_LC_1_21_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_21_lut_LC_1_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_21_lut_LC_1_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_21_lut_LC_1_21_3 (
            .in0(_gnd_net_),
            .in1(N__30963),
            .in2(N__54725),
            .in3(N__21720),
            .lcout(n2382),
            .ltout(),
            .carryin(n12714),
            .carryout(n12715),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_22_lut_LC_1_21_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1570_22_lut_LC_1_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_22_lut_LC_1_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1570_22_lut_LC_1_21_4 (
            .in0(_gnd_net_),
            .in1(N__25695),
            .in2(N__54723),
            .in3(N__21771),
            .lcout(n2381),
            .ltout(),
            .carryin(n12715),
            .carryout(n12716),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1570_23_lut_LC_1_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1570_23_lut_LC_1_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1570_23_lut_LC_1_21_5.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1570_23_lut_LC_1_21_5 (
            .in0(N__54324),
            .in1(N__35765),
            .in2(N__25812),
            .in3(N__21768),
            .lcout(n2412),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_2_lut_LC_1_22_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_2_lut_LC_1_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_2_lut_LC_1_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_2_lut_LC_1_22_0 (
            .in0(_gnd_net_),
            .in1(N__33501),
            .in2(_gnd_net_),
            .in3(N__21765),
            .lcout(n2901),
            .ltout(),
            .carryin(bfn_1_22_0_),
            .carryout(n12811),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_3_lut_LC_1_22_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_3_lut_LC_1_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_3_lut_LC_1_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_3_lut_LC_1_22_1 (
            .in0(_gnd_net_),
            .in1(N__54708),
            .in2(N__26577),
            .in3(N__21762),
            .lcout(n2900),
            .ltout(),
            .carryin(n12811),
            .carryout(n12812),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_4_lut_LC_1_22_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_4_lut_LC_1_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_4_lut_LC_1_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_4_lut_LC_1_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29460),
            .in3(N__21759),
            .lcout(n2899),
            .ltout(),
            .carryin(n12812),
            .carryout(n12813),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_5_lut_LC_1_22_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_5_lut_LC_1_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_5_lut_LC_1_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_5_lut_LC_1_22_3 (
            .in0(_gnd_net_),
            .in1(N__54709),
            .in2(N__29649),
            .in3(N__21756),
            .lcout(n2898),
            .ltout(),
            .carryin(n12813),
            .carryout(n12814),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_6_lut_LC_1_22_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_6_lut_LC_1_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_6_lut_LC_1_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_6_lut_LC_1_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26544),
            .in3(N__21753),
            .lcout(n2897),
            .ltout(),
            .carryin(n12814),
            .carryout(n12815),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_7_lut_LC_1_22_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_7_lut_LC_1_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_7_lut_LC_1_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_7_lut_LC_1_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29884),
            .in3(N__21750),
            .lcout(n2896),
            .ltout(),
            .carryin(n12815),
            .carryout(n12816),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_8_lut_LC_1_22_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_8_lut_LC_1_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_8_lut_LC_1_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_8_lut_LC_1_22_6 (
            .in0(_gnd_net_),
            .in1(N__22757),
            .in2(N__55030),
            .in3(N__21747),
            .lcout(n2895),
            .ltout(),
            .carryin(n12816),
            .carryout(n12817),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_9_lut_LC_1_22_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_9_lut_LC_1_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_9_lut_LC_1_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_9_lut_LC_1_22_7 (
            .in0(_gnd_net_),
            .in1(N__54713),
            .in2(N__24584),
            .in3(N__21798),
            .lcout(n2894),
            .ltout(),
            .carryin(n12817),
            .carryout(n12818),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_10_lut_LC_1_23_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_10_lut_LC_1_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_10_lut_LC_1_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_10_lut_LC_1_23_0 (
            .in0(_gnd_net_),
            .in1(N__54283),
            .in2(N__29732),
            .in3(N__21795),
            .lcout(n2893),
            .ltout(),
            .carryin(bfn_1_23_0_),
            .carryout(n12819),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_11_lut_LC_1_23_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_11_lut_LC_1_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_11_lut_LC_1_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_11_lut_LC_1_23_1 (
            .in0(_gnd_net_),
            .in1(N__26740),
            .in2(N__54705),
            .in3(N__21792),
            .lcout(n2892),
            .ltout(),
            .carryin(n12819),
            .carryout(n12820),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_12_lut_LC_1_23_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_12_lut_LC_1_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_12_lut_LC_1_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_12_lut_LC_1_23_2 (
            .in0(_gnd_net_),
            .in1(N__54287),
            .in2(N__29336),
            .in3(N__21789),
            .lcout(n2891),
            .ltout(),
            .carryin(n12820),
            .carryout(n12821),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_13_lut_LC_1_23_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_13_lut_LC_1_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_13_lut_LC_1_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_13_lut_LC_1_23_3 (
            .in0(_gnd_net_),
            .in1(N__54292),
            .in2(N__24621),
            .in3(N__21786),
            .lcout(n2890),
            .ltout(),
            .carryin(n12821),
            .carryout(n12822),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_14_lut_LC_1_23_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_14_lut_LC_1_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_14_lut_LC_1_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_14_lut_LC_1_23_4 (
            .in0(_gnd_net_),
            .in1(N__54288),
            .in2(N__24542),
            .in3(N__21783),
            .lcout(n2889),
            .ltout(),
            .carryin(n12822),
            .carryout(n12823),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_15_lut_LC_1_23_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_15_lut_LC_1_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_15_lut_LC_1_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_15_lut_LC_1_23_5 (
            .in0(_gnd_net_),
            .in1(N__54293),
            .in2(N__29831),
            .in3(N__21780),
            .lcout(n2888),
            .ltout(),
            .carryin(n12823),
            .carryout(n12824),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_16_lut_LC_1_23_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_16_lut_LC_1_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_16_lut_LC_1_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_16_lut_LC_1_23_6 (
            .in0(_gnd_net_),
            .in1(N__24309),
            .in2(N__54707),
            .in3(N__21777),
            .lcout(n2887),
            .ltout(),
            .carryin(n12824),
            .carryout(n12825),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_17_lut_LC_1_23_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_17_lut_LC_1_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_17_lut_LC_1_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_17_lut_LC_1_23_7 (
            .in0(_gnd_net_),
            .in1(N__26844),
            .in2(N__54706),
            .in3(N__21774),
            .lcout(n2886),
            .ltout(),
            .carryin(n12825),
            .carryout(n12826),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_18_lut_LC_1_24_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_18_lut_LC_1_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_18_lut_LC_1_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_18_lut_LC_1_24_0 (
            .in0(_gnd_net_),
            .in1(N__26292),
            .in2(N__54240),
            .in3(N__21825),
            .lcout(n2885),
            .ltout(),
            .carryin(bfn_1_24_0_),
            .carryout(n12827),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_19_lut_LC_1_24_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_19_lut_LC_1_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_19_lut_LC_1_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_19_lut_LC_1_24_1 (
            .in0(_gnd_net_),
            .in1(N__27235),
            .in2(N__55275),
            .in3(N__21822),
            .lcout(n2884),
            .ltout(),
            .carryin(n12827),
            .carryout(n12828),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_20_lut_LC_1_24_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_20_lut_LC_1_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_20_lut_LC_1_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_20_lut_LC_1_24_2 (
            .in0(_gnd_net_),
            .in1(N__26337),
            .in2(N__54241),
            .in3(N__21819),
            .lcout(n2883),
            .ltout(),
            .carryin(n12828),
            .carryout(n12829),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_21_lut_LC_1_24_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_21_lut_LC_1_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_21_lut_LC_1_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_21_lut_LC_1_24_3 (
            .in0(_gnd_net_),
            .in1(N__53834),
            .in2(N__26504),
            .in3(N__21816),
            .lcout(n2882),
            .ltout(),
            .carryin(n12829),
            .carryout(n12830),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_22_lut_LC_1_24_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_22_lut_LC_1_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_22_lut_LC_1_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_22_lut_LC_1_24_4 (
            .in0(_gnd_net_),
            .in1(N__29767),
            .in2(N__54242),
            .in3(N__21813),
            .lcout(n2881),
            .ltout(),
            .carryin(n12830),
            .carryout(n12831),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_23_lut_LC_1_24_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_23_lut_LC_1_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_23_lut_LC_1_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_23_lut_LC_1_24_5 (
            .in0(_gnd_net_),
            .in1(N__26447),
            .in2(N__55276),
            .in3(N__21810),
            .lcout(n2880),
            .ltout(),
            .carryin(n12831),
            .carryout(n12832),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_24_lut_LC_1_24_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_24_lut_LC_1_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_24_lut_LC_1_24_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_24_lut_LC_1_24_6 (
            .in0(_gnd_net_),
            .in1(N__26471),
            .in2(N__54243),
            .in3(N__21807),
            .lcout(n2879),
            .ltout(),
            .carryin(n12832),
            .carryout(n12833),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_25_lut_LC_1_24_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_25_lut_LC_1_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_25_lut_LC_1_24_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_25_lut_LC_1_24_7 (
            .in0(_gnd_net_),
            .in1(N__26418),
            .in2(N__55277),
            .in3(N__21804),
            .lcout(n2878),
            .ltout(),
            .carryin(n12833),
            .carryout(n12834),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_26_lut_LC_1_25_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_26_lut_LC_1_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_26_lut_LC_1_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_26_lut_LC_1_25_0 (
            .in0(_gnd_net_),
            .in1(N__26901),
            .in2(N__54654),
            .in3(N__21801),
            .lcout(n2877),
            .ltout(),
            .carryin(bfn_1_25_0_),
            .carryout(n12835),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_27_lut_LC_1_25_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1905_27_lut_LC_1_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_27_lut_LC_1_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1905_27_lut_LC_1_25_1 (
            .in0(_gnd_net_),
            .in1(N__26402),
            .in2(N__54655),
            .in3(N__21858),
            .lcout(n2876),
            .ltout(),
            .carryin(n12835),
            .carryout(n12836),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1905_28_lut_LC_1_25_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1905_28_lut_LC_1_25_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1905_28_lut_LC_1_25_2.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1905_28_lut_LC_1_25_2 (
            .in0(N__54236),
            .in1(N__34352),
            .in2(N__26367),
            .in3(N__21855),
            .lcout(n2907),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1914_3_lut_LC_1_25_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1914_3_lut_LC_1_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1914_3_lut_LC_1_25_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1914_3_lut_LC_1_25_4 (
            .in0(_gnd_net_),
            .in1(N__26500),
            .in2(N__34333),
            .in3(N__21852),
            .lcout(n2914),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1932_3_lut_LC_1_25_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1932_3_lut_LC_1_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1932_3_lut_LC_1_25_5.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1932_3_lut_LC_1_25_5 (
            .in0(N__26572),
            .in1(_gnd_net_),
            .in2(N__21846),
            .in3(N__34316),
            .lcout(n2932),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1847_3_lut_LC_1_25_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1847_3_lut_LC_1_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1847_3_lut_LC_1_25_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 encoder0_position_31__I_0_i1847_3_lut_LC_1_25_6 (
            .in0(_gnd_net_),
            .in1(N__36411),
            .in2(N__22365),
            .in3(N__22845),
            .lcout(n2815),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1778_3_lut_LC_1_25_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1778_3_lut_LC_1_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1778_3_lut_LC_1_25_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1778_3_lut_LC_1_25_7 (
            .in0(_gnd_net_),
            .in1(N__22245),
            .in2(N__29688),
            .in3(N__36295),
            .lcout(n2714),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.reg_out_i0_i0_LC_1_26_0 .C_ON=1'b0;
    defparam \debounce.reg_out_i0_i0_LC_1_26_0 .SEQ_MODE=4'b1000;
    defparam \debounce.reg_out_i0_i0_LC_1_26_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \debounce.reg_out_i0_i0_LC_1_26_0  (
            .in0(N__46927),
            .in1(N__21921),
            .in2(_gnd_net_),
            .in3(N__38870),
            .lcout(h3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56199),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1908_3_lut_LC_1_26_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1908_3_lut_LC_1_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1908_3_lut_LC_1_26_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1908_3_lut_LC_1_26_1 (
            .in0(_gnd_net_),
            .in1(N__21834),
            .in2(N__34335),
            .in3(N__26403),
            .lcout(n2908),
            .ltout(n2908_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1975_3_lut_LC_1_26_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1975_3_lut_LC_1_26_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1975_3_lut_LC_1_26_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1975_3_lut_LC_1_26_2 (
            .in0(N__34513),
            .in1(_gnd_net_),
            .in2(N__21828),
            .in3(N__23028),
            .lcout(n3007),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1865_3_lut_LC_1_26_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1865_3_lut_LC_1_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1865_3_lut_LC_1_26_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1865_3_lut_LC_1_26_3 (
            .in0(N__22296),
            .in1(N__33539),
            .in2(_gnd_net_),
            .in3(N__36417),
            .lcout(n2833),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1927_3_lut_LC_1_26_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1927_3_lut_LC_1_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1927_3_lut_LC_1_26_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1927_3_lut_LC_1_26_4 (
            .in0(_gnd_net_),
            .in1(N__21879),
            .in2(N__22761),
            .in3(N__34328),
            .lcout(n2927),
            .ltout(n2927_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1994_3_lut_LC_1_26_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1994_3_lut_LC_1_26_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1994_3_lut_LC_1_26_5.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1994_3_lut_LC_1_26_5 (
            .in0(N__22881),
            .in1(_gnd_net_),
            .in2(N__21867),
            .in3(N__34512),
            .lcout(n3026),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1993_3_lut_LC_1_27_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1993_3_lut_LC_1_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1993_3_lut_LC_1_27_0.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1993_3_lut_LC_1_27_0 (
            .in0(N__22962),
            .in1(_gnd_net_),
            .in2(N__34509),
            .in3(N__26781),
            .lcout(n3025),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1990_3_lut_LC_1_27_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1990_3_lut_LC_1_27_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1990_3_lut_LC_1_27_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1990_3_lut_LC_1_27_1 (
            .in0(_gnd_net_),
            .in1(N__29301),
            .in2(N__22941),
            .in3(N__34483),
            .lcout(n3022),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1985_3_lut_LC_1_27_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1985_3_lut_LC_1_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1985_3_lut_LC_1_27_2.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i1985_3_lut_LC_1_27_2 (
            .in0(N__26817),
            .in1(N__23004),
            .in2(N__34511),
            .in3(_gnd_net_),
            .lcout(n3017),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1992_3_lut_LC_1_27_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1992_3_lut_LC_1_27_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1992_3_lut_LC_1_27_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1992_3_lut_LC_1_27_3 (
            .in0(_gnd_net_),
            .in1(N__22953),
            .in2(N__29715),
            .in3(N__34493),
            .lcout(n3024),
            .ltout(n3024_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_166_LC_1_27_4.C_ON=1'b0;
    defparam i1_4_lut_adj_166_LC_1_27_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_166_LC_1_27_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_166_LC_1_27_4 (
            .in0(N__24736),
            .in1(N__24935),
            .in2(N__21864),
            .in3(N__24778),
            .lcout(),
            .ltout(n14730_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_168_LC_1_27_5.C_ON=1'b0;
    defparam i1_4_lut_adj_168_LC_1_27_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_168_LC_1_27_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_168_LC_1_27_5 (
            .in0(N__24880),
            .in1(N__27278),
            .in2(N__21861),
            .in3(N__21897),
            .lcout(n14736),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1989_3_lut_LC_1_27_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1989_3_lut_LC_1_27_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1989_3_lut_LC_1_27_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1989_3_lut_LC_1_27_6 (
            .in0(_gnd_net_),
            .in1(N__22929),
            .in2(N__34510),
            .in3(N__26682),
            .lcout(n3021),
            .ltout(n3021_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_165_LC_1_27_7.C_ON=1'b0;
    defparam i1_3_lut_adj_165_LC_1_27_7.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_165_LC_1_27_7.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_165_LC_1_27_7 (
            .in0(_gnd_net_),
            .in1(N__25006),
            .in2(N__21900),
            .in3(N__24830),
            .lcout(n14728),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_174_LC_1_28_0.C_ON=1'b0;
    defparam i1_4_lut_adj_174_LC_1_28_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_174_LC_1_28_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_174_LC_1_28_0 (
            .in0(N__27968),
            .in1(N__32905),
            .in2(N__30811),
            .in3(N__27802),
            .lcout(),
            .ltout(n14150_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_176_LC_1_28_1.C_ON=1'b0;
    defparam i1_4_lut_adj_176_LC_1_28_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_176_LC_1_28_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_176_LC_1_28_1 (
            .in0(N__30658),
            .in1(N__21885),
            .in2(N__21891),
            .in3(N__21975),
            .lcout(n14156),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1977_3_lut_LC_1_28_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1977_3_lut_LC_1_28_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1977_3_lut_LC_1_28_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1977_3_lut_LC_1_28_3 (
            .in0(_gnd_net_),
            .in1(N__27072),
            .in2(N__22974),
            .in3(N__34514),
            .lcout(n3009),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2062_3_lut_LC_1_28_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2062_3_lut_LC_1_28_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2062_3_lut_LC_1_28_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2062_3_lut_LC_1_28_4 (
            .in0(_gnd_net_),
            .in1(N__24804),
            .in2(N__30597),
            .in3(N__34710),
            .lcout(n3126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2064_3_lut_LC_1_28_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2064_3_lut_LC_1_28_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2064_3_lut_LC_1_28_5.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i2064_3_lut_LC_1_28_5 (
            .in0(N__24843),
            .in1(_gnd_net_),
            .in2(N__34716),
            .in3(N__29958),
            .lcout(n3128),
            .ltout(n3128_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_175_LC_1_28_6.C_ON=1'b0;
    defparam i1_4_lut_adj_175_LC_1_28_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_175_LC_1_28_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_175_LC_1_28_6 (
            .in0(N__27676),
            .in1(N__27751),
            .in2(N__21888),
            .in3(N__27735),
            .lcout(n14148),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.reg_B_i0_LC_1_28_7 .C_ON=1'b0;
    defparam \debounce.reg_B_i0_LC_1_28_7 .SEQ_MODE=4'b1000;
    defparam \debounce.reg_B_i0_LC_1_28_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debounce.reg_B_i0_LC_1_28_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21942),
            .lcout(reg_B_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56203),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2054_3_lut_LC_1_29_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2054_3_lut_LC_1_29_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2054_3_lut_LC_1_29_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i2054_3_lut_LC_1_29_0 (
            .in0(_gnd_net_),
            .in1(N__30623),
            .in2(N__34708),
            .in3(N__24903),
            .lcout(n3118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2060_3_lut_LC_1_29_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2060_3_lut_LC_1_29_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2060_3_lut_LC_1_29_2.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i2060_3_lut_LC_1_29_2 (
            .in0(N__24746),
            .in1(_gnd_net_),
            .in2(N__34709),
            .in3(N__24723),
            .lcout(n3124),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2056_3_lut_LC_1_29_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2056_3_lut_LC_1_29_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2056_3_lut_LC_1_29_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2056_3_lut_LC_1_29_3 (
            .in0(_gnd_net_),
            .in1(N__24951),
            .in2(N__24978),
            .in3(N__34681),
            .lcout(n3120),
            .ltout(n3120_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2123_3_lut_LC_1_29_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2123_3_lut_LC_1_29_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2123_3_lut_LC_1_29_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2123_3_lut_LC_1_29_4 (
            .in0(_gnd_net_),
            .in1(N__23085),
            .in2(N__21981),
            .in3(N__34911),
            .lcout(n3219),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2058_3_lut_LC_1_29_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2058_3_lut_LC_1_29_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2058_3_lut_LC_1_29_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2058_3_lut_LC_1_29_5 (
            .in0(_gnd_net_),
            .in1(N__30560),
            .in2(N__25035),
            .in3(N__34686),
            .lcout(n3122),
            .ltout(n3122_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_173_LC_1_29_6.C_ON=1'b0;
    defparam i1_4_lut_adj_173_LC_1_29_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_173_LC_1_29_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_173_LC_1_29_6 (
            .in0(N__30883),
            .in1(N__23096),
            .in2(N__21978),
            .in3(N__27544),
            .lcout(n14146),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2059_3_lut_LC_1_29_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2059_3_lut_LC_1_29_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2059_3_lut_LC_1_29_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2059_3_lut_LC_1_29_7 (
            .in0(_gnd_net_),
            .in1(N__24707),
            .in2(N__24687),
            .in3(N__34682),
            .lcout(n3123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.reg_B_i2_LC_1_30_0 .C_ON=1'b0;
    defparam \debounce.reg_B_i2_LC_1_30_0 .SEQ_MODE=4'b1000;
    defparam \debounce.reg_B_i2_LC_1_30_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \debounce.reg_B_i2_LC_1_30_0  (
            .in0(N__21969),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(reg_B_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56207),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.reg_B_i1_LC_1_30_1 .C_ON=1'b0;
    defparam \debounce.reg_B_i1_LC_1_30_1 .SEQ_MODE=4'b1000;
    defparam \debounce.reg_B_i1_LC_1_30_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \debounce.reg_B_i1_LC_1_30_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21959),
            .lcout(reg_B_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56207),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.i2_4_lut_LC_1_30_2 .C_ON=1'b0;
    defparam \debounce.i2_4_lut_LC_1_30_2 .SEQ_MODE=4'b0000;
    defparam \debounce.i2_4_lut_LC_1_30_2 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \debounce.i2_4_lut_LC_1_30_2  (
            .in0(N__21968),
            .in1(N__38885),
            .in2(N__21960),
            .in3(N__22070),
            .lcout(),
            .ltout(\debounce.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.i3_4_lut_LC_1_30_3 .C_ON=1'b0;
    defparam \debounce.i3_4_lut_LC_1_30_3 .SEQ_MODE=4'b0000;
    defparam \debounce.i3_4_lut_LC_1_30_3 .LUT_INIT=16'b1111011011111111;
    LogicCell40 \debounce.i3_4_lut_LC_1_30_3  (
            .in0(N__21941),
            .in1(N__21920),
            .in2(N__21903),
            .in3(N__38857),
            .lcout(\debounce.cnt_next_9__N_424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.i7_4_lut_LC_1_30_4 .C_ON=1'b0;
    defparam \debounce.i7_4_lut_LC_1_30_4 .SEQ_MODE=4'b0000;
    defparam \debounce.i7_4_lut_LC_1_30_4 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \debounce.i7_4_lut_LC_1_30_4  (
            .in0(N__21995),
            .in1(N__22149),
            .in2(N__22128),
            .in3(N__22193),
            .lcout(\debounce.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.i6_4_lut_LC_1_30_5 .C_ON=1'b0;
    defparam \debounce.i6_4_lut_LC_1_30_5 .SEQ_MODE=4'b0000;
    defparam \debounce.i6_4_lut_LC_1_30_5 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \debounce.i6_4_lut_LC_1_30_5  (
            .in0(N__22163),
            .in1(N__22058),
            .in2(N__22029),
            .in3(N__22043),
            .lcout(),
            .ltout(\debounce.n16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.i9_4_lut_LC_1_30_6 .C_ON=1'b0;
    defparam \debounce.i9_4_lut_LC_1_30_6 .SEQ_MODE=4'b0000;
    defparam \debounce.i9_4_lut_LC_1_30_6 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \debounce.i9_4_lut_LC_1_30_6  (
            .in0(N__22010),
            .in1(N__22178),
            .in2(N__22080),
            .in3(N__22077),
            .lcout(n14129),
            .ltout(n14129_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.reg_out_i0_i2_LC_1_30_7 .C_ON=1'b0;
    defparam \debounce.reg_out_i0_i2_LC_1_30_7 .SEQ_MODE=4'b1000;
    defparam \debounce.reg_out_i0_i2_LC_1_30_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \debounce.reg_out_i0_i2_LC_1_30_7  (
            .in0(N__22071),
            .in1(_gnd_net_),
            .in2(N__22062),
            .in3(N__46866),
            .lcout(h1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56207),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.cnt_reg_665__i0_LC_1_31_0 .C_ON=1'b1;
    defparam \debounce.cnt_reg_665__i0_LC_1_31_0 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_665__i0_LC_1_31_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_665__i0_LC_1_31_0  (
            .in0(_gnd_net_),
            .in1(N__22059),
            .in2(_gnd_net_),
            .in3(N__22047),
            .lcout(\debounce.cnt_reg_0 ),
            .ltout(),
            .carryin(bfn_1_31_0_),
            .carryout(\debounce.n13013 ),
            .clk(N__56208),
            .ce(),
            .sr(N__22106));
    defparam \debounce.cnt_reg_665__i1_LC_1_31_1 .C_ON=1'b1;
    defparam \debounce.cnt_reg_665__i1_LC_1_31_1 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_665__i1_LC_1_31_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_665__i1_LC_1_31_1  (
            .in0(_gnd_net_),
            .in1(N__22044),
            .in2(_gnd_net_),
            .in3(N__22032),
            .lcout(\debounce.cnt_reg_1 ),
            .ltout(),
            .carryin(\debounce.n13013 ),
            .carryout(\debounce.n13014 ),
            .clk(N__56208),
            .ce(),
            .sr(N__22106));
    defparam \debounce.cnt_reg_665__i2_LC_1_31_2 .C_ON=1'b1;
    defparam \debounce.cnt_reg_665__i2_LC_1_31_2 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_665__i2_LC_1_31_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_665__i2_LC_1_31_2  (
            .in0(_gnd_net_),
            .in1(N__22028),
            .in2(_gnd_net_),
            .in3(N__22014),
            .lcout(\debounce.cnt_reg_2 ),
            .ltout(),
            .carryin(\debounce.n13014 ),
            .carryout(\debounce.n13015 ),
            .clk(N__56208),
            .ce(),
            .sr(N__22106));
    defparam \debounce.cnt_reg_665__i3_LC_1_31_3 .C_ON=1'b1;
    defparam \debounce.cnt_reg_665__i3_LC_1_31_3 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_665__i3_LC_1_31_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_665__i3_LC_1_31_3  (
            .in0(_gnd_net_),
            .in1(N__22011),
            .in2(_gnd_net_),
            .in3(N__21999),
            .lcout(\debounce.cnt_reg_3 ),
            .ltout(),
            .carryin(\debounce.n13015 ),
            .carryout(\debounce.n13016 ),
            .clk(N__56208),
            .ce(),
            .sr(N__22106));
    defparam \debounce.cnt_reg_665__i4_LC_1_31_4 .C_ON=1'b1;
    defparam \debounce.cnt_reg_665__i4_LC_1_31_4 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_665__i4_LC_1_31_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_665__i4_LC_1_31_4  (
            .in0(_gnd_net_),
            .in1(N__21996),
            .in2(_gnd_net_),
            .in3(N__21984),
            .lcout(\debounce.cnt_reg_4 ),
            .ltout(),
            .carryin(\debounce.n13016 ),
            .carryout(\debounce.n13017 ),
            .clk(N__56208),
            .ce(),
            .sr(N__22106));
    defparam \debounce.cnt_reg_665__i5_LC_1_31_5 .C_ON=1'b1;
    defparam \debounce.cnt_reg_665__i5_LC_1_31_5 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_665__i5_LC_1_31_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_665__i5_LC_1_31_5  (
            .in0(_gnd_net_),
            .in1(N__22194),
            .in2(_gnd_net_),
            .in3(N__22182),
            .lcout(\debounce.cnt_reg_5 ),
            .ltout(),
            .carryin(\debounce.n13017 ),
            .carryout(\debounce.n13018 ),
            .clk(N__56208),
            .ce(),
            .sr(N__22106));
    defparam \debounce.cnt_reg_665__i6_LC_1_31_6 .C_ON=1'b1;
    defparam \debounce.cnt_reg_665__i6_LC_1_31_6 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_665__i6_LC_1_31_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_665__i6_LC_1_31_6  (
            .in0(_gnd_net_),
            .in1(N__22179),
            .in2(_gnd_net_),
            .in3(N__22167),
            .lcout(\debounce.cnt_reg_6 ),
            .ltout(),
            .carryin(\debounce.n13018 ),
            .carryout(\debounce.n13019 ),
            .clk(N__56208),
            .ce(),
            .sr(N__22106));
    defparam \debounce.cnt_reg_665__i7_LC_1_31_7 .C_ON=1'b1;
    defparam \debounce.cnt_reg_665__i7_LC_1_31_7 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_665__i7_LC_1_31_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_665__i7_LC_1_31_7  (
            .in0(_gnd_net_),
            .in1(N__22164),
            .in2(_gnd_net_),
            .in3(N__22152),
            .lcout(\debounce.cnt_reg_7 ),
            .ltout(),
            .carryin(\debounce.n13019 ),
            .carryout(\debounce.n13020 ),
            .clk(N__56208),
            .ce(),
            .sr(N__22106));
    defparam \debounce.cnt_reg_665__i8_LC_1_32_0 .C_ON=1'b1;
    defparam \debounce.cnt_reg_665__i8_LC_1_32_0 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_665__i8_LC_1_32_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_665__i8_LC_1_32_0  (
            .in0(_gnd_net_),
            .in1(N__22148),
            .in2(_gnd_net_),
            .in3(N__22134),
            .lcout(\debounce.cnt_reg_8 ),
            .ltout(),
            .carryin(bfn_1_32_0_),
            .carryout(\debounce.n13021 ),
            .clk(N__56210),
            .ce(),
            .sr(N__22110));
    defparam \debounce.cnt_reg_665__i9_LC_1_32_1 .C_ON=1'b0;
    defparam \debounce.cnt_reg_665__i9_LC_1_32_1 .SEQ_MODE=4'b1000;
    defparam \debounce.cnt_reg_665__i9_LC_1_32_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \debounce.cnt_reg_665__i9_LC_1_32_1  (
            .in0(_gnd_net_),
            .in1(N__22124),
            .in2(_gnd_net_),
            .in3(N__22131),
            .lcout(\debounce.cnt_reg_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56210),
            .ce(),
            .sr(N__22110));
    defparam encoder0_position_31__I_0_add_1771_2_lut_LC_2_13_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_2_lut_LC_2_13_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_2_lut_LC_2_13_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_2_lut_LC_2_13_0 (
            .in0(_gnd_net_),
            .in1(N__33582),
            .in2(_gnd_net_),
            .in3(N__22089),
            .lcout(n2701),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(n12762),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_3_lut_LC_2_13_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_3_lut_LC_2_13_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_3_lut_LC_2_13_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_3_lut_LC_2_13_1 (
            .in0(_gnd_net_),
            .in1(N__26265),
            .in2(N__55563),
            .in3(N__22086),
            .lcout(n2700),
            .ltout(),
            .carryin(n12762),
            .carryout(n12763),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_4_lut_LC_2_13_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_4_lut_LC_2_13_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_4_lut_LC_2_13_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_4_lut_LC_2_13_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29259),
            .in3(N__22083),
            .lcout(n2699),
            .ltout(),
            .carryin(n12763),
            .carryout(n12764),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_5_lut_LC_2_13_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_5_lut_LC_2_13_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_5_lut_LC_2_13_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_5_lut_LC_2_13_3 (
            .in0(_gnd_net_),
            .in1(N__55436),
            .in2(N__29196),
            .in3(N__22224),
            .lcout(n2698),
            .ltout(),
            .carryin(n12764),
            .carryout(n12765),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_6_lut_LC_2_13_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_6_lut_LC_2_13_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_6_lut_LC_2_13_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_6_lut_LC_2_13_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29439),
            .in3(N__22221),
            .lcout(n2697),
            .ltout(),
            .carryin(n12765),
            .carryout(n12766),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_7_lut_LC_2_13_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_7_lut_LC_2_13_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_7_lut_LC_2_13_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_7_lut_LC_2_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29508),
            .in3(N__22218),
            .lcout(n2696),
            .ltout(),
            .carryin(n12766),
            .carryout(n12767),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_8_lut_LC_2_13_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_8_lut_LC_2_13_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_8_lut_LC_2_13_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_8_lut_LC_2_13_6 (
            .in0(_gnd_net_),
            .in1(N__55562),
            .in2(N__23589),
            .in3(N__22215),
            .lcout(n2695),
            .ltout(),
            .carryin(n12767),
            .carryout(n12768),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_9_lut_LC_2_13_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_9_lut_LC_2_13_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_9_lut_LC_2_13_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_9_lut_LC_2_13_7 (
            .in0(_gnd_net_),
            .in1(N__55437),
            .in2(N__29076),
            .in3(N__22212),
            .lcout(n2694),
            .ltout(),
            .carryin(n12768),
            .carryout(n12769),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_10_lut_LC_2_14_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_10_lut_LC_2_14_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_10_lut_LC_2_14_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_10_lut_LC_2_14_0 (
            .in0(_gnd_net_),
            .in1(N__55426),
            .in2(N__26037),
            .in3(N__22209),
            .lcout(n2693),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(n12770),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_11_lut_LC_2_14_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_11_lut_LC_2_14_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_11_lut_LC_2_14_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_11_lut_LC_2_14_1 (
            .in0(_gnd_net_),
            .in1(N__55433),
            .in2(N__25971),
            .in3(N__22206),
            .lcout(n2692),
            .ltout(),
            .carryin(n12770),
            .carryout(n12771),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_12_lut_LC_2_14_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_12_lut_LC_2_14_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_12_lut_LC_2_14_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_12_lut_LC_2_14_2 (
            .in0(_gnd_net_),
            .in1(N__55427),
            .in2(N__33921),
            .in3(N__22203),
            .lcout(n2691),
            .ltout(),
            .carryin(n12771),
            .carryout(n12772),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_13_lut_LC_2_14_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_13_lut_LC_2_14_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_13_lut_LC_2_14_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_13_lut_LC_2_14_3 (
            .in0(_gnd_net_),
            .in1(N__24128),
            .in2(N__55535),
            .in3(N__22200),
            .lcout(n2690),
            .ltout(),
            .carryin(n12772),
            .carryout(n12773),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_14_lut_LC_2_14_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_14_lut_LC_2_14_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_14_lut_LC_2_14_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_14_lut_LC_2_14_4 (
            .in0(_gnd_net_),
            .in1(N__55431),
            .in2(N__23676),
            .in3(N__22197),
            .lcout(n2689),
            .ltout(),
            .carryin(n12773),
            .carryout(n12774),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_15_lut_LC_2_14_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_15_lut_LC_2_14_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_15_lut_LC_2_14_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_15_lut_LC_2_14_5 (
            .in0(_gnd_net_),
            .in1(N__55434),
            .in2(N__23880),
            .in3(N__22263),
            .lcout(n2688),
            .ltout(),
            .carryin(n12774),
            .carryout(n12775),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_16_lut_LC_2_14_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_16_lut_LC_2_14_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_16_lut_LC_2_14_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_16_lut_LC_2_14_6 (
            .in0(_gnd_net_),
            .in1(N__55432),
            .in2(N__29394),
            .in3(N__22260),
            .lcout(n2687),
            .ltout(),
            .carryin(n12775),
            .carryout(n12776),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_17_lut_LC_2_14_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_17_lut_LC_2_14_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_17_lut_LC_2_14_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_17_lut_LC_2_14_7 (
            .in0(_gnd_net_),
            .in1(N__55435),
            .in2(N__26148),
            .in3(N__22257),
            .lcout(n2686),
            .ltout(),
            .carryin(n12776),
            .carryout(n12777),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_18_lut_LC_2_15_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_18_lut_LC_2_15_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_18_lut_LC_2_15_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_18_lut_LC_2_15_0 (
            .in0(_gnd_net_),
            .in1(N__26235),
            .in2(N__55551),
            .in3(N__22254),
            .lcout(n2685),
            .ltout(),
            .carryin(bfn_2_15_0_),
            .carryout(n12778),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_19_lut_LC_2_15_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_19_lut_LC_2_15_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_19_lut_LC_2_15_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_19_lut_LC_2_15_1 (
            .in0(_gnd_net_),
            .in1(N__25997),
            .in2(N__55555),
            .in3(N__22251),
            .lcout(n2684),
            .ltout(),
            .carryin(n12778),
            .carryout(n12779),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_20_lut_LC_2_15_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_20_lut_LC_2_15_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_20_lut_LC_2_15_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_20_lut_LC_2_15_2 (
            .in0(_gnd_net_),
            .in1(N__32628),
            .in2(N__55552),
            .in3(N__22248),
            .lcout(n2683),
            .ltout(),
            .carryin(n12779),
            .carryout(n12780),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_21_lut_LC_2_15_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_21_lut_LC_2_15_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_21_lut_LC_2_15_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_21_lut_LC_2_15_3 (
            .in0(_gnd_net_),
            .in1(N__29684),
            .in2(N__55556),
            .in3(N__22233),
            .lcout(n2682),
            .ltout(),
            .carryin(n12780),
            .carryout(n12781),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_22_lut_LC_2_15_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_22_lut_LC_2_15_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_22_lut_LC_2_15_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_22_lut_LC_2_15_4 (
            .in0(_gnd_net_),
            .in1(N__26208),
            .in2(N__55553),
            .in3(N__22230),
            .lcout(n2681),
            .ltout(),
            .carryin(n12781),
            .carryout(n12782),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_23_lut_LC_2_15_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_23_lut_LC_2_15_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_23_lut_LC_2_15_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_23_lut_LC_2_15_5 (
            .in0(_gnd_net_),
            .in1(N__26175),
            .in2(N__55557),
            .in3(N__22227),
            .lcout(n2680),
            .ltout(),
            .carryin(n12782),
            .carryout(n12783),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_24_lut_LC_2_15_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_24_lut_LC_2_15_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_24_lut_LC_2_15_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_24_lut_LC_2_15_6 (
            .in0(_gnd_net_),
            .in1(N__29544),
            .in2(N__55554),
            .in3(N__22305),
            .lcout(n2679),
            .ltout(),
            .carryin(n12783),
            .carryout(n12784),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_25_lut_LC_2_15_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1771_25_lut_LC_2_15_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_25_lut_LC_2_15_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_25_lut_LC_2_15_7 (
            .in0(_gnd_net_),
            .in1(N__32559),
            .in2(N__55558),
            .in3(N__22302),
            .lcout(n2678),
            .ltout(),
            .carryin(n12784),
            .carryout(n12785),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1771_26_lut_LC_2_16_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1771_26_lut_LC_2_16_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1771_26_lut_LC_2_16_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1771_26_lut_LC_2_16_0 (
            .in0(_gnd_net_),
            .in1(N__54743),
            .in2(N__32736),
            .in3(N__22299),
            .lcout(n2677),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_2_lut_LC_2_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_2_lut_LC_2_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_2_lut_LC_2_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_2_lut_LC_2_17_0 (
            .in0(_gnd_net_),
            .in1(N__33540),
            .in2(_gnd_net_),
            .in3(N__22281),
            .lcout(n2801),
            .ltout(),
            .carryin(bfn_2_17_0_),
            .carryout(n12786),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_3_lut_LC_2_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_3_lut_LC_2_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_3_lut_LC_2_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_3_lut_LC_2_17_1 (
            .in0(_gnd_net_),
            .in1(N__55493),
            .in2(N__26628),
            .in3(N__22278),
            .lcout(n2800),
            .ltout(),
            .carryin(n12786),
            .carryout(n12787),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_4_lut_LC_2_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_4_lut_LC_2_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_4_lut_LC_2_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_4_lut_LC_2_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24078),
            .in3(N__22275),
            .lcout(n2799),
            .ltout(),
            .carryin(n12787),
            .carryout(n12788),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_5_lut_LC_2_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_5_lut_LC_2_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_5_lut_LC_2_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_5_lut_LC_2_17_3 (
            .in0(_gnd_net_),
            .in1(N__55494),
            .in2(N__24369),
            .in3(N__22272),
            .lcout(n2798),
            .ltout(),
            .carryin(n12788),
            .carryout(n12789),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_6_lut_LC_2_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_6_lut_LC_2_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_6_lut_LC_2_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_6_lut_LC_2_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23838),
            .in3(N__22269),
            .lcout(n2797),
            .ltout(),
            .carryin(n12789),
            .carryout(n12790),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_7_lut_LC_2_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_7_lut_LC_2_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_7_lut_LC_2_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_7_lut_LC_2_17_5 (
            .in0(_gnd_net_),
            .in1(N__23916),
            .in2(_gnd_net_),
            .in3(N__22266),
            .lcout(n2796),
            .ltout(),
            .carryin(n12790),
            .carryout(n12791),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_8_lut_LC_2_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_8_lut_LC_2_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_8_lut_LC_2_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_8_lut_LC_2_17_6 (
            .in0(_gnd_net_),
            .in1(N__55496),
            .in2(N__23733),
            .in3(N__22332),
            .lcout(n2795),
            .ltout(),
            .carryin(n12791),
            .carryout(n12792),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_9_lut_LC_2_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_9_lut_LC_2_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_9_lut_LC_2_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_9_lut_LC_2_17_7 (
            .in0(_gnd_net_),
            .in1(N__55495),
            .in2(N__23562),
            .in3(N__22329),
            .lcout(n2794),
            .ltout(),
            .carryin(n12792),
            .carryout(n12793),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_10_lut_LC_2_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_10_lut_LC_2_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_10_lut_LC_2_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_10_lut_LC_2_18_0 (
            .in0(_gnd_net_),
            .in1(N__55349),
            .in2(N__23715),
            .in3(N__22326),
            .lcout(n2793),
            .ltout(),
            .carryin(bfn_2_18_0_),
            .carryout(n12794),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_11_lut_LC_2_18_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_11_lut_LC_2_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_11_lut_LC_2_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_11_lut_LC_2_18_1 (
            .in0(_gnd_net_),
            .in1(N__55355),
            .in2(N__22698),
            .in3(N__22323),
            .lcout(n2792),
            .ltout(),
            .carryin(n12794),
            .carryout(n12795),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_12_lut_LC_2_18_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_12_lut_LC_2_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_12_lut_LC_2_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_12_lut_LC_2_18_2 (
            .in0(_gnd_net_),
            .in1(N__55350),
            .in2(N__23637),
            .in3(N__22320),
            .lcout(n2791),
            .ltout(),
            .carryin(n12795),
            .carryout(n12796),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_13_lut_LC_2_18_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_13_lut_LC_2_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_13_lut_LC_2_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_13_lut_LC_2_18_3 (
            .in0(_gnd_net_),
            .in1(N__55356),
            .in2(N__22512),
            .in3(N__22317),
            .lcout(n2790),
            .ltout(),
            .carryin(n12796),
            .carryout(n12797),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_14_lut_LC_2_18_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_14_lut_LC_2_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_14_lut_LC_2_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_14_lut_LC_2_18_4 (
            .in0(_gnd_net_),
            .in1(N__55351),
            .in2(N__24102),
            .in3(N__22314),
            .lcout(n2789),
            .ltout(),
            .carryin(n12797),
            .carryout(n12798),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_15_lut_LC_2_18_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_15_lut_LC_2_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_15_lut_LC_2_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_15_lut_LC_2_18_5 (
            .in0(_gnd_net_),
            .in1(N__55357),
            .in2(N__23756),
            .in3(N__22311),
            .lcout(n2788),
            .ltout(),
            .carryin(n12798),
            .carryout(n12799),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_16_lut_LC_2_18_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_16_lut_LC_2_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_16_lut_LC_2_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_16_lut_LC_2_18_6 (
            .in0(_gnd_net_),
            .in1(N__24227),
            .in2(N__55492),
            .in3(N__22308),
            .lcout(n2787),
            .ltout(),
            .carryin(n12799),
            .carryout(n12800),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_17_lut_LC_2_18_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_17_lut_LC_2_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_17_lut_LC_2_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_17_lut_LC_2_18_7 (
            .in0(_gnd_net_),
            .in1(N__23990),
            .in2(N__55491),
            .in3(N__22374),
            .lcout(n2786),
            .ltout(),
            .carryin(n12800),
            .carryout(n12801),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_18_lut_LC_2_19_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_18_lut_LC_2_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_18_lut_LC_2_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_18_lut_LC_2_19_0 (
            .in0(_gnd_net_),
            .in1(N__24165),
            .in2(N__55526),
            .in3(N__22371),
            .lcout(n2785),
            .ltout(),
            .carryin(bfn_2_19_0_),
            .carryout(n12802),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_19_lut_LC_2_19_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_19_lut_LC_2_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_19_lut_LC_2_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_19_lut_LC_2_19_1 (
            .in0(_gnd_net_),
            .in1(N__23952),
            .in2(N__55530),
            .in3(N__22368),
            .lcout(n2784),
            .ltout(),
            .carryin(n12802),
            .carryout(n12803),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_20_lut_LC_2_19_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_20_lut_LC_2_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_20_lut_LC_2_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_20_lut_LC_2_19_2 (
            .in0(_gnd_net_),
            .in1(N__22844),
            .in2(N__55527),
            .in3(N__22350),
            .lcout(n2783),
            .ltout(),
            .carryin(n12803),
            .carryout(n12804),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_21_lut_LC_2_19_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_21_lut_LC_2_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_21_lut_LC_2_19_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_21_lut_LC_2_19_3 (
            .in0(_gnd_net_),
            .in1(N__22582),
            .in2(N__55531),
            .in3(N__22347),
            .lcout(n2782),
            .ltout(),
            .carryin(n12804),
            .carryout(n12805),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_22_lut_LC_2_19_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_22_lut_LC_2_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_22_lut_LC_2_19_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_22_lut_LC_2_19_4 (
            .in0(_gnd_net_),
            .in1(N__24279),
            .in2(N__55528),
            .in3(N__22344),
            .lcout(n2781),
            .ltout(),
            .carryin(n12805),
            .carryout(n12806),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_23_lut_LC_2_19_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_23_lut_LC_2_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_23_lut_LC_2_19_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_23_lut_LC_2_19_5 (
            .in0(_gnd_net_),
            .in1(N__24417),
            .in2(N__55532),
            .in3(N__22341),
            .lcout(n2780),
            .ltout(),
            .carryin(n12806),
            .carryout(n12807),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_24_lut_LC_2_19_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_24_lut_LC_2_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_24_lut_LC_2_19_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_24_lut_LC_2_19_6 (
            .in0(_gnd_net_),
            .in1(N__26106),
            .in2(N__55529),
            .in3(N__22338),
            .lcout(n2779),
            .ltout(),
            .carryin(n12807),
            .carryout(n12808),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_25_lut_LC_2_19_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_25_lut_LC_2_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_25_lut_LC_2_19_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_25_lut_LC_2_19_7 (
            .in0(_gnd_net_),
            .in1(N__24039),
            .in2(N__55533),
            .in3(N__22335),
            .lcout(n2778),
            .ltout(),
            .carryin(n12808),
            .carryout(n12809),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_26_lut_LC_2_20_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1838_26_lut_LC_2_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_26_lut_LC_2_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1838_26_lut_LC_2_20_0 (
            .in0(_gnd_net_),
            .in1(N__24463),
            .in2(N__55547),
            .in3(N__22452),
            .lcout(n2777),
            .ltout(),
            .carryin(bfn_2_20_0_),
            .carryout(n12810),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1838_27_lut_LC_2_20_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1838_27_lut_LC_2_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1838_27_lut_LC_2_20_1.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1838_27_lut_LC_2_20_1 (
            .in0(N__53967),
            .in1(N__22799),
            .in2(N__36491),
            .in3(N__22449),
            .lcout(n2808),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1779_3_lut_LC_2_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1779_3_lut_LC_2_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1779_3_lut_LC_2_20_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1779_3_lut_LC_2_20_4 (
            .in0(_gnd_net_),
            .in1(N__32624),
            .in2(N__36293),
            .in3(N__22446),
            .lcout(n2715),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1773_3_lut_LC_2_20_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1773_3_lut_LC_2_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1773_3_lut_LC_2_20_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1773_3_lut_LC_2_20_5 (
            .in0(_gnd_net_),
            .in1(N__32732),
            .in2(N__22437),
            .in3(N__36275),
            .lcout(n2709),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1774_3_lut_LC_2_20_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1774_3_lut_LC_2_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1774_3_lut_LC_2_20_6.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1774_3_lut_LC_2_20_6 (
            .in0(N__32555),
            .in1(_gnd_net_),
            .in2(N__36294),
            .in3(N__22422),
            .lcout(n2710),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13045_1_lut_LC_2_20_7.C_ON=1'b0;
    defparam i13045_1_lut_LC_2_20_7.SEQ_MODE=4'b0000;
    defparam i13045_1_lut_LC_2_20_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 i13045_1_lut_LC_2_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35744),
            .lcout(n15775),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1861_3_lut_LC_2_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1861_3_lut_LC_2_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1861_3_lut_LC_2_21_0.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1861_3_lut_LC_2_21_0 (
            .in0(_gnd_net_),
            .in1(N__22413),
            .in2(N__36453),
            .in3(N__23831),
            .lcout(n2829),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1790_3_lut_LC_2_21_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1790_3_lut_LC_2_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1790_3_lut_LC_2_21_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1790_3_lut_LC_2_21_1 (
            .in0(_gnd_net_),
            .in1(N__29069),
            .in2(N__22404),
            .in3(N__36262),
            .lcout(n2726),
            .ltout(n2726_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1857_3_lut_LC_2_21_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1857_3_lut_LC_2_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1857_3_lut_LC_2_21_2.LUT_INIT=16'b1110010011100100;
    LogicCell40 encoder0_position_31__I_0_i1857_3_lut_LC_2_21_2 (
            .in0(N__36422),
            .in1(N__22389),
            .in2(N__22377),
            .in3(_gnd_net_),
            .lcout(n2825),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1717_3_lut_LC_2_21_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1717_3_lut_LC_2_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1717_3_lut_LC_2_21_3.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1717_3_lut_LC_2_21_3 (
            .in0(N__34086),
            .in1(_gnd_net_),
            .in2(N__32484),
            .in3(N__36095),
            .lcout(n2621),
            .ltout(n2621_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1784_3_lut_LC_2_21_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1784_3_lut_LC_2_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1784_3_lut_LC_2_21_4.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1784_3_lut_LC_2_21_4 (
            .in0(N__36266),
            .in1(_gnd_net_),
            .in2(N__22566),
            .in3(N__22563),
            .lcout(n2720),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1792_3_lut_LC_2_21_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1792_3_lut_LC_2_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1792_3_lut_LC_2_21_6.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1792_3_lut_LC_2_21_6 (
            .in0(_gnd_net_),
            .in1(N__29501),
            .in2(N__36292),
            .in3(N__22551),
            .lcout(n2728),
            .ltout(n2728_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1859_3_lut_LC_2_21_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1859_3_lut_LC_2_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1859_3_lut_LC_2_21_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1859_3_lut_LC_2_21_7 (
            .in0(_gnd_net_),
            .in1(N__22536),
            .in2(N__22527),
            .in3(N__36418),
            .lcout(n2827),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_54_LC_2_22_0.C_ON=1'b0;
    defparam i1_4_lut_adj_54_LC_2_22_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_54_LC_2_22_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_54_LC_2_22_0 (
            .in0(N__22502),
            .in1(N__23551),
            .in2(N__22690),
            .in3(N__24220),
            .lcout(n14346),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1787_3_lut_LC_2_22_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1787_3_lut_LC_2_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1787_3_lut_LC_2_22_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1787_3_lut_LC_2_22_1 (
            .in0(_gnd_net_),
            .in1(N__33917),
            .in2(N__22524),
            .in3(N__36234),
            .lcout(n2723),
            .ltout(n2723_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1854_3_lut_LC_2_22_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1854_3_lut_LC_2_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1854_3_lut_LC_2_22_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1854_3_lut_LC_2_22_2 (
            .in0(_gnd_net_),
            .in1(N__22491),
            .in2(N__22479),
            .in3(N__36423),
            .lcout(n2822),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1789_3_lut_LC_2_22_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1789_3_lut_LC_2_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1789_3_lut_LC_2_22_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1789_3_lut_LC_2_22_3 (
            .in0(_gnd_net_),
            .in1(N__22476),
            .in2(N__26033),
            .in3(N__36235),
            .lcout(n2725),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1793_3_lut_LC_2_22_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1793_3_lut_LC_2_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1793_3_lut_LC_2_22_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1793_3_lut_LC_2_22_4 (
            .in0(_gnd_net_),
            .in1(N__29434),
            .in2(N__36279),
            .in3(N__22467),
            .lcout(n2729),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1777_3_lut_LC_2_22_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1777_3_lut_LC_2_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1777_3_lut_LC_2_22_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1777_3_lut_LC_2_22_5 (
            .in0(_gnd_net_),
            .in1(N__26207),
            .in2(N__22665),
            .in3(N__36239),
            .lcout(n2713),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1858_3_lut_LC_2_22_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1858_3_lut_LC_2_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1858_3_lut_LC_2_22_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1858_3_lut_LC_2_22_6 (
            .in0(_gnd_net_),
            .in1(N__23552),
            .in2(N__22650),
            .in3(N__36424),
            .lcout(n2826),
            .ltout(n2826_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_61_LC_2_22_7.C_ON=1'b0;
    defparam i1_4_lut_adj_61_LC_2_22_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_61_LC_2_22_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_61_LC_2_22_7 (
            .in0(N__22756),
            .in1(N__24577),
            .in2(N__22635),
            .in3(N__24535),
            .lcout(n14688),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_59_LC_2_23_0.C_ON=1'b0;
    defparam i1_4_lut_adj_59_LC_2_23_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_59_LC_2_23_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_59_LC_2_23_0 (
            .in0(N__23886),
            .in1(N__22583),
            .in2(N__22843),
            .in3(N__22605),
            .lcout(),
            .ltout(n14362_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_60_LC_2_23_1.C_ON=1'b0;
    defparam i1_4_lut_adj_60_LC_2_23_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_60_LC_2_23_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_60_LC_2_23_1 (
            .in0(N__24278),
            .in1(N__26098),
            .in2(N__22632),
            .in3(N__24415),
            .lcout(n14368),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1853_3_lut_LC_2_23_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1853_3_lut_LC_2_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1853_3_lut_LC_2_23_2.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1853_3_lut_LC_2_23_2 (
            .in0(_gnd_net_),
            .in1(N__24092),
            .in2(N__36445),
            .in3(N__22629),
            .lcout(n2821),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_56_LC_2_23_3.C_ON=1'b0;
    defparam i1_3_lut_adj_56_LC_2_23_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_56_LC_2_23_3.LUT_INIT=16'b1111111111111010;
    LogicCell40 i1_3_lut_adj_56_LC_2_23_3 (
            .in0(N__24091),
            .in1(_gnd_net_),
            .in2(N__22617),
            .in3(N__23983),
            .lcout(),
            .ltout(n14350_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_57_LC_2_23_4.C_ON=1'b0;
    defparam i1_4_lut_adj_57_LC_2_23_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_57_LC_2_23_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_57_LC_2_23_4 (
            .in0(N__23694),
            .in1(N__24157),
            .in2(N__22608),
            .in3(N__23945),
            .lcout(n14356),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1846_3_lut_LC_2_23_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1846_3_lut_LC_2_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1846_3_lut_LC_2_23_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1846_3_lut_LC_2_23_5 (
            .in0(_gnd_net_),
            .in1(N__22599),
            .in2(N__22587),
            .in3(N__36408),
            .lcout(n2814),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1849_3_lut_LC_2_23_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1849_3_lut_LC_2_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1849_3_lut_LC_2_23_6.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1849_3_lut_LC_2_23_6 (
            .in0(_gnd_net_),
            .in1(N__24158),
            .in2(N__36446),
            .in3(N__22872),
            .lcout(n2817),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1780_3_lut_LC_2_23_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1780_3_lut_LC_2_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1780_3_lut_LC_2_23_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1780_3_lut_LC_2_23_7 (
            .in0(_gnd_net_),
            .in1(N__22860),
            .in2(N__25998),
            .in3(N__36258),
            .lcout(n2716),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1775_3_lut_LC_2_24_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1775_3_lut_LC_2_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1775_3_lut_LC_2_24_0.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1775_3_lut_LC_2_24_0 (
            .in0(N__29540),
            .in1(_gnd_net_),
            .in2(N__22818),
            .in3(N__36245),
            .lcout(n2711),
            .ltout(n2711_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12595_4_lut_LC_2_24_1.C_ON=1'b0;
    defparam i12595_4_lut_LC_2_24_1.SEQ_MODE=4'b0000;
    defparam i12595_4_lut_LC_2_24_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12595_4_lut_LC_2_24_1 (
            .in0(N__22800),
            .in1(N__24467),
            .in2(N__22785),
            .in3(N__22782),
            .lcout(n2742),
            .ltout(n2742_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1860_3_lut_LC_2_24_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1860_3_lut_LC_2_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1860_3_lut_LC_2_24_2.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1860_3_lut_LC_2_24_2 (
            .in0(_gnd_net_),
            .in1(N__22776),
            .in2(N__22764),
            .in3(N__23915),
            .lcout(n2828),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12592_1_lut_LC_2_24_3.C_ON=1'b0;
    defparam i12592_1_lut_LC_2_24_3.SEQ_MODE=4'b0000;
    defparam i12592_1_lut_LC_2_24_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12592_1_lut_LC_2_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36437),
            .lcout(n15322),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1852_3_lut_LC_2_24_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1852_3_lut_LC_2_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1852_3_lut_LC_2_24_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1852_3_lut_LC_2_24_4 (
            .in0(_gnd_net_),
            .in1(N__23757),
            .in2(N__36457),
            .in3(N__22731),
            .lcout(n2820),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1783_3_lut_LC_2_24_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1783_3_lut_LC_2_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1783_3_lut_LC_2_24_5.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1783_3_lut_LC_2_24_5 (
            .in0(_gnd_net_),
            .in1(N__29387),
            .in2(N__36280),
            .in3(N__22719),
            .lcout(n2719),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1856_3_lut_LC_2_24_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1856_3_lut_LC_2_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1856_3_lut_LC_2_24_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1856_3_lut_LC_2_24_6 (
            .in0(_gnd_net_),
            .in1(N__22707),
            .in2(N__36456),
            .in3(N__22694),
            .lcout(n2824),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1855_3_lut_LC_2_24_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1855_3_lut_LC_2_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1855_3_lut_LC_2_24_7.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1855_3_lut_LC_2_24_7 (
            .in0(N__22911),
            .in1(_gnd_net_),
            .in2(N__23636),
            .in3(N__36438),
            .lcout(n2823),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_2_lut_LC_2_25_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_2_lut_LC_2_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_2_lut_LC_2_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_2_lut_LC_2_25_0 (
            .in0(_gnd_net_),
            .in1(N__35178),
            .in2(_gnd_net_),
            .in3(N__22902),
            .lcout(n3001),
            .ltout(),
            .carryin(bfn_2_25_0_),
            .carryout(n12837),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_3_lut_LC_2_25_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_3_lut_LC_2_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_3_lut_LC_2_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_3_lut_LC_2_25_1 (
            .in0(_gnd_net_),
            .in1(N__30222),
            .in2(N__55083),
            .in3(N__22899),
            .lcout(n3000),
            .ltout(),
            .carryin(n12837),
            .carryout(n12838),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_4_lut_LC_2_25_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_4_lut_LC_2_25_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_4_lut_LC_2_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_4_lut_LC_2_25_2 (
            .in0(_gnd_net_),
            .in1(N__30130),
            .in2(_gnd_net_),
            .in3(N__22896),
            .lcout(n2999),
            .ltout(),
            .carryin(n12838),
            .carryout(n12839),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_5_lut_LC_2_25_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_5_lut_LC_2_25_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_5_lut_LC_2_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_5_lut_LC_2_25_3 (
            .in0(_gnd_net_),
            .in1(N__30007),
            .in2(N__55084),
            .in3(N__22893),
            .lcout(n2998),
            .ltout(),
            .carryin(n12839),
            .carryout(n12840),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_6_lut_LC_2_25_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_6_lut_LC_2_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_6_lut_LC_2_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_6_lut_LC_2_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29598),
            .in3(N__22890),
            .lcout(n2997),
            .ltout(),
            .carryin(n12840),
            .carryout(n12841),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_7_lut_LC_2_25_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_7_lut_LC_2_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_7_lut_LC_2_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_7_lut_LC_2_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27167),
            .in3(N__22887),
            .lcout(n2996),
            .ltout(),
            .carryin(n12841),
            .carryout(n12842),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_8_lut_LC_2_25_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_8_lut_LC_2_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_8_lut_LC_2_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_8_lut_LC_2_25_6 (
            .in0(_gnd_net_),
            .in1(N__29856),
            .in2(N__55066),
            .in3(N__22884),
            .lcout(n2995),
            .ltout(),
            .carryin(n12842),
            .carryout(n12843),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_9_lut_LC_2_25_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_9_lut_LC_2_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_9_lut_LC_2_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_9_lut_LC_2_25_7 (
            .in0(_gnd_net_),
            .in1(N__26795),
            .in2(N__55085),
            .in3(N__22875),
            .lcout(n2994),
            .ltout(),
            .carryin(n12843),
            .carryout(n12844),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_10_lut_LC_2_26_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_10_lut_LC_2_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_10_lut_LC_2_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_10_lut_LC_2_26_0 (
            .in0(_gnd_net_),
            .in1(N__26774),
            .in2(N__55062),
            .in3(N__22956),
            .lcout(n2993),
            .ltout(),
            .carryin(bfn_2_26_0_),
            .carryout(n12845),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_11_lut_LC_2_26_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_11_lut_LC_2_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_11_lut_LC_2_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_11_lut_LC_2_26_1 (
            .in0(_gnd_net_),
            .in1(N__29708),
            .in2(N__55080),
            .in3(N__22947),
            .lcout(n2992),
            .ltout(),
            .carryin(n12845),
            .carryout(n12846),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_12_lut_LC_2_26_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_12_lut_LC_2_26_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_12_lut_LC_2_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_12_lut_LC_2_26_2 (
            .in0(_gnd_net_),
            .in1(N__29562),
            .in2(N__55063),
            .in3(N__22944),
            .lcout(n2991),
            .ltout(),
            .carryin(n12846),
            .carryout(n12847),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_13_lut_LC_2_26_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_13_lut_LC_2_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_13_lut_LC_2_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_13_lut_LC_2_26_3 (
            .in0(_gnd_net_),
            .in1(N__54813),
            .in2(N__29300),
            .in3(N__22932),
            .lcout(n2990),
            .ltout(),
            .carryin(n12847),
            .carryout(n12848),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_14_lut_LC_2_26_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_14_lut_LC_2_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_14_lut_LC_2_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_14_lut_LC_2_26_4 (
            .in0(_gnd_net_),
            .in1(N__26675),
            .in2(N__55064),
            .in3(N__22923),
            .lcout(n2989),
            .ltout(),
            .carryin(n12848),
            .carryout(n12849),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_15_lut_LC_2_26_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_15_lut_LC_2_26_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_15_lut_LC_2_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_15_lut_LC_2_26_5 (
            .in0(_gnd_net_),
            .in1(N__26699),
            .in2(N__55081),
            .in3(N__22920),
            .lcout(n2988),
            .ltout(),
            .carryin(n12849),
            .carryout(n12850),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_16_lut_LC_2_26_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_16_lut_LC_2_26_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_16_lut_LC_2_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_16_lut_LC_2_26_6 (
            .in0(_gnd_net_),
            .in1(N__30179),
            .in2(N__55065),
            .in3(N__22917),
            .lcout(n2987),
            .ltout(),
            .carryin(n12850),
            .carryout(n12851),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_17_lut_LC_2_26_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_17_lut_LC_2_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_17_lut_LC_2_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_17_lut_LC_2_26_7 (
            .in0(_gnd_net_),
            .in1(N__26654),
            .in2(N__55082),
            .in3(N__22914),
            .lcout(n2986),
            .ltout(),
            .carryin(n12851),
            .carryout(n12852),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_18_lut_LC_2_27_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_18_lut_LC_2_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_18_lut_LC_2_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_18_lut_LC_2_27_0 (
            .in0(_gnd_net_),
            .in1(N__26813),
            .in2(N__55058),
            .in3(N__22998),
            .lcout(n2985),
            .ltout(),
            .carryin(bfn_2_27_0_),
            .carryout(n12853),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_19_lut_LC_2_27_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_19_lut_LC_2_27_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_19_lut_LC_2_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_19_lut_LC_2_27_1 (
            .in0(_gnd_net_),
            .in1(N__30368),
            .in2(N__55076),
            .in3(N__22995),
            .lcout(n2984),
            .ltout(),
            .carryin(n12853),
            .carryout(n12854),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_20_lut_LC_2_27_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_20_lut_LC_2_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_20_lut_LC_2_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_20_lut_LC_2_27_2 (
            .in0(_gnd_net_),
            .in1(N__27204),
            .in2(N__55059),
            .in3(N__22992),
            .lcout(n2983),
            .ltout(),
            .carryin(n12854),
            .carryout(n12855),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_21_lut_LC_2_27_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_21_lut_LC_2_27_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_21_lut_LC_2_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_21_lut_LC_2_27_3 (
            .in0(_gnd_net_),
            .in1(N__27123),
            .in2(N__55077),
            .in3(N__22989),
            .lcout(n2982),
            .ltout(),
            .carryin(n12855),
            .carryout(n12856),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_22_lut_LC_2_27_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_22_lut_LC_2_27_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_22_lut_LC_2_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_22_lut_LC_2_27_4 (
            .in0(_gnd_net_),
            .in1(N__27093),
            .in2(N__55060),
            .in3(N__22986),
            .lcout(n2981),
            .ltout(),
            .carryin(n12856),
            .carryout(n12857),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_23_lut_LC_2_27_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_23_lut_LC_2_27_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_23_lut_LC_2_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_23_lut_LC_2_27_5 (
            .in0(_gnd_net_),
            .in1(N__30294),
            .in2(N__55078),
            .in3(N__22983),
            .lcout(n2980),
            .ltout(),
            .carryin(n12857),
            .carryout(n12858),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_24_lut_LC_2_27_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_24_lut_LC_2_27_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_24_lut_LC_2_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_24_lut_LC_2_27_6 (
            .in0(_gnd_net_),
            .in1(N__27042),
            .in2(N__55061),
            .in3(N__22980),
            .lcout(n2979),
            .ltout(),
            .carryin(n12858),
            .carryout(n12859),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_25_lut_LC_2_27_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_25_lut_LC_2_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_25_lut_LC_2_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_25_lut_LC_2_27_7 (
            .in0(_gnd_net_),
            .in1(N__26937),
            .in2(N__55079),
            .in3(N__22977),
            .lcout(n2978),
            .ltout(),
            .carryin(n12859),
            .carryout(n12860),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_26_lut_LC_2_28_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_26_lut_LC_2_28_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_26_lut_LC_2_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_26_lut_LC_2_28_0 (
            .in0(_gnd_net_),
            .in1(N__27071),
            .in2(N__55057),
            .in3(N__22965),
            .lcout(n2977),
            .ltout(),
            .carryin(bfn_2_28_0_),
            .carryout(n12861),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_27_lut_LC_2_28_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_27_lut_LC_2_28_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_27_lut_LC_2_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_27_lut_LC_2_28_1 (
            .in0(_gnd_net_),
            .in1(N__54792),
            .in2(N__26979),
            .in3(N__23031),
            .lcout(n2976),
            .ltout(),
            .carryin(n12861),
            .carryout(n12862),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_28_lut_LC_2_28_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1972_28_lut_LC_2_28_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_28_lut_LC_2_28_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1972_28_lut_LC_2_28_2 (
            .in0(_gnd_net_),
            .in1(N__54793),
            .in2(N__27030),
            .in3(N__23019),
            .lcout(n2975),
            .ltout(),
            .carryin(n12862),
            .carryout(n12863),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1972_29_lut_LC_2_28_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1972_29_lut_LC_2_28_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1972_29_lut_LC_2_28_3.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1972_29_lut_LC_2_28_3 (
            .in0(N__54794),
            .in1(N__27002),
            .in2(N__34532),
            .in3(N__23016),
            .lcout(n3006),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2061_3_lut_LC_2_28_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2061_3_lut_LC_2_28_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2061_3_lut_LC_2_28_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2061_3_lut_LC_2_28_4 (
            .in0(_gnd_net_),
            .in1(N__24788),
            .in2(N__24762),
            .in3(N__34649),
            .lcout(n3125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2055_3_lut_LC_2_28_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2055_3_lut_LC_2_28_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2055_3_lut_LC_2_28_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2055_3_lut_LC_2_28_5 (
            .in0(_gnd_net_),
            .in1(N__24912),
            .in2(N__34695),
            .in3(N__24934),
            .lcout(n3119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2057_3_lut_LC_2_28_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2057_3_lut_LC_2_28_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2057_3_lut_LC_2_28_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2057_3_lut_LC_2_28_6 (
            .in0(_gnd_net_),
            .in1(N__25010),
            .in2(N__24990),
            .in3(N__34653),
            .lcout(n3121),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2052_3_lut_LC_2_28_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2052_3_lut_LC_2_28_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2052_3_lut_LC_2_28_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2052_3_lut_LC_2_28_7 (
            .in0(_gnd_net_),
            .in1(N__24864),
            .in2(N__34696),
            .in3(N__24884),
            .lcout(n3116),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_2_lut_LC_2_29_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_2_lut_LC_2_29_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_2_lut_LC_2_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_2_lut_LC_2_29_0 (
            .in0(_gnd_net_),
            .in1(N__34170),
            .in2(_gnd_net_),
            .in3(N__23013),
            .lcout(n3201),
            .ltout(),
            .carryin(bfn_2_29_0_),
            .carryout(n12892),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_3_lut_LC_2_29_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_3_lut_LC_2_29_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_3_lut_LC_2_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_3_lut_LC_2_29_1 (
            .in0(_gnd_net_),
            .in1(N__54572),
            .in2(N__30432),
            .in3(N__23010),
            .lcout(n3200),
            .ltout(),
            .carryin(n12892),
            .carryout(n12893),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_4_lut_LC_2_29_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_4_lut_LC_2_29_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_4_lut_LC_2_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_4_lut_LC_2_29_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30510),
            .in3(N__23007),
            .lcout(n3199),
            .ltout(),
            .carryin(n12893),
            .carryout(n12894),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_5_lut_LC_2_29_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_5_lut_LC_2_29_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_5_lut_LC_2_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_5_lut_LC_2_29_3 (
            .in0(_gnd_net_),
            .in1(N__54573),
            .in2(N__30396),
            .in3(N__23058),
            .lcout(n3198),
            .ltout(),
            .carryin(n12894),
            .carryout(n12895),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_6_lut_LC_2_29_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_6_lut_LC_2_29_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_6_lut_LC_2_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_6_lut_LC_2_29_4 (
            .in0(_gnd_net_),
            .in1(N__32957),
            .in2(_gnd_net_),
            .in3(N__23055),
            .lcout(n3197),
            .ltout(),
            .carryin(n12895),
            .carryout(n12896),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_7_lut_LC_2_29_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_7_lut_LC_2_29_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_7_lut_LC_2_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_7_lut_LC_2_29_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30492),
            .in3(N__23052),
            .lcout(n3196),
            .ltout(),
            .carryin(n12896),
            .carryout(n12897),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_8_lut_LC_2_29_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_8_lut_LC_2_29_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_8_lut_LC_2_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_8_lut_LC_2_29_6 (
            .in0(_gnd_net_),
            .in1(N__54582),
            .in2(N__28007),
            .in3(N__23049),
            .lcout(n3195),
            .ltout(),
            .carryin(n12897),
            .carryout(n12898),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_9_lut_LC_2_29_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_9_lut_LC_2_29_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_9_lut_LC_2_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_9_lut_LC_2_29_7 (
            .in0(_gnd_net_),
            .in1(N__27733),
            .in2(N__54879),
            .in3(N__23046),
            .lcout(n3194),
            .ltout(),
            .carryin(n12898),
            .carryout(n12899),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_10_lut_LC_2_30_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_10_lut_LC_2_30_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_10_lut_LC_2_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_10_lut_LC_2_30_0 (
            .in0(_gnd_net_),
            .in1(N__54556),
            .in2(N__32916),
            .in3(N__23043),
            .lcout(n3193),
            .ltout(),
            .carryin(bfn_2_30_0_),
            .carryout(n12900),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_11_lut_LC_2_30_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_11_lut_LC_2_30_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_11_lut_LC_2_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_11_lut_LC_2_30_1 (
            .in0(_gnd_net_),
            .in1(N__54564),
            .in2(N__27764),
            .in3(N__23040),
            .lcout(n3192),
            .ltout(),
            .carryin(n12900),
            .carryout(n12901),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_12_lut_LC_2_30_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_12_lut_LC_2_30_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_12_lut_LC_2_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_12_lut_LC_2_30_2 (
            .in0(_gnd_net_),
            .in1(N__54557),
            .in2(N__30812),
            .in3(N__23037),
            .lcout(n3191),
            .ltout(),
            .carryin(n12901),
            .carryout(n12902),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_13_lut_LC_2_30_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_13_lut_LC_2_30_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_13_lut_LC_2_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_13_lut_LC_2_30_3 (
            .in0(_gnd_net_),
            .in1(N__54565),
            .in2(N__27551),
            .in3(N__23034),
            .lcout(n3190),
            .ltout(),
            .carryin(n12902),
            .carryout(n12903),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_14_lut_LC_2_30_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_14_lut_LC_2_30_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_14_lut_LC_2_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_14_lut_LC_2_30_4 (
            .in0(_gnd_net_),
            .in1(N__30692),
            .in2(N__54877),
            .in3(N__23103),
            .lcout(n3189),
            .ltout(),
            .carryin(n12903),
            .carryout(n12904),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_15_lut_LC_2_30_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_15_lut_LC_2_30_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_15_lut_LC_2_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_15_lut_LC_2_30_5 (
            .in0(_gnd_net_),
            .in1(N__27809),
            .in2(N__54875),
            .in3(N__23100),
            .lcout(n3188),
            .ltout(),
            .carryin(n12904),
            .carryout(n12905),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_16_lut_LC_2_30_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_16_lut_LC_2_30_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_16_lut_LC_2_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_16_lut_LC_2_30_6 (
            .in0(_gnd_net_),
            .in1(N__23097),
            .in2(N__54878),
            .in3(N__23079),
            .lcout(n3187),
            .ltout(),
            .carryin(n12905),
            .carryout(n12906),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_17_lut_LC_2_30_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_17_lut_LC_2_30_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_17_lut_LC_2_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_17_lut_LC_2_30_7 (
            .in0(_gnd_net_),
            .in1(N__27683),
            .in2(N__54876),
            .in3(N__23076),
            .lcout(n3186),
            .ltout(),
            .carryin(n12906),
            .carryout(n12907),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_18_lut_LC_2_31_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_18_lut_LC_2_31_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_18_lut_LC_2_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_18_lut_LC_2_31_0 (
            .in0(_gnd_net_),
            .in1(N__30890),
            .in2(N__54871),
            .in3(N__23073),
            .lcout(n3185),
            .ltout(),
            .carryin(bfn_2_31_0_),
            .carryout(n12908),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_19_lut_LC_2_31_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_19_lut_LC_2_31_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_19_lut_LC_2_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_19_lut_LC_2_31_1 (
            .in0(_gnd_net_),
            .in1(N__27969),
            .in2(N__54726),
            .in3(N__23070),
            .lcout(n3184),
            .ltout(),
            .carryin(n12908),
            .carryout(n12909),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_20_lut_LC_2_31_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_20_lut_LC_2_31_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_20_lut_LC_2_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_20_lut_LC_2_31_2 (
            .in0(_gnd_net_),
            .in1(N__30665),
            .in2(N__54872),
            .in3(N__23067),
            .lcout(n3183),
            .ltout(),
            .carryin(n12909),
            .carryout(n12910),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_21_lut_LC_2_31_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_21_lut_LC_2_31_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_21_lut_LC_2_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_21_lut_LC_2_31_3 (
            .in0(_gnd_net_),
            .in1(N__30038),
            .in2(N__54727),
            .in3(N__23064),
            .lcout(n3182),
            .ltout(),
            .carryin(n12910),
            .carryout(n12911),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_22_lut_LC_2_31_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_22_lut_LC_2_31_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_22_lut_LC_2_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_22_lut_LC_2_31_4 (
            .in0(_gnd_net_),
            .in1(N__27914),
            .in2(N__54873),
            .in3(N__23061),
            .lcout(n3181),
            .ltout(),
            .carryin(n12911),
            .carryout(n12912),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_23_lut_LC_2_31_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_23_lut_LC_2_31_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_23_lut_LC_2_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_23_lut_LC_2_31_5 (
            .in0(_gnd_net_),
            .in1(N__27882),
            .in2(N__54728),
            .in3(N__23130),
            .lcout(n3180),
            .ltout(),
            .carryin(n12912),
            .carryout(n12913),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_24_lut_LC_2_31_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_24_lut_LC_2_31_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_24_lut_LC_2_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_24_lut_LC_2_31_6 (
            .in0(_gnd_net_),
            .in1(N__30738),
            .in2(N__54874),
            .in3(N__23127),
            .lcout(n3179),
            .ltout(),
            .carryin(n12913),
            .carryout(n12914),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_25_lut_LC_2_31_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_25_lut_LC_2_31_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_25_lut_LC_2_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_25_lut_LC_2_31_7 (
            .in0(_gnd_net_),
            .in1(N__31064),
            .in2(N__54729),
            .in3(N__23124),
            .lcout(n3178),
            .ltout(),
            .carryin(n12914),
            .carryout(n12915),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_26_lut_LC_2_32_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_26_lut_LC_2_32_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_26_lut_LC_2_32_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_26_lut_LC_2_32_0 (
            .in0(_gnd_net_),
            .in1(N__31028),
            .in2(N__54325),
            .in3(N__23121),
            .lcout(n3177),
            .ltout(),
            .carryin(bfn_2_32_0_),
            .carryout(n12916),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_27_lut_LC_2_32_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_27_lut_LC_2_32_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_27_lut_LC_2_32_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_27_lut_LC_2_32_1 (
            .in0(_gnd_net_),
            .in1(N__30852),
            .in2(N__54328),
            .in3(N__23118),
            .lcout(n3176),
            .ltout(),
            .carryin(n12916),
            .carryout(n12917),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_28_lut_LC_2_32_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_28_lut_LC_2_32_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_28_lut_LC_2_32_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_28_lut_LC_2_32_2 (
            .in0(_gnd_net_),
            .in1(N__27843),
            .in2(N__54326),
            .in3(N__23115),
            .lcout(n3175),
            .ltout(),
            .carryin(n12917),
            .carryout(n12918),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_29_lut_LC_2_32_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_29_lut_LC_2_32_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_29_lut_LC_2_32_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_29_lut_LC_2_32_3 (
            .in0(_gnd_net_),
            .in1(N__28076),
            .in2(N__54329),
            .in3(N__23112),
            .lcout(n3174),
            .ltout(),
            .carryin(n12918),
            .carryout(n12919),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_30_lut_LC_2_32_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2106_30_lut_LC_2_32_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_30_lut_LC_2_32_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2106_30_lut_LC_2_32_4 (
            .in0(_gnd_net_),
            .in1(N__28058),
            .in2(N__54327),
            .in3(N__23109),
            .lcout(n3173),
            .ltout(),
            .carryin(n12919),
            .carryout(n12920),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2106_31_lut_LC_2_32_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_2106_31_lut_LC_2_32_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2106_31_lut_LC_2_32_5.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_2106_31_lut_LC_2_32_5 (
            .in0(N__53935),
            .in1(N__28040),
            .in2(N__34940),
            .in3(N__23106),
            .lcout(n3204),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_2_lut_LC_3_14_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_2_lut_LC_3_14_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_2_lut_LC_3_14_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_2_lut_LC_3_14_0 (
            .in0(_gnd_net_),
            .in1(N__38206),
            .in2(_gnd_net_),
            .in3(N__23157),
            .lcout(n2301),
            .ltout(),
            .carryin(bfn_3_14_0_),
            .carryout(n12676),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_3_lut_LC_3_14_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_3_lut_LC_3_14_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_3_lut_LC_3_14_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_3_lut_LC_3_14_1 (
            .in0(_gnd_net_),
            .in1(N__55543),
            .in2(N__23238),
            .in3(N__23154),
            .lcout(n2300),
            .ltout(),
            .carryin(n12676),
            .carryout(n12677),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_4_lut_LC_3_14_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_4_lut_LC_3_14_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_4_lut_LC_3_14_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_4_lut_LC_3_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25235),
            .in3(N__23151),
            .lcout(n2299),
            .ltout(),
            .carryin(n12677),
            .carryout(n12678),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_5_lut_LC_3_14_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_5_lut_LC_3_14_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_5_lut_LC_3_14_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_5_lut_LC_3_14_3 (
            .in0(_gnd_net_),
            .in1(N__55544),
            .in2(N__25208),
            .in3(N__23148),
            .lcout(n2298),
            .ltout(),
            .carryin(n12678),
            .carryout(n12679),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_6_lut_LC_3_14_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_6_lut_LC_3_14_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_6_lut_LC_3_14_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_6_lut_LC_3_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28386),
            .in3(N__23145),
            .lcout(n2297),
            .ltout(),
            .carryin(n12679),
            .carryout(n12680),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_7_lut_LC_3_14_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_7_lut_LC_3_14_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_7_lut_LC_3_14_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_7_lut_LC_3_14_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25152),
            .in3(N__23142),
            .lcout(n2296),
            .ltout(),
            .carryin(n12680),
            .carryout(n12681),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_8_lut_LC_3_14_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_8_lut_LC_3_14_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_8_lut_LC_3_14_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_8_lut_LC_3_14_6 (
            .in0(_gnd_net_),
            .in1(N__55546),
            .in2(N__25400),
            .in3(N__23139),
            .lcout(n2295),
            .ltout(),
            .carryin(n12681),
            .carryout(n12682),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_9_lut_LC_3_14_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_9_lut_LC_3_14_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_9_lut_LC_3_14_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_9_lut_LC_3_14_7 (
            .in0(_gnd_net_),
            .in1(N__55545),
            .in2(N__28254),
            .in3(N__23136),
            .lcout(n2294),
            .ltout(),
            .carryin(n12682),
            .carryout(n12683),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_10_lut_LC_3_15_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_10_lut_LC_3_15_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_10_lut_LC_3_15_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_10_lut_LC_3_15_0 (
            .in0(_gnd_net_),
            .in1(N__55540),
            .in2(N__25376),
            .in3(N__23133),
            .lcout(n2293),
            .ltout(),
            .carryin(bfn_3_15_0_),
            .carryout(n12684),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_11_lut_LC_3_15_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_11_lut_LC_3_15_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_11_lut_LC_3_15_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_11_lut_LC_3_15_1 (
            .in0(_gnd_net_),
            .in1(N__55419),
            .in2(N__25349),
            .in3(N__23184),
            .lcout(n2292),
            .ltout(),
            .carryin(n12684),
            .carryout(n12685),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_12_lut_LC_3_15_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_12_lut_LC_3_15_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_12_lut_LC_3_15_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_12_lut_LC_3_15_2 (
            .in0(_gnd_net_),
            .in1(N__55541),
            .in2(N__28305),
            .in3(N__23181),
            .lcout(n2291),
            .ltout(),
            .carryin(n12685),
            .carryout(n12686),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_13_lut_LC_3_15_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_13_lut_LC_3_15_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_13_lut_LC_3_15_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_13_lut_LC_3_15_3 (
            .in0(_gnd_net_),
            .in1(N__55420),
            .in2(N__28341),
            .in3(N__23178),
            .lcout(n2290),
            .ltout(),
            .carryin(n12686),
            .carryout(n12687),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_14_lut_LC_3_15_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_14_lut_LC_3_15_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_14_lut_LC_3_15_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_14_lut_LC_3_15_4 (
            .in0(_gnd_net_),
            .in1(N__55542),
            .in2(N__23310),
            .in3(N__23175),
            .lcout(n2289),
            .ltout(),
            .carryin(n12687),
            .carryout(n12688),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_15_lut_LC_3_15_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_15_lut_LC_3_15_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_15_lut_LC_3_15_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_15_lut_LC_3_15_5 (
            .in0(_gnd_net_),
            .in1(N__55421),
            .in2(N__25178),
            .in3(N__23172),
            .lcout(n2288),
            .ltout(),
            .carryin(n12688),
            .carryout(n12689),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_16_lut_LC_3_15_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_16_lut_LC_3_15_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_16_lut_LC_3_15_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_16_lut_LC_3_15_6 (
            .in0(_gnd_net_),
            .in1(N__25494),
            .in2(N__55534),
            .in3(N__23169),
            .lcout(n2287),
            .ltout(),
            .carryin(n12689),
            .carryout(n12690),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_17_lut_LC_3_15_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_17_lut_LC_3_15_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_17_lut_LC_3_15_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_17_lut_LC_3_15_7 (
            .in0(_gnd_net_),
            .in1(N__55425),
            .in2(N__23349),
            .in3(N__23166),
            .lcout(n2286),
            .ltout(),
            .carryin(n12690),
            .carryout(n12691),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_18_lut_LC_3_16_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_18_lut_LC_3_16_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_18_lut_LC_3_16_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_18_lut_LC_3_16_0 (
            .in0(_gnd_net_),
            .in1(N__54732),
            .in2(N__25539),
            .in3(N__23163),
            .lcout(n2285),
            .ltout(),
            .carryin(bfn_3_16_0_),
            .carryout(n12692),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_19_lut_LC_3_16_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_19_lut_LC_3_16_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_19_lut_LC_3_16_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_19_lut_LC_3_16_1 (
            .in0(_gnd_net_),
            .in1(N__54736),
            .in2(N__28539),
            .in3(N__23160),
            .lcout(n2284),
            .ltout(),
            .carryin(n12692),
            .carryout(n12693),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_20_lut_LC_3_16_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_20_lut_LC_3_16_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_20_lut_LC_3_16_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_20_lut_LC_3_16_2 (
            .in0(_gnd_net_),
            .in1(N__30992),
            .in2(N__55035),
            .in3(N__23247),
            .lcout(n2283),
            .ltout(),
            .carryin(n12693),
            .carryout(n12694),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_21_lut_LC_3_16_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1503_21_lut_LC_3_16_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_21_lut_LC_3_16_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1503_21_lut_LC_3_16_3 (
            .in0(_gnd_net_),
            .in1(N__28488),
            .in2(N__55034),
            .in3(N__23244),
            .lcout(n2282),
            .ltout(),
            .carryin(n12694),
            .carryout(n12695),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1503_22_lut_LC_3_16_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1503_22_lut_LC_3_16_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1503_22_lut_LC_3_16_4.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1503_22_lut_LC_3_16_4 (
            .in0(N__25578),
            .in1(N__35612),
            .in2(N__55036),
            .in3(N__23241),
            .lcout(n2313),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10000_4_lut_LC_3_16_6.C_ON=1'b0;
    defparam i10000_4_lut_LC_3_16_6.SEQ_MODE=4'b0000;
    defparam i10000_4_lut_LC_3_16_6.LUT_INIT=16'b1111111010101010;
    LogicCell40 i10000_4_lut_LC_3_16_6 (
            .in0(N__25201),
            .in1(N__38210),
            .in2(N__23234),
            .in3(N__25231),
            .lcout(n11977),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1457_3_lut_LC_3_17_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1457_3_lut_LC_3_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1457_3_lut_LC_3_17_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i1457_3_lut_LC_3_17_0 (
            .in0(N__33633),
            .in1(N__25317),
            .in2(_gnd_net_),
            .in3(N__35447),
            .lcout(n2233),
            .ltout(n2233_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1524_3_lut_LC_3_17_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1524_3_lut_LC_3_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1524_3_lut_LC_3_17_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1524_3_lut_LC_3_17_1 (
            .in0(_gnd_net_),
            .in1(N__23217),
            .in2(N__23208),
            .in3(N__35574),
            .lcout(n2332),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1523_3_lut_LC_3_17_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1523_3_lut_LC_3_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1523_3_lut_LC_3_17_2.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i1523_3_lut_LC_3_17_2 (
            .in0(N__25236),
            .in1(N__23205),
            .in2(N__35595),
            .in3(_gnd_net_),
            .lcout(n2331),
            .ltout(n2331_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9994_4_lut_LC_3_17_3.C_ON=1'b0;
    defparam i9994_4_lut_LC_3_17_3.SEQ_MODE=4'b0000;
    defparam i9994_4_lut_LC_3_17_3.LUT_INIT=16'b1111111011110000;
    LogicCell40 i9994_4_lut_LC_3_17_3 (
            .in0(N__38345),
            .in1(N__29104),
            .in2(N__23196),
            .in3(N__28720),
            .lcout(n11971),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1525_3_lut_LC_3_17_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1525_3_lut_LC_3_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1525_3_lut_LC_3_17_4.LUT_INIT=16'b1100101011001010;
    LogicCell40 encoder0_position_31__I_0_i1525_3_lut_LC_3_17_4 (
            .in0(N__23193),
            .in1(N__38211),
            .in2(N__35594),
            .in3(_gnd_net_),
            .lcout(n2333),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_38_LC_3_17_5.C_ON=1'b0;
    defparam i1_4_lut_adj_38_LC_3_17_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_38_LC_3_17_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_38_LC_3_17_5 (
            .in0(N__28336),
            .in1(N__23303),
            .in2(N__25177),
            .in3(N__25323),
            .lcout(n14594),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13018_1_lut_LC_3_17_6.C_ON=1'b0;
    defparam i13018_1_lut_LC_3_17_6.SEQ_MODE=4'b0000;
    defparam i13018_1_lut_LC_3_17_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 i13018_1_lut_LC_3_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35596),
            .in3(_gnd_net_),
            .lcout(n15748),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1446_3_lut_LC_3_18_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1446_3_lut_LC_3_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1446_3_lut_LC_3_18_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1446_3_lut_LC_3_18_0 (
            .in0(_gnd_net_),
            .in1(N__25440),
            .in2(N__31200),
            .in3(N__35436),
            .lcout(n2222),
            .ltout(n2222_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1513_3_lut_LC_3_18_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1513_3_lut_LC_3_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1513_3_lut_LC_3_18_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1513_3_lut_LC_3_18_1 (
            .in0(N__35538),
            .in1(_gnd_net_),
            .in2(N__23292),
            .in3(N__23289),
            .lcout(n2321),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1515_3_lut_LC_3_18_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1515_3_lut_LC_3_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1515_3_lut_LC_3_18_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1515_3_lut_LC_3_18_2 (
            .in0(_gnd_net_),
            .in1(N__23280),
            .in2(N__28304),
            .in3(N__35537),
            .lcout(n2323),
            .ltout(n2323_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_42_LC_3_18_3.C_ON=1'b0;
    defparam i1_4_lut_adj_42_LC_3_18_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_42_LC_3_18_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_42_LC_3_18_3 (
            .in0(N__28849),
            .in1(N__25636),
            .in2(N__23271),
            .in3(N__28774),
            .lcout(n14382),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1443_3_lut_LC_3_18_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1443_3_lut_LC_3_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1443_3_lut_LC_3_18_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1443_3_lut_LC_3_18_4 (
            .in0(_gnd_net_),
            .in1(N__25416),
            .in2(N__33114),
            .in3(N__35437),
            .lcout(n2219),
            .ltout(n2219_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1510_3_lut_LC_3_18_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1510_3_lut_LC_3_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1510_3_lut_LC_3_18_5.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1510_3_lut_LC_3_18_5 (
            .in0(N__35539),
            .in1(_gnd_net_),
            .in2(N__23268),
            .in3(N__23265),
            .lcout(n2318),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1514_3_lut_LC_3_18_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1514_3_lut_LC_3_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1514_3_lut_LC_3_18_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1514_3_lut_LC_3_18_6 (
            .in0(_gnd_net_),
            .in1(N__23256),
            .in2(N__28340),
            .in3(N__35533),
            .lcout(n2322),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1517_3_lut_LC_3_18_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1517_3_lut_LC_3_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1517_3_lut_LC_3_18_7.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1517_3_lut_LC_3_18_7 (
            .in0(_gnd_net_),
            .in1(N__25377),
            .in2(N__35573),
            .in3(N__23406),
            .lcout(n2325),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1522_3_lut_LC_3_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1522_3_lut_LC_3_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1522_3_lut_LC_3_19_0.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1522_3_lut_LC_3_19_0 (
            .in0(N__23397),
            .in1(_gnd_net_),
            .in2(N__35588),
            .in3(N__25212),
            .lcout(n2330),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1519_rep_17_3_lut_LC_3_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1519_rep_17_3_lut_LC_3_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1519_rep_17_3_lut_LC_3_19_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1519_rep_17_3_lut_LC_3_19_1 (
            .in0(_gnd_net_),
            .in1(N__23388),
            .in2(N__25404),
            .in3(N__35554),
            .lcout(n2327),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1520_3_lut_LC_3_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1520_3_lut_LC_3_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1520_3_lut_LC_3_19_2.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1520_3_lut_LC_3_19_2 (
            .in0(N__25151),
            .in1(_gnd_net_),
            .in2(N__35587),
            .in3(N__23379),
            .lcout(n2328),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_39_LC_3_19_3.C_ON=1'b0;
    defparam i1_2_lut_adj_39_LC_3_19_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_39_LC_3_19_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 i1_2_lut_adj_39_LC_3_19_3 (
            .in0(_gnd_net_),
            .in1(N__25150),
            .in2(_gnd_net_),
            .in3(N__28384),
            .lcout(),
            .ltout(n14808_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_40_LC_3_19_4.C_ON=1'b0;
    defparam i1_4_lut_adj_40_LC_3_19_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_40_LC_3_19_4.LUT_INIT=16'b1111111111101010;
    LogicCell40 i1_4_lut_adj_40_LC_3_19_4 (
            .in0(N__25486),
            .in1(N__23370),
            .in2(N__23361),
            .in3(N__23358),
            .lcout(),
            .ltout(n14598_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_41_LC_3_19_5.C_ON=1'b0;
    defparam i1_4_lut_adj_41_LC_3_19_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_41_LC_3_19_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_41_LC_3_19_5 (
            .in0(N__25529),
            .in1(N__23342),
            .in2(N__23331),
            .in3(N__28531),
            .lcout(),
            .ltout(n14604_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13021_4_lut_LC_3_19_6.C_ON=1'b0;
    defparam i13021_4_lut_LC_3_19_6.SEQ_MODE=4'b0000;
    defparam i13021_4_lut_LC_3_19_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 i13021_4_lut_LC_3_19_6 (
            .in0(N__30985),
            .in1(N__28484),
            .in2(N__23328),
            .in3(N__25574),
            .lcout(n2247),
            .ltout(n2247_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1521_3_lut_LC_3_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1521_3_lut_LC_3_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1521_3_lut_LC_3_19_7.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1521_3_lut_LC_3_19_7 (
            .in0(_gnd_net_),
            .in1(N__28385),
            .in2(N__23325),
            .in3(N__23322),
            .lcout(n2329),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1512_3_lut_LC_3_20_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1512_3_lut_LC_3_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1512_3_lut_LC_3_20_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1512_3_lut_LC_3_20_0 (
            .in0(_gnd_net_),
            .in1(N__23523),
            .in2(N__25185),
            .in3(N__35561),
            .lcout(n2320),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12484_3_lut_LC_3_20_1.C_ON=1'b0;
    defparam i12484_3_lut_LC_3_20_1.SEQ_MODE=4'b0000;
    defparam i12484_3_lut_LC_3_20_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 i12484_3_lut_LC_3_20_1 (
            .in0(_gnd_net_),
            .in1(N__23514),
            .in2(N__23462),
            .in3(N__35716),
            .lcout(n2423),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1511_3_lut_LC_3_20_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1511_3_lut_LC_3_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1511_3_lut_LC_3_20_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1511_3_lut_LC_3_20_2 (
            .in0(N__23505),
            .in1(N__25490),
            .in2(_gnd_net_),
            .in3(N__35562),
            .lcout(n2319),
            .ltout(n2319_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1578_3_lut_LC_3_20_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1578_3_lut_LC_3_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1578_3_lut_LC_3_20_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1578_3_lut_LC_3_20_3 (
            .in0(_gnd_net_),
            .in1(N__23496),
            .in2(N__23487),
            .in3(N__35717),
            .lcout(n2418),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_46_LC_3_20_4.C_ON=1'b0;
    defparam i1_4_lut_adj_46_LC_3_20_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_46_LC_3_20_4.LUT_INIT=16'b1111111110000000;
    LogicCell40 i1_4_lut_adj_46_LC_3_20_4 (
            .in0(N__25894),
            .in1(N__23484),
            .in2(N__28831),
            .in3(N__23412),
            .lcout(n14392),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12483_3_lut_LC_3_20_5.C_ON=1'b0;
    defparam i12483_3_lut_LC_3_20_5.SEQ_MODE=4'b0000;
    defparam i12483_3_lut_LC_3_20_5.LUT_INIT=16'b1100101011001010;
    LogicCell40 i12483_3_lut_LC_3_20_5 (
            .in0(N__23475),
            .in1(N__25353),
            .in2(N__35589),
            .in3(_gnd_net_),
            .lcout(n2324),
            .ltout(n2324_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_43_LC_3_20_6.C_ON=1'b0;
    defparam i1_4_lut_adj_43_LC_3_20_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_43_LC_3_20_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_43_LC_3_20_6 (
            .in0(N__25864),
            .in1(N__25774),
            .in2(N__23442),
            .in3(N__28681),
            .lcout(),
            .ltout(n14384_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_45_LC_3_20_7.C_ON=1'b0;
    defparam i1_4_lut_adj_45_LC_3_20_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_45_LC_3_20_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_45_LC_3_20_7 (
            .in0(N__25618),
            .in1(N__23435),
            .in2(N__23424),
            .in3(N__23421),
            .lcout(n14390),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1718_3_lut_LC_3_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1718_3_lut_LC_3_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1718_3_lut_LC_3_21_0.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1718_3_lut_LC_3_21_0 (
            .in0(N__32499),
            .in1(_gnd_net_),
            .in2(N__36102),
            .in3(N__32513),
            .lcout(n2622),
            .ltout(n2622_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1785_3_lut_LC_3_21_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1785_3_lut_LC_3_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1785_3_lut_LC_3_21_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1785_3_lut_LC_3_21_1 (
            .in0(_gnd_net_),
            .in1(N__23772),
            .in2(N__23760),
            .in3(N__36268),
            .lcout(n2721),
            .ltout(n2721_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_55_LC_3_21_2.C_ON=1'b0;
    defparam i1_4_lut_adj_55_LC_3_21_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_55_LC_3_21_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_55_LC_3_21_2 (
            .in0(N__23726),
            .in1(N__23708),
            .in2(N__23697),
            .in3(N__23620),
            .lcout(n14348),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1719_3_lut_LC_3_21_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1719_3_lut_LC_3_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1719_3_lut_LC_3_21_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1719_3_lut_LC_3_21_3 (
            .in0(_gnd_net_),
            .in1(N__32070),
            .in2(N__32090),
            .in3(N__36094),
            .lcout(n2623),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1575_3_lut_LC_3_21_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1575_3_lut_LC_3_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1575_3_lut_LC_3_21_4.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1575_3_lut_LC_3_21_4 (
            .in0(N__23685),
            .in1(_gnd_net_),
            .in2(N__35745),
            .in3(N__25727),
            .lcout(n2415),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1724_3_lut_LC_3_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1724_3_lut_LC_3_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1724_3_lut_LC_3_21_5.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1724_3_lut_LC_3_21_5 (
            .in0(N__32244),
            .in1(_gnd_net_),
            .in2(N__32217),
            .in3(N__36090),
            .lcout(n2628),
            .ltout(n2628_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_32_LC_3_21_6.C_ON=1'b0;
    defparam i1_4_lut_adj_32_LC_3_21_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_32_LC_3_21_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_32_LC_3_21_6 (
            .in0(N__26017),
            .in1(N__23666),
            .in2(N__23655),
            .in3(N__33907),
            .lcout(n14668),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1788_3_lut_LC_3_21_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1788_3_lut_LC_3_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1788_3_lut_LC_3_21_7.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i1788_3_lut_LC_3_21_7 (
            .in0(_gnd_net_),
            .in1(N__36267),
            .in2(N__25964),
            .in3(N__23652),
            .lcout(n2724),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1791_3_lut_LC_3_22_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1791_3_lut_LC_3_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1791_3_lut_LC_3_22_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1791_3_lut_LC_3_22_0 (
            .in0(_gnd_net_),
            .in1(N__23604),
            .in2(N__23582),
            .in3(N__36224),
            .lcout(n2727),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1796_3_lut_LC_3_22_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1796_3_lut_LC_3_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1796_3_lut_LC_3_22_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1796_3_lut_LC_3_22_1 (
            .in0(_gnd_net_),
            .in1(N__23538),
            .in2(N__36276),
            .in3(N__26261),
            .lcout(n2732),
            .ltout(n2732_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9980_3_lut_LC_3_22_2.C_ON=1'b0;
    defparam i9980_3_lut_LC_3_22_2.SEQ_MODE=4'b0000;
    defparam i9980_3_lut_LC_3_22_2.LUT_INIT=16'b1111000011000000;
    LogicCell40 i9980_3_lut_LC_3_22_2 (
            .in0(_gnd_net_),
            .in1(N__26614),
            .in2(N__23919),
            .in3(N__33523),
            .lcout(),
            .ltout(n11957_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_58_LC_3_22_3.C_ON=1'b0;
    defparam i1_4_lut_adj_58_LC_3_22_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_58_LC_3_22_3.LUT_INIT=16'b1000100010000000;
    LogicCell40 i1_4_lut_adj_58_LC_3_22_3 (
            .in0(N__23905),
            .in1(N__23827),
            .in2(N__23889),
            .in3(N__24352),
            .lcout(n13808),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_50_LC_3_22_4.C_ON=1'b0;
    defparam i1_4_lut_adj_50_LC_3_22_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_50_LC_3_22_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_50_LC_3_22_4 (
            .in0(N__29383),
            .in1(N__23870),
            .in2(N__26231),
            .in3(N__23859),
            .lcout(n14674),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1794_3_lut_LC_3_22_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1794_3_lut_LC_3_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1794_3_lut_LC_3_22_5.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1794_3_lut_LC_3_22_5 (
            .in0(_gnd_net_),
            .in1(N__29195),
            .in2(N__36277),
            .in3(N__23853),
            .lcout(n2730),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1795_3_lut_LC_3_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1795_3_lut_LC_3_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1795_3_lut_LC_3_22_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1795_3_lut_LC_3_22_7 (
            .in0(N__23811),
            .in1(_gnd_net_),
            .in2(N__36278),
            .in3(N__29252),
            .lcout(n2731),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1797_3_lut_LC_3_23_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1797_3_lut_LC_3_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1797_3_lut_LC_3_23_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i1797_3_lut_LC_3_23_1 (
            .in0(N__33577),
            .in1(N__23796),
            .in2(_gnd_net_),
            .in3(N__36240),
            .lcout(n2733),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_28_LC_3_23_2.C_ON=1'b0;
    defparam i1_4_lut_adj_28_LC_3_23_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_28_LC_3_23_2.LUT_INIT=16'b1111111011101110;
    LogicCell40 i1_4_lut_adj_28_LC_3_23_2 (
            .in0(N__26134),
            .in1(N__24124),
            .in2(N__26244),
            .in3(N__25827),
            .lcout(),
            .ltout(n14650_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_31_LC_3_23_3.C_ON=1'b0;
    defparam i1_4_lut_adj_31_LC_3_23_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_31_LC_3_23_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_31_LC_3_23_3 (
            .in0(N__29683),
            .in1(N__32617),
            .in2(N__23778),
            .in3(N__25932),
            .lcout(),
            .ltout(n14654_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_34_LC_3_23_4.C_ON=1'b0;
    defparam i1_4_lut_adj_34_LC_3_23_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_34_LC_3_23_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_34_LC_3_23_4 (
            .in0(N__26164),
            .in1(N__26191),
            .in2(N__23775),
            .in3(N__29533),
            .lcout(),
            .ltout(n14660_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12565_4_lut_LC_3_23_5.C_ON=1'b0;
    defparam i12565_4_lut_LC_3_23_5.SEQ_MODE=4'b0000;
    defparam i12565_4_lut_LC_3_23_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12565_4_lut_LC_3_23_5 (
            .in0(N__32548),
            .in1(N__32722),
            .in2(N__24189),
            .in3(N__24186),
            .lcout(n2643),
            .ltout(n2643_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1782_3_lut_LC_3_23_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1782_3_lut_LC_3_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1782_3_lut_LC_3_23_6.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1782_3_lut_LC_3_23_6 (
            .in0(N__26135),
            .in1(_gnd_net_),
            .in2(N__24180),
            .in3(N__24177),
            .lcout(n2718),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1786_3_lut_LC_3_23_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1786_3_lut_LC_3_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1786_3_lut_LC_3_23_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1786_3_lut_LC_3_23_7 (
            .in0(_gnd_net_),
            .in1(N__24144),
            .in2(N__24129),
            .in3(N__36241),
            .lcout(n2722),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1863_3_lut_LC_3_24_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1863_3_lut_LC_3_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1863_3_lut_LC_3_24_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1863_3_lut_LC_3_24_0 (
            .in0(_gnd_net_),
            .in1(N__24074),
            .in2(N__24054),
            .in3(N__36427),
            .lcout(n2831),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1842_3_lut_LC_3_24_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1842_3_lut_LC_3_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1842_3_lut_LC_3_24_1.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1842_3_lut_LC_3_24_1 (
            .in0(N__24035),
            .in1(_gnd_net_),
            .in2(N__36455),
            .in3(N__24021),
            .lcout(n2810),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1850_3_lut_LC_3_24_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1850_3_lut_LC_3_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1850_3_lut_LC_3_24_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1850_3_lut_LC_3_24_2 (
            .in0(_gnd_net_),
            .in1(N__24003),
            .in2(N__23991),
            .in3(N__36429),
            .lcout(n2818),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1781_3_lut_LC_3_24_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1781_3_lut_LC_3_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1781_3_lut_LC_3_24_3.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1781_3_lut_LC_3_24_3 (
            .in0(N__26230),
            .in1(_gnd_net_),
            .in2(N__36281),
            .in3(N__23967),
            .lcout(n2717),
            .ltout(n2717_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1848_3_lut_LC_3_24_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1848_3_lut_LC_3_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1848_3_lut_LC_3_24_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1848_3_lut_LC_3_24_4 (
            .in0(_gnd_net_),
            .in1(N__23934),
            .in2(N__23922),
            .in3(N__36430),
            .lcout(n2816),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1844_3_lut_LC_3_24_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1844_3_lut_LC_3_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1844_3_lut_LC_3_24_5.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1844_3_lut_LC_3_24_5 (
            .in0(_gnd_net_),
            .in1(N__24416),
            .in2(N__36454),
            .in3(N__24393),
            .lcout(n2812),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1862_3_lut_LC_3_24_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1862_3_lut_LC_3_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1862_3_lut_LC_3_24_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1862_3_lut_LC_3_24_6 (
            .in0(_gnd_net_),
            .in1(N__24381),
            .in2(N__24368),
            .in3(N__36428),
            .lcout(n2830),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1776_3_lut_LC_3_24_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1776_3_lut_LC_3_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1776_3_lut_LC_3_24_7.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1776_3_lut_LC_3_24_7 (
            .in0(_gnd_net_),
            .in1(N__26168),
            .in2(N__36282),
            .in3(N__24336),
            .lcout(n2712),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1919_3_lut_LC_3_25_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1919_3_lut_LC_3_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1919_3_lut_LC_3_25_0.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i1919_3_lut_LC_3_25_0 (
            .in0(N__24308),
            .in1(N__24321),
            .in2(N__34323),
            .in3(_gnd_net_),
            .lcout(n2919),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_62_LC_3_25_1.C_ON=1'b0;
    defparam i1_4_lut_adj_62_LC_3_25_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_62_LC_3_25_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_62_LC_3_25_1 (
            .in0(N__24616),
            .in1(N__29329),
            .in2(N__26750),
            .in3(N__29827),
            .lcout(),
            .ltout(n14690_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_63_LC_3_25_2.C_ON=1'b0;
    defparam i1_4_lut_adj_63_LC_3_25_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_63_LC_3_25_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_63_LC_3_25_2 (
            .in0(N__24307),
            .in1(N__26833),
            .in2(N__24294),
            .in3(N__24291),
            .lcout(),
            .ltout(n14696_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_65_LC_3_25_3.C_ON=1'b0;
    defparam i1_4_lut_adj_65_LC_3_25_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_65_LC_3_25_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_65_LC_3_25_3 (
            .in0(N__27239),
            .in1(N__26281),
            .in2(N__24282),
            .in3(N__26514),
            .lcout(n14702),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1845_3_lut_LC_3_25_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1845_3_lut_LC_3_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1845_3_lut_LC_3_25_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1845_3_lut_LC_3_25_4 (
            .in0(_gnd_net_),
            .in1(N__24277),
            .in2(N__24246),
            .in3(N__36410),
            .lcout(n2813),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1851_3_lut_LC_3_25_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1851_3_lut_LC_3_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1851_3_lut_LC_3_25_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1851_3_lut_LC_3_25_6 (
            .in0(_gnd_net_),
            .in1(N__24231),
            .in2(N__24204),
            .in3(N__36409),
            .lcout(n2819),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1922_3_lut_LC_3_25_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1922_3_lut_LC_3_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1922_3_lut_LC_3_25_7.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1922_3_lut_LC_3_25_7 (
            .in0(N__24617),
            .in1(_gnd_net_),
            .in2(N__24603),
            .in3(N__34293),
            .lcout(n2922),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1926_3_lut_LC_3_26_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1926_3_lut_LC_3_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1926_3_lut_LC_3_26_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1926_3_lut_LC_3_26_0 (
            .in0(_gnd_net_),
            .in1(N__24588),
            .in2(N__24561),
            .in3(N__34277),
            .lcout(n2926),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1921_3_lut_LC_3_26_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1921_3_lut_LC_3_26_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1921_3_lut_LC_3_26_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1921_3_lut_LC_3_26_2 (
            .in0(_gnd_net_),
            .in1(N__24546),
            .in2(N__24519),
            .in3(N__34278),
            .lcout(n2921),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1982_3_lut_LC_3_26_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1982_3_lut_LC_3_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1982_3_lut_LC_3_26_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1982_3_lut_LC_3_26_3 (
            .in0(_gnd_net_),
            .in1(N__27118),
            .in2(N__24504),
            .in3(N__34461),
            .lcout(n3014),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1986_3_lut_LC_3_26_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1986_3_lut_LC_3_26_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1986_3_lut_LC_3_26_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1986_3_lut_LC_3_26_5 (
            .in0(_gnd_net_),
            .in1(N__26655),
            .in2(N__24495),
            .in3(N__34460),
            .lcout(n3018),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i16_1_lut_LC_3_26_6.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i16_1_lut_LC_3_26_6.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i16_1_lut_LC_3_26_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i16_1_lut_LC_3_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46500),
            .lcout(n10_adj_582),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1911_3_lut_LC_3_26_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1911_3_lut_LC_3_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1911_3_lut_LC_3_26_7.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1911_3_lut_LC_3_26_7 (
            .in0(_gnd_net_),
            .in1(N__26472),
            .in2(N__34320),
            .in3(N__24486),
            .lcout(n2911),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1841_3_lut_LC_3_27_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1841_3_lut_LC_3_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1841_3_lut_LC_3_27_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1841_3_lut_LC_3_27_0 (
            .in0(_gnd_net_),
            .in1(N__24471),
            .in2(N__24444),
            .in3(N__36458),
            .lcout(n2809),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1996_3_lut_LC_3_27_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1996_3_lut_LC_3_27_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1996_3_lut_LC_3_27_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1996_3_lut_LC_3_27_1 (
            .in0(_gnd_net_),
            .in1(N__24426),
            .in2(N__27168),
            .in3(N__34453),
            .lcout(n3028),
            .ltout(n3028_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2063_3_lut_LC_3_27_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2063_3_lut_LC_3_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2063_3_lut_LC_3_27_2.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i2063_3_lut_LC_3_27_2 (
            .in0(N__24813),
            .in1(_gnd_net_),
            .in2(N__24672),
            .in3(N__34603),
            .lcout(n3127),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1988_3_lut_LC_3_27_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1988_3_lut_LC_3_27_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1988_3_lut_LC_3_27_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1988_3_lut_LC_3_27_3 (
            .in0(_gnd_net_),
            .in1(N__26700),
            .in2(N__24669),
            .in3(N__34454),
            .lcout(n3020),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1912_3_lut_LC_3_27_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1912_3_lut_LC_3_27_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1912_3_lut_LC_3_27_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1912_3_lut_LC_3_27_4 (
            .in0(_gnd_net_),
            .in1(N__24660),
            .in2(N__26448),
            .in3(N__34332),
            .lcout(n2912),
            .ltout(n2912_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1979_3_lut_LC_3_27_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1979_3_lut_LC_3_27_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1979_3_lut_LC_3_27_5.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1979_3_lut_LC_3_27_5 (
            .in0(N__24648),
            .in1(_gnd_net_),
            .in2(N__24642),
            .in3(N__34459),
            .lcout(n3011),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12654_1_lut_LC_3_27_6.C_ON=1'b0;
    defparam i12654_1_lut_LC_3_27_6.SEQ_MODE=4'b0000;
    defparam i12654_1_lut_LC_3_27_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12654_1_lut_LC_3_27_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34502),
            .in3(_gnd_net_),
            .lcout(n15384),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1983_3_lut_LC_3_27_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1983_3_lut_LC_3_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1983_3_lut_LC_3_27_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1983_3_lut_LC_3_27_7 (
            .in0(_gnd_net_),
            .in1(N__27200),
            .in2(N__24639),
            .in3(N__34458),
            .lcout(n3015),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_2_lut_LC_3_28_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_2_lut_LC_3_28_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_2_lut_LC_3_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_2_lut_LC_3_28_0 (
            .in0(_gnd_net_),
            .in1(N__41570),
            .in2(_gnd_net_),
            .in3(N__24630),
            .lcout(n3101),
            .ltout(),
            .carryin(bfn_3_28_0_),
            .carryout(n12864),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_3_lut_LC_3_28_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_3_lut_LC_3_28_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_3_lut_LC_3_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_3_lut_LC_3_28_1 (
            .in0(_gnd_net_),
            .in1(N__54443),
            .in2(N__30099),
            .in3(N__24627),
            .lcout(n3100),
            .ltout(),
            .carryin(n12864),
            .carryout(n12865),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_4_lut_LC_3_28_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_4_lut_LC_3_28_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_4_lut_LC_3_28_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_4_lut_LC_3_28_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30078),
            .in3(N__24624),
            .lcout(n3099),
            .ltout(),
            .carryin(n12865),
            .carryout(n12866),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_5_lut_LC_3_28_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_5_lut_LC_3_28_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_5_lut_LC_3_28_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_5_lut_LC_3_28_3 (
            .in0(_gnd_net_),
            .in1(N__54444),
            .in2(N__29931),
            .in3(N__24849),
            .lcout(n3098),
            .ltout(),
            .carryin(n12866),
            .carryout(n12867),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_6_lut_LC_3_28_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_6_lut_LC_3_28_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_6_lut_LC_3_28_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_6_lut_LC_3_28_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29979),
            .in3(N__24846),
            .lcout(n3097),
            .ltout(),
            .carryin(n12867),
            .carryout(n12868),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_7_lut_LC_3_28_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_7_lut_LC_3_28_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_7_lut_LC_3_28_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_7_lut_LC_3_28_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29954),
            .in3(N__24834),
            .lcout(n3096),
            .ltout(),
            .carryin(n12868),
            .carryout(n12869),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_8_lut_LC_3_28_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_8_lut_LC_3_28_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_8_lut_LC_3_28_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_8_lut_LC_3_28_6 (
            .in0(_gnd_net_),
            .in1(N__54446),
            .in2(N__24831),
            .in3(N__24807),
            .lcout(n3095),
            .ltout(),
            .carryin(n12869),
            .carryout(n12870),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_9_lut_LC_3_28_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_9_lut_LC_3_28_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_9_lut_LC_3_28_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_9_lut_LC_3_28_7 (
            .in0(_gnd_net_),
            .in1(N__54445),
            .in2(N__30587),
            .in3(N__24795),
            .lcout(n3094),
            .ltout(),
            .carryin(n12870),
            .carryout(n12871),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_10_lut_LC_3_29_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_10_lut_LC_3_29_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_10_lut_LC_3_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_10_lut_LC_3_29_0 (
            .in0(_gnd_net_),
            .in1(N__54574),
            .in2(N__24792),
            .in3(N__24753),
            .lcout(n3093),
            .ltout(),
            .carryin(bfn_3_29_0_),
            .carryout(n12872),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_11_lut_LC_3_29_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_11_lut_LC_3_29_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_11_lut_LC_3_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_11_lut_LC_3_29_1 (
            .in0(_gnd_net_),
            .in1(N__54578),
            .in2(N__24750),
            .in3(N__24714),
            .lcout(n3092),
            .ltout(),
            .carryin(n12872),
            .carryout(n12873),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_12_lut_LC_3_29_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_12_lut_LC_3_29_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_12_lut_LC_3_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_12_lut_LC_3_29_2 (
            .in0(_gnd_net_),
            .in1(N__54575),
            .in2(N__24711),
            .in3(N__24675),
            .lcout(n3091),
            .ltout(),
            .carryin(n12873),
            .carryout(n12874),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_13_lut_LC_3_29_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_13_lut_LC_3_29_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_13_lut_LC_3_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_13_lut_LC_3_29_3 (
            .in0(_gnd_net_),
            .in1(N__54579),
            .in2(N__30561),
            .in3(N__25020),
            .lcout(n3090),
            .ltout(),
            .carryin(n12874),
            .carryout(n12875),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_14_lut_LC_3_29_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_14_lut_LC_3_29_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_14_lut_LC_3_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_14_lut_LC_3_29_4 (
            .in0(_gnd_net_),
            .in1(N__54576),
            .in2(N__25017),
            .in3(N__24981),
            .lcout(n3089),
            .ltout(),
            .carryin(n12875),
            .carryout(n12876),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_15_lut_LC_3_29_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_15_lut_LC_3_29_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_15_lut_LC_3_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_15_lut_LC_3_29_5 (
            .in0(_gnd_net_),
            .in1(N__54580),
            .in2(N__24977),
            .in3(N__24942),
            .lcout(n3088),
            .ltout(),
            .carryin(n12876),
            .carryout(n12877),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_16_lut_LC_3_29_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_16_lut_LC_3_29_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_16_lut_LC_3_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_16_lut_LC_3_29_6 (
            .in0(_gnd_net_),
            .in1(N__54577),
            .in2(N__24939),
            .in3(N__24906),
            .lcout(n3087),
            .ltout(),
            .carryin(n12877),
            .carryout(n12878),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_17_lut_LC_3_29_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_17_lut_LC_3_29_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_17_lut_LC_3_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_17_lut_LC_3_29_7 (
            .in0(_gnd_net_),
            .in1(N__54581),
            .in2(N__30624),
            .in3(N__24894),
            .lcout(n3086),
            .ltout(),
            .carryin(n12878),
            .carryout(n12879),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_18_lut_LC_3_30_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_18_lut_LC_3_30_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_18_lut_LC_3_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_18_lut_LC_3_30_0 (
            .in0(_gnd_net_),
            .in1(N__27282),
            .in2(N__54864),
            .in3(N__24891),
            .lcout(n3085),
            .ltout(),
            .carryin(bfn_3_30_0_),
            .carryout(n12880),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_19_lut_LC_3_30_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_19_lut_LC_3_30_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_19_lut_LC_3_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_19_lut_LC_3_30_1 (
            .in0(_gnd_net_),
            .in1(N__24888),
            .in2(N__54868),
            .in3(N__24855),
            .lcout(n3084),
            .ltout(),
            .carryin(n12880),
            .carryout(n12881),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_20_lut_LC_3_30_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_20_lut_LC_3_30_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_20_lut_LC_3_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_20_lut_LC_3_30_2 (
            .in0(_gnd_net_),
            .in1(N__30323),
            .in2(N__54865),
            .in3(N__24852),
            .lcout(n3083),
            .ltout(),
            .carryin(n12881),
            .carryout(n12882),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_21_lut_LC_3_30_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_21_lut_LC_3_30_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_21_lut_LC_3_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_21_lut_LC_3_30_3 (
            .in0(_gnd_net_),
            .in1(N__27494),
            .in2(N__54869),
            .in3(N__25062),
            .lcout(n3082),
            .ltout(),
            .carryin(n12882),
            .carryout(n12883),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_22_lut_LC_3_30_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_22_lut_LC_3_30_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_22_lut_LC_3_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_22_lut_LC_3_30_4 (
            .in0(_gnd_net_),
            .in1(N__27462),
            .in2(N__54866),
            .in3(N__25059),
            .lcout(n3081),
            .ltout(),
            .carryin(n12883),
            .carryout(n12884),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_23_lut_LC_3_30_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_23_lut_LC_3_30_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_23_lut_LC_3_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_23_lut_LC_3_30_5 (
            .in0(_gnd_net_),
            .in1(N__27587),
            .in2(N__54870),
            .in3(N__25056),
            .lcout(n3080),
            .ltout(),
            .carryin(n12884),
            .carryout(n12885),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_24_lut_LC_3_30_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_24_lut_LC_3_30_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_24_lut_LC_3_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_24_lut_LC_3_30_6 (
            .in0(_gnd_net_),
            .in1(N__30251),
            .in2(N__54867),
            .in3(N__25053),
            .lcout(n3079),
            .ltout(),
            .carryin(n12885),
            .carryout(n12886),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_25_lut_LC_3_30_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_25_lut_LC_3_30_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_25_lut_LC_3_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_25_lut_LC_3_30_7 (
            .in0(_gnd_net_),
            .in1(N__54534),
            .in2(N__27431),
            .in3(N__25050),
            .lcout(n3078),
            .ltout(),
            .carryin(n12886),
            .carryout(n12887),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_26_lut_LC_3_31_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_26_lut_LC_3_31_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_26_lut_LC_3_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_26_lut_LC_3_31_0 (
            .in0(_gnd_net_),
            .in1(N__28208),
            .in2(N__54860),
            .in3(N__25047),
            .lcout(n3077),
            .ltout(),
            .carryin(bfn_3_31_0_),
            .carryout(n12888),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_27_lut_LC_3_31_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_27_lut_LC_3_31_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_27_lut_LC_3_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_27_lut_LC_3_31_1 (
            .in0(_gnd_net_),
            .in1(N__27404),
            .in2(N__54862),
            .in3(N__25044),
            .lcout(n3076),
            .ltout(),
            .carryin(n12888),
            .carryout(n12889),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_28_lut_LC_3_31_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_28_lut_LC_3_31_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_28_lut_LC_3_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_28_lut_LC_3_31_2 (
            .in0(_gnd_net_),
            .in1(N__27347),
            .in2(N__54861),
            .in3(N__25041),
            .lcout(n3075),
            .ltout(),
            .carryin(n12889),
            .carryout(n12890),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_29_lut_LC_3_31_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2039_29_lut_LC_3_31_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_29_lut_LC_3_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2039_29_lut_LC_3_31_3 (
            .in0(_gnd_net_),
            .in1(N__27323),
            .in2(N__54863),
            .in3(N__25038),
            .lcout(n3074),
            .ltout(),
            .carryin(n12890),
            .carryout(n12891),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2039_30_lut_LC_3_31_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_2039_30_lut_LC_3_31_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2039_30_lut_LC_3_31_4.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_2039_30_lut_LC_3_31_4 (
            .in0(N__54515),
            .in1(N__34739),
            .in2(N__27369),
            .in3(N__25128),
            .lcout(n3105),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2043_3_lut_LC_3_31_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2043_3_lut_LC_3_31_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2043_3_lut_LC_3_31_5.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i2043_3_lut_LC_3_31_5 (
            .in0(N__27348),
            .in1(_gnd_net_),
            .in2(N__25125),
            .in3(N__34664),
            .lcout(n3107),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2050_3_lut_LC_3_31_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2050_3_lut_LC_3_31_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2050_3_lut_LC_3_31_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2050_3_lut_LC_3_31_6 (
            .in0(_gnd_net_),
            .in1(N__25116),
            .in2(N__34697),
            .in3(N__27498),
            .lcout(n3114),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2042_3_lut_LC_3_31_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2042_3_lut_LC_3_31_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2042_3_lut_LC_3_31_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2042_3_lut_LC_3_31_7 (
            .in0(_gnd_net_),
            .in1(N__27324),
            .in2(N__25110),
            .in3(N__34665),
            .lcout(n3106),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2109_3_lut_LC_3_32_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2109_3_lut_LC_3_32_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2109_3_lut_LC_3_32_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i2109_3_lut_LC_3_32_0 (
            .in0(_gnd_net_),
            .in1(N__28059),
            .in2(N__34906),
            .in3(N__25101),
            .lcout(n3205),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12721_1_lut_LC_3_32_1.C_ON=1'b0;
    defparam i12721_1_lut_LC_3_32_1.SEQ_MODE=4'b0000;
    defparam i12721_1_lut_LC_3_32_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12721_1_lut_LC_3_32_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34858),
            .lcout(n15451),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2110_3_lut_LC_3_32_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2110_3_lut_LC_3_32_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2110_3_lut_LC_3_32_2.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2110_3_lut_LC_3_32_2 (
            .in0(_gnd_net_),
            .in1(N__25095),
            .in2(N__34907),
            .in3(N__28077),
            .lcout(n3206),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2047_3_lut_LC_3_32_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2047_3_lut_LC_3_32_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2047_3_lut_LC_3_32_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2047_3_lut_LC_3_32_3 (
            .in0(_gnd_net_),
            .in1(N__25089),
            .in2(N__30258),
            .in3(N__34698),
            .lcout(n3111),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2046_3_lut_LC_3_32_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2046_3_lut_LC_3_32_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2046_3_lut_LC_3_32_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2046_3_lut_LC_3_32_5 (
            .in0(_gnd_net_),
            .in1(N__27432),
            .in2(N__25080),
            .in3(N__34699),
            .lcout(n3110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2044_3_lut_LC_3_32_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2044_3_lut_LC_3_32_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2044_3_lut_LC_3_32_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2044_3_lut_LC_3_32_6 (
            .in0(_gnd_net_),
            .in1(N__25068),
            .in2(N__34714),
            .in3(N__27405),
            .lcout(n3108),
            .ltout(n3108_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2111_3_lut_LC_3_32_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2111_3_lut_LC_3_32_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2111_3_lut_LC_3_32_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2111_3_lut_LC_3_32_7 (
            .in0(_gnd_net_),
            .in1(N__25245),
            .in2(N__25239),
            .in3(N__34862),
            .lcout(n3207),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1456_3_lut_LC_4_15_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1456_3_lut_LC_4_15_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1456_3_lut_LC_4_15_0.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1456_3_lut_LC_4_15_0 (
            .in0(_gnd_net_),
            .in1(N__25308),
            .in2(N__35446),
            .in3(N__33677),
            .lcout(n2232),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1455_3_lut_LC_4_15_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1455_3_lut_LC_4_15_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1455_3_lut_LC_4_15_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1455_3_lut_LC_4_15_6 (
            .in0(_gnd_net_),
            .in1(N__25296),
            .in2(N__35445),
            .in3(N__33705),
            .lcout(n2231),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_33_LC_4_16_0.C_ON=1'b0;
    defparam i1_4_lut_adj_33_LC_4_16_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_33_LC_4_16_0.LUT_INIT=16'b1100000010000000;
    LogicCell40 i1_4_lut_adj_33_LC_4_16_0 (
            .in0(N__28097),
            .in1(N__28150),
            .in2(N__25271),
            .in3(N__33645),
            .lcout(n13787),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1450_3_lut_LC_4_16_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1450_3_lut_LC_4_16_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1450_3_lut_LC_4_16_1.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1450_3_lut_LC_4_16_1 (
            .in0(N__25467),
            .in1(_gnd_net_),
            .in2(N__28128),
            .in3(N__35419),
            .lcout(n2226),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1445_3_lut_LC_4_16_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1445_3_lut_LC_4_16_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1445_3_lut_LC_4_16_2.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1445_3_lut_LC_4_16_2 (
            .in0(_gnd_net_),
            .in1(N__28455),
            .in2(N__35444),
            .in3(N__25431),
            .lcout(n2221),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1449_rep_20_3_lut_LC_4_16_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1449_rep_20_3_lut_LC_4_16_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1449_rep_20_3_lut_LC_4_16_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1449_rep_20_3_lut_LC_4_16_3 (
            .in0(_gnd_net_),
            .in1(N__25458),
            .in2(N__28611),
            .in3(N__35418),
            .lcout(n2225),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1453_3_lut_LC_4_16_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1453_3_lut_LC_4_16_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1453_3_lut_LC_4_16_4.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1453_3_lut_LC_4_16_4 (
            .in0(_gnd_net_),
            .in1(N__25281),
            .in2(N__35443),
            .in3(N__28151),
            .lcout(n2229),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1385_3_lut_LC_4_16_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1385_3_lut_LC_4_16_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1385_3_lut_LC_4_16_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1385_3_lut_LC_4_16_5 (
            .in0(_gnd_net_),
            .in1(N__33777),
            .in2(N__31170),
            .in3(N__35298),
            .lcout(n2129),
            .ltout(n2129_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1452_3_lut_LC_4_16_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1452_3_lut_LC_4_16_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1452_3_lut_LC_4_16_6.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1452_3_lut_LC_4_16_6 (
            .in0(N__35420),
            .in1(_gnd_net_),
            .in2(N__25407),
            .in3(N__25254),
            .lcout(n2228),
            .ltout(n2228_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_37_LC_4_16_7.C_ON=1'b0;
    defparam i1_4_lut_adj_37_LC_4_16_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_37_LC_4_16_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_37_LC_4_16_7 (
            .in0(N__25369),
            .in1(N__25342),
            .in2(N__25326),
            .in3(N__28356),
            .lcout(n14588),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_2_lut_LC_4_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_2_lut_LC_4_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_2_lut_LC_4_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_2_lut_LC_4_17_0 (
            .in0(_gnd_net_),
            .in1(N__33632),
            .in2(_gnd_net_),
            .in3(N__25311),
            .lcout(n2201),
            .ltout(),
            .carryin(bfn_4_17_0_),
            .carryout(n12657),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_3_lut_LC_4_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_3_lut_LC_4_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_3_lut_LC_4_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_3_lut_LC_4_17_1 (
            .in0(_gnd_net_),
            .in1(N__55453),
            .in2(N__33678),
            .in3(N__25299),
            .lcout(n2200),
            .ltout(),
            .carryin(n12657),
            .carryout(n12658),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_4_lut_LC_4_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_4_lut_LC_4_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_4_lut_LC_4_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_4_lut_LC_4_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33704),
            .in3(N__25287),
            .lcout(n2199),
            .ltout(),
            .carryin(n12658),
            .carryout(n12659),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_5_lut_LC_4_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_5_lut_LC_4_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_5_lut_LC_4_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_5_lut_LC_4_17_3 (
            .in0(_gnd_net_),
            .in1(N__55454),
            .in2(N__28101),
            .in3(N__25284),
            .lcout(n2198),
            .ltout(),
            .carryin(n12659),
            .carryout(n12660),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_6_lut_LC_4_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_6_lut_LC_4_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_6_lut_LC_4_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_6_lut_LC_4_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28155),
            .in3(N__25275),
            .lcout(n2197),
            .ltout(),
            .carryin(n12660),
            .carryout(n12661),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_7_lut_LC_4_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_7_lut_LC_4_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_7_lut_LC_4_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_7_lut_LC_4_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25272),
            .in3(N__25248),
            .lcout(n2196),
            .ltout(),
            .carryin(n12661),
            .carryout(n12662),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_8_lut_LC_4_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_8_lut_LC_4_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_8_lut_LC_4_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_8_lut_LC_4_17_6 (
            .in0(_gnd_net_),
            .in1(N__54351),
            .in2(N__28224),
            .in3(N__25470),
            .lcout(n2195),
            .ltout(),
            .carryin(n12662),
            .carryout(n12663),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_9_lut_LC_4_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_9_lut_LC_4_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_9_lut_LC_4_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_9_lut_LC_4_17_7 (
            .in0(_gnd_net_),
            .in1(N__55455),
            .in2(N__28127),
            .in3(N__25461),
            .lcout(n2194),
            .ltout(),
            .carryin(n12663),
            .carryout(n12664),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_10_lut_LC_4_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_10_lut_LC_4_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_10_lut_LC_4_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_10_lut_LC_4_18_0 (
            .in0(_gnd_net_),
            .in1(N__55444),
            .in2(N__28607),
            .in3(N__25449),
            .lcout(n2193),
            .ltout(),
            .carryin(bfn_4_18_0_),
            .carryout(n12665),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_11_lut_LC_4_18_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_11_lut_LC_4_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_11_lut_LC_4_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_11_lut_LC_4_18_1 (
            .in0(_gnd_net_),
            .in1(N__54346),
            .in2(N__28574),
            .in3(N__25446),
            .lcout(n2192),
            .ltout(),
            .carryin(n12665),
            .carryout(n12666),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_12_lut_LC_4_18_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_12_lut_LC_4_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_12_lut_LC_4_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_12_lut_LC_4_18_2 (
            .in0(_gnd_net_),
            .in1(N__55445),
            .in2(N__28425),
            .in3(N__25443),
            .lcout(n2191),
            .ltout(),
            .carryin(n12666),
            .carryout(n12667),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_13_lut_LC_4_18_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_13_lut_LC_4_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_13_lut_LC_4_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_13_lut_LC_4_18_3 (
            .in0(_gnd_net_),
            .in1(N__54347),
            .in2(N__31199),
            .in3(N__25434),
            .lcout(n2190),
            .ltout(),
            .carryin(n12667),
            .carryout(n12668),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_14_lut_LC_4_18_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_14_lut_LC_4_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_14_lut_LC_4_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_14_lut_LC_4_18_4 (
            .in0(_gnd_net_),
            .in1(N__55446),
            .in2(N__28451),
            .in3(N__25422),
            .lcout(n2189),
            .ltout(),
            .carryin(n12668),
            .carryout(n12669),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_15_lut_LC_4_18_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_15_lut_LC_4_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_15_lut_LC_4_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_15_lut_LC_4_18_5 (
            .in0(_gnd_net_),
            .in1(N__31313),
            .in2(N__55538),
            .in3(N__25419),
            .lcout(n2188),
            .ltout(),
            .carryin(n12669),
            .carryout(n12670),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_16_lut_LC_4_18_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_16_lut_LC_4_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_16_lut_LC_4_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_16_lut_LC_4_18_6 (
            .in0(_gnd_net_),
            .in1(N__33110),
            .in2(N__54731),
            .in3(N__25410),
            .lcout(n2187),
            .ltout(),
            .carryin(n12670),
            .carryout(n12671),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_17_lut_LC_4_18_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_17_lut_LC_4_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_17_lut_LC_4_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_17_lut_LC_4_18_7 (
            .in0(_gnd_net_),
            .in1(N__33227),
            .in2(N__55539),
            .in3(N__25593),
            .lcout(n2186),
            .ltout(),
            .carryin(n12671),
            .carryout(n12672),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_18_lut_LC_4_19_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_18_lut_LC_4_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_18_lut_LC_4_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_18_lut_LC_4_19_0 (
            .in0(_gnd_net_),
            .in1(N__28891),
            .in2(N__55536),
            .in3(N__25590),
            .lcout(n2185),
            .ltout(),
            .carryin(bfn_4_19_0_),
            .carryout(n12673),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_19_lut_LC_4_19_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_19_lut_LC_4_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_19_lut_LC_4_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_19_lut_LC_4_19_1 (
            .in0(_gnd_net_),
            .in1(N__31355),
            .in2(N__54730),
            .in3(N__25587),
            .lcout(n2184),
            .ltout(),
            .carryin(n12673),
            .carryout(n12674),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_20_lut_LC_4_19_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1436_20_lut_LC_4_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_20_lut_LC_4_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1436_20_lut_LC_4_19_2 (
            .in0(_gnd_net_),
            .in1(N__28499),
            .in2(N__55537),
            .in3(N__25584),
            .lcout(n2183),
            .ltout(),
            .carryin(n12674),
            .carryout(n12675),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1436_21_lut_LC_4_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1436_21_lut_LC_4_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1436_21_lut_LC_4_19_3.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1436_21_lut_LC_4_19_3 (
            .in0(N__54345),
            .in1(N__35462),
            .in2(N__31224),
            .in3(N__25581),
            .lcout(n2214),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1518_3_lut_LC_4_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1518_3_lut_LC_4_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1518_3_lut_LC_4_19_4.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1518_3_lut_LC_4_19_4 (
            .in0(N__28246),
            .in1(_gnd_net_),
            .in2(N__25563),
            .in3(N__35540),
            .lcout(n2326),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1442_3_lut_LC_4_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1442_3_lut_LC_4_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1442_3_lut_LC_4_19_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1442_3_lut_LC_4_19_5 (
            .in0(_gnd_net_),
            .in1(N__33228),
            .in2(N__25548),
            .in3(N__35417),
            .lcout(n2218),
            .ltout(n2218_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1509_3_lut_LC_4_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1509_3_lut_LC_4_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1509_3_lut_LC_4_19_6.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1509_3_lut_LC_4_19_6 (
            .in0(N__25518),
            .in1(_gnd_net_),
            .in2(N__25506),
            .in3(N__35541),
            .lcout(n2317),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1444_3_lut_LC_4_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1444_3_lut_LC_4_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1444_3_lut_LC_4_19_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1444_3_lut_LC_4_19_7 (
            .in0(_gnd_net_),
            .in1(N__31314),
            .in2(N__25503),
            .in3(N__35416),
            .lcout(n2220),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_47_LC_4_20_0.C_ON=1'b0;
    defparam i1_4_lut_adj_47_LC_4_20_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_47_LC_4_20_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_47_LC_4_20_0 (
            .in0(N__25723),
            .in1(N__28972),
            .in2(N__29017),
            .in3(N__25818),
            .lcout(),
            .ltout(n14398_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13048_4_lut_LC_4_20_1.C_ON=1'b0;
    defparam i13048_4_lut_LC_4_20_1.SEQ_MODE=4'b0000;
    defparam i13048_4_lut_LC_4_20_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 i13048_4_lut_LC_4_20_1 (
            .in0(N__25805),
            .in1(N__30952),
            .in2(N__25785),
            .in3(N__25688),
            .lcout(n2346),
            .ltout(n2346_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12485_3_lut_LC_4_20_2.C_ON=1'b0;
    defparam i12485_3_lut_LC_4_20_2.SEQ_MODE=4'b0000;
    defparam i12485_3_lut_LC_4_20_2.LUT_INIT=16'b1010111110100000;
    LogicCell40 i12485_3_lut_LC_4_20_2 (
            .in0(N__25778),
            .in1(_gnd_net_),
            .in2(N__25758),
            .in3(N__25755),
            .lcout(n2426),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1508_3_lut_LC_4_20_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1508_3_lut_LC_4_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1508_3_lut_LC_4_20_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1508_3_lut_LC_4_20_3 (
            .in0(_gnd_net_),
            .in1(N__25743),
            .in2(N__28535),
            .in3(N__35566),
            .lcout(n2316),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1506_3_lut_LC_4_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1506_3_lut_LC_4_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1506_3_lut_LC_4_20_4.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1506_3_lut_LC_4_20_4 (
            .in0(_gnd_net_),
            .in1(N__25707),
            .in2(N__35590),
            .in3(N__28483),
            .lcout(n2314),
            .ltout(n2314_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1573_3_lut_LC_4_20_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1573_3_lut_LC_4_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1573_3_lut_LC_4_20_5.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1573_3_lut_LC_4_20_5 (
            .in0(N__35708),
            .in1(_gnd_net_),
            .in2(N__25677),
            .in3(N__25674),
            .lcout(n2413),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1584_3_lut_LC_4_20_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1584_3_lut_LC_4_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1584_3_lut_LC_4_20_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1584_3_lut_LC_4_20_6 (
            .in0(_gnd_net_),
            .in1(N__25662),
            .in2(N__25652),
            .in3(N__35704),
            .lcout(n2424),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1579_3_lut_LC_4_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1579_3_lut_LC_4_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1579_3_lut_LC_4_20_7.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1579_3_lut_LC_4_20_7 (
            .in0(_gnd_net_),
            .in1(N__25622),
            .in2(N__35740),
            .in3(N__25602),
            .lcout(n2419),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1574_3_lut_LC_4_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1574_3_lut_LC_4_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1574_3_lut_LC_4_21_0.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1574_3_lut_LC_4_21_0 (
            .in0(N__25926),
            .in1(_gnd_net_),
            .in2(N__35742),
            .in3(N__30962),
            .lcout(n2414),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1588_3_lut_LC_4_21_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1588_3_lut_LC_4_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1588_3_lut_LC_4_21_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1588_3_lut_LC_4_21_1 (
            .in0(_gnd_net_),
            .in1(N__25917),
            .in2(N__25905),
            .in3(N__35709),
            .lcout(n2428),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1587_3_lut_LC_4_21_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1587_3_lut_LC_4_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1587_3_lut_LC_4_21_2.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1587_3_lut_LC_4_21_2 (
            .in0(_gnd_net_),
            .in1(N__25874),
            .in2(N__35741),
            .in3(N__25848),
            .lcout(n2427),
            .ltout(n2427_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_48_LC_4_21_3.C_ON=1'b0;
    defparam i1_4_lut_adj_48_LC_4_21_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_48_LC_4_21_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_48_LC_4_21_3 (
            .in0(N__33968),
            .in1(N__31798),
            .in2(N__25836),
            .in3(N__31420),
            .lcout(),
            .ltout(n14620_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_49_LC_4_21_4.C_ON=1'b0;
    defparam i1_3_lut_adj_49_LC_4_21_4.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_49_LC_4_21_4.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_49_LC_4_21_4 (
            .in0(_gnd_net_),
            .in1(N__31498),
            .in2(N__25833),
            .in3(N__34102),
            .lcout(n14622),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1654_3_lut_LC_4_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1654_3_lut_LC_4_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1654_3_lut_LC_4_21_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1654_3_lut_LC_4_21_5 (
            .in0(_gnd_net_),
            .in1(N__31464),
            .in2(N__31449),
            .in3(N__35911),
            .lcout(n2526),
            .ltout(n2526_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1721_3_lut_LC_4_21_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1721_3_lut_LC_4_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1721_3_lut_LC_4_21_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1721_3_lut_LC_4_21_6 (
            .in0(_gnd_net_),
            .in1(N__32109),
            .in2(N__25830),
            .in3(N__36097),
            .lcout(n2625),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_4_21_7.C_ON=1'b0;
    defparam i1_2_lut_LC_4_21_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_4_21_7.LUT_INIT=16'b1111000000000000;
    LogicCell40 i1_2_lut_LC_4_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29438),
            .in3(N__29500),
            .lcout(n14816),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1647_3_lut_LC_4_22_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1647_3_lut_LC_4_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1647_3_lut_LC_4_22_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1647_3_lut_LC_4_22_0 (
            .in0(_gnd_net_),
            .in1(N__31710),
            .in2(N__31728),
            .in3(N__35862),
            .lcout(n2519),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1652_3_lut_LC_4_22_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1652_3_lut_LC_4_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1652_3_lut_LC_4_22_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1652_3_lut_LC_4_22_1 (
            .in0(_gnd_net_),
            .in1(N__31404),
            .in2(N__35898),
            .in3(N__31430),
            .lcout(n2524),
            .ltout(n2524_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_154_LC_4_22_2.C_ON=1'b0;
    defparam i1_3_lut_adj_154_LC_4_22_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_154_LC_4_22_2.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_154_LC_4_22_2 (
            .in0(_gnd_net_),
            .in1(N__32189),
            .in2(N__26055),
            .in3(N__32120),
            .lcout(),
            .ltout(n14574_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_159_LC_4_22_3.C_ON=1'b0;
    defparam i1_4_lut_adj_159_LC_4_22_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_159_LC_4_22_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_159_LC_4_22_3 (
            .in0(N__32404),
            .in1(N__26046),
            .in2(N__26052),
            .in3(N__32661),
            .lcout(n14117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1651_3_lut_LC_4_22_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1651_3_lut_LC_4_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1651_3_lut_LC_4_22_4.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1651_3_lut_LC_4_22_4 (
            .in0(N__31808),
            .in1(_gnd_net_),
            .in2(N__31785),
            .in3(N__35861),
            .lcout(n2523),
            .ltout(n2523_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_156_LC_4_22_5.C_ON=1'b0;
    defparam i1_3_lut_adj_156_LC_4_22_5.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_156_LC_4_22_5.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_156_LC_4_22_5 (
            .in0(_gnd_net_),
            .in1(N__32156),
            .in2(N__26049),
            .in3(N__32446),
            .lcout(n14576),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1655_3_lut_LC_4_22_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1655_3_lut_LC_4_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1655_3_lut_LC_4_22_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1655_3_lut_LC_4_22_6 (
            .in0(_gnd_net_),
            .in1(N__31502),
            .in2(N__31482),
            .in3(N__35860),
            .lcout(n2527),
            .ltout(n2527_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1722_3_lut_LC_4_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1722_3_lut_LC_4_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1722_3_lut_LC_4_22_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1722_3_lut_LC_4_22_7 (
            .in0(_gnd_net_),
            .in1(N__32145),
            .in2(N__26040),
            .in3(N__36068),
            .lcout(n2626),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1713_3_lut_LC_4_23_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1713_3_lut_LC_4_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1713_3_lut_LC_4_23_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1713_3_lut_LC_4_23_0 (
            .in0(_gnd_net_),
            .in1(N__33840),
            .in2(N__32370),
            .in3(N__36048),
            .lcout(n2617),
            .ltout(n2617_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_29_LC_4_23_1.C_ON=1'b0;
    defparam i1_3_lut_adj_29_LC_4_23_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_29_LC_4_23_1.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_29_LC_4_23_1 (
            .in0(_gnd_net_),
            .in1(N__25963),
            .in2(N__25935),
            .in3(N__29059),
            .lcout(n14812),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1729_3_lut_LC_4_23_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1729_3_lut_LC_4_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1729_3_lut_LC_4_23_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i1729_3_lut_LC_4_23_2 (
            .in0(N__35145),
            .in1(N__31881),
            .in2(_gnd_net_),
            .in3(N__36044),
            .lcout(n2633),
            .ltout(n2633_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10082_4_lut_LC_4_23_3.C_ON=1'b0;
    defparam i10082_4_lut_LC_4_23_3.SEQ_MODE=4'b0000;
    defparam i10082_4_lut_LC_4_23_3.LUT_INIT=16'b1111111010101010;
    LogicCell40 i10082_4_lut_LC_4_23_3 (
            .in0(N__29182),
            .in1(N__33581),
            .in2(N__26247),
            .in3(N__29239),
            .lcout(n12059),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1714_3_lut_LC_4_23_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1714_3_lut_LC_4_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1714_3_lut_LC_4_23_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1714_3_lut_LC_4_23_4 (
            .in0(_gnd_net_),
            .in1(N__32408),
            .in2(N__32388),
            .in3(N__36049),
            .lcout(n2618),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1710_3_lut_LC_4_23_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1710_3_lut_LC_4_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1710_3_lut_LC_4_23_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1710_3_lut_LC_4_23_5 (
            .in0(N__32858),
            .in1(_gnd_net_),
            .in2(N__36086),
            .in3(N__32844),
            .lcout(n2614),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1709_3_lut_LC_4_23_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1709_3_lut_LC_4_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1709_3_lut_LC_4_23_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1709_3_lut_LC_4_23_6 (
            .in0(_gnd_net_),
            .in1(N__32822),
            .in2(N__32802),
            .in3(N__36050),
            .lcout(n2613),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1715_3_lut_LC_4_23_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1715_3_lut_LC_4_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1715_3_lut_LC_4_23_7.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1715_3_lut_LC_4_23_7 (
            .in0(N__32450),
            .in1(_gnd_net_),
            .in2(N__36085),
            .in3(N__32430),
            .lcout(n2619),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1929_3_lut_LC_4_24_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1929_3_lut_LC_4_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1929_3_lut_LC_4_24_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1929_3_lut_LC_4_24_0 (
            .in0(_gnd_net_),
            .in1(N__26118),
            .in2(N__26540),
            .in3(N__34301),
            .lcout(n2929),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1843_3_lut_LC_4_24_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1843_3_lut_LC_4_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1843_3_lut_LC_4_24_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1843_3_lut_LC_4_24_3 (
            .in0(_gnd_net_),
            .in1(N__26102),
            .in2(N__26082),
            .in3(N__36426),
            .lcout(n2811),
            .ltout(n2811_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1910_3_lut_LC_4_24_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1910_3_lut_LC_4_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1910_3_lut_LC_4_24_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1910_3_lut_LC_4_24_4 (
            .in0(_gnd_net_),
            .in1(N__26067),
            .in2(N__26058),
            .in3(N__34302),
            .lcout(n2910),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1864_3_lut_LC_4_24_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1864_3_lut_LC_4_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1864_3_lut_LC_4_24_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1864_3_lut_LC_4_24_5 (
            .in0(_gnd_net_),
            .in1(N__26618),
            .in2(N__26598),
            .in3(N__36425),
            .lcout(n2832),
            .ltout(n2832_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9976_3_lut_LC_4_24_6.C_ON=1'b0;
    defparam i9976_3_lut_LC_4_24_6.SEQ_MODE=4'b0000;
    defparam i9976_3_lut_LC_4_24_6.LUT_INIT=16'b1111000011000000;
    LogicCell40 i9976_3_lut_LC_4_24_6 (
            .in0(_gnd_net_),
            .in1(N__33496),
            .in2(N__26580),
            .in3(N__26573),
            .lcout(),
            .ltout(n11953_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_64_LC_4_24_7.C_ON=1'b0;
    defparam i1_4_lut_adj_64_LC_4_24_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_64_LC_4_24_7.LUT_INIT=16'b1100100000000000;
    LogicCell40 i1_4_lut_adj_64_LC_4_24_7 (
            .in0(N__29635),
            .in1(N__26533),
            .in2(N__26517),
            .in3(N__29888),
            .lcout(n13857),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_66_LC_4_25_0.C_ON=1'b0;
    defparam i1_4_lut_adj_66_LC_4_25_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_66_LC_4_25_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_66_LC_4_25_0 (
            .in0(N__29774),
            .in1(N__26332),
            .in2(N__26508),
            .in3(N__26478),
            .lcout(),
            .ltout(n14708_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_67_LC_4_25_1.C_ON=1'b0;
    defparam i1_4_lut_adj_67_LC_4_25_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_67_LC_4_25_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_67_LC_4_25_1 (
            .in0(N__26464),
            .in1(N__26434),
            .in2(N__26421),
            .in3(N__26414),
            .lcout(),
            .ltout(n14714_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12626_4_lut_LC_4_25_2.C_ON=1'b0;
    defparam i12626_4_lut_LC_4_25_2.SEQ_MODE=4'b0000;
    defparam i12626_4_lut_LC_4_25_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12626_4_lut_LC_4_25_2 (
            .in0(N__26395),
            .in1(N__26893),
            .in2(N__26370),
            .in3(N__26366),
            .lcout(n2841),
            .ltout(n2841_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1915_3_lut_LC_4_25_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1915_3_lut_LC_4_25_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1915_3_lut_LC_4_25_3.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1915_3_lut_LC_4_25_3 (
            .in0(N__26333),
            .in1(_gnd_net_),
            .in2(N__26319),
            .in3(N__26316),
            .lcout(n2915),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1917_3_lut_LC_4_25_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1917_3_lut_LC_4_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1917_3_lut_LC_4_25_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1917_3_lut_LC_4_25_4 (
            .in0(_gnd_net_),
            .in1(N__26304),
            .in2(N__26291),
            .in3(N__34297),
            .lcout(n2917),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2049_3_lut_LC_4_25_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2049_3_lut_LC_4_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2049_3_lut_LC_4_25_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2049_3_lut_LC_4_25_5 (
            .in0(_gnd_net_),
            .in1(N__26913),
            .in2(N__27461),
            .in3(N__34659),
            .lcout(n3113),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1909_3_lut_LC_4_25_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1909_3_lut_LC_4_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1909_3_lut_LC_4_25_7.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1909_3_lut_LC_4_25_7 (
            .in0(N__26894),
            .in1(_gnd_net_),
            .in2(N__34324),
            .in3(N__26880),
            .lcout(n2909),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1976_3_lut_LC_4_26_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1976_3_lut_LC_4_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1976_3_lut_LC_4_26_0.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1976_3_lut_LC_4_26_0 (
            .in0(N__26971),
            .in1(_gnd_net_),
            .in2(N__26871),
            .in3(N__34479),
            .lcout(n3008),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1918_3_lut_LC_4_26_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1918_3_lut_LC_4_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1918_3_lut_LC_4_26_1.LUT_INIT=16'b1110010011100100;
    LogicCell40 encoder0_position_31__I_0_i1918_3_lut_LC_4_26_1 (
            .in0(N__34290),
            .in1(N__26856),
            .in2(N__26843),
            .in3(_gnd_net_),
            .lcout(n2918),
            .ltout(n2918_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_155_LC_4_26_2.C_ON=1'b0;
    defparam i1_4_lut_adj_155_LC_4_26_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_155_LC_4_26_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_155_LC_4_26_2 (
            .in0(N__26796),
            .in1(N__26773),
            .in2(N__26757),
            .in3(N__29277),
            .lcout(n14216),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1924_3_lut_LC_4_26_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1924_3_lut_LC_4_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1924_3_lut_LC_4_26_3.LUT_INIT=16'b1101100011011000;
    LogicCell40 encoder0_position_31__I_0_i1924_3_lut_LC_4_26_3 (
            .in0(N__34292),
            .in1(N__26754),
            .in2(N__26715),
            .in3(_gnd_net_),
            .lcout(n2924),
            .ltout(n2924_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_69_LC_4_26_4.C_ON=1'b0;
    defparam i1_4_lut_adj_69_LC_4_26_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_69_LC_4_26_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_69_LC_4_26_4 (
            .in0(N__26698),
            .in1(N__26674),
            .in2(N__26658),
            .in3(N__26653),
            .lcout(),
            .ltout(n14212_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_161_LC_4_26_5.C_ON=1'b0;
    defparam i1_4_lut_adj_161_LC_4_26_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_161_LC_4_26_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_161_LC_4_26_5 (
            .in0(N__27196),
            .in1(N__30355),
            .in2(N__26637),
            .in3(N__26634),
            .lcout(n14222),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12622_1_lut_LC_4_26_6.C_ON=1'b0;
    defparam i12622_1_lut_LC_4_26_6.SEQ_MODE=4'b0000;
    defparam i12622_1_lut_LC_4_26_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12622_1_lut_LC_4_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34289),
            .lcout(n15352),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1916_3_lut_LC_4_26_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1916_3_lut_LC_4_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1916_3_lut_LC_4_26_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_i1916_3_lut_LC_4_26_7 (
            .in0(N__34291),
            .in1(N__27243),
            .in2(_gnd_net_),
            .in3(N__27216),
            .lcout(n2916),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1981_3_lut_LC_4_27_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1981_3_lut_LC_4_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1981_3_lut_LC_4_27_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1981_3_lut_LC_4_27_0 (
            .in0(_gnd_net_),
            .in1(N__27092),
            .in2(N__27180),
            .in3(N__34474),
            .lcout(n3013),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_162_LC_4_27_1.C_ON=1'b0;
    defparam i1_4_lut_adj_162_LC_4_27_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_162_LC_4_27_1.LUT_INIT=16'b1111111110000000;
    LogicCell40 i1_4_lut_adj_162_LC_4_27_1 (
            .in0(N__29590),
            .in1(N__30198),
            .in2(N__27166),
            .in3(N__27129),
            .lcout(),
            .ltout(n14224_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_163_LC_4_27_2.C_ON=1'b0;
    defparam i1_4_lut_adj_163_LC_4_27_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_163_LC_4_27_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_163_LC_4_27_2 (
            .in0(N__30286),
            .in1(N__27119),
            .in2(N__27096),
            .in3(N__27091),
            .lcout(),
            .ltout(n14230_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_164_LC_4_27_3.C_ON=1'b0;
    defparam i1_4_lut_adj_164_LC_4_27_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_164_LC_4_27_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_164_LC_4_27_3 (
            .in0(N__27064),
            .in1(N__26935),
            .in2(N__27045),
            .in3(N__27041),
            .lcout(),
            .ltout(n14236_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12658_4_lut_LC_4_27_4.C_ON=1'b0;
    defparam i12658_4_lut_LC_4_27_4.SEQ_MODE=4'b0000;
    defparam i12658_4_lut_LC_4_27_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12658_4_lut_LC_4_27_4 (
            .in0(N__27026),
            .in1(N__27003),
            .in2(N__26982),
            .in3(N__26972),
            .lcout(n2940),
            .ltout(n2940_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1997_3_lut_LC_4_27_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1997_3_lut_LC_4_27_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1997_3_lut_LC_4_27_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1997_3_lut_LC_4_27_5 (
            .in0(N__29591),
            .in1(_gnd_net_),
            .in2(N__26952),
            .in3(N__26949),
            .lcout(n3029),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1978_3_lut_LC_4_27_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1978_3_lut_LC_4_27_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1978_3_lut_LC_4_27_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_i1978_3_lut_LC_4_27_6 (
            .in0(N__26936),
            .in1(N__34475),
            .in2(_gnd_net_),
            .in3(N__26922),
            .lcout(n3010),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1995_3_lut_LC_4_27_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1995_3_lut_LC_4_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1995_3_lut_LC_4_27_7.LUT_INIT=16'b1111101001010000;
    LogicCell40 encoder0_position_31__I_0_i1995_3_lut_LC_4_27_7 (
            .in0(N__34473),
            .in1(_gnd_net_),
            .in2(N__27528),
            .in3(N__29852),
            .lcout(n3027),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2000_3_lut_LC_4_28_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2000_3_lut_LC_4_28_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2000_3_lut_LC_4_28_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2000_3_lut_LC_4_28_0 (
            .in0(_gnd_net_),
            .in1(N__30221),
            .in2(N__27513),
            .in3(N__34462),
            .lcout(n3032),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_170_LC_4_28_1.C_ON=1'b0;
    defparam i1_4_lut_adj_170_LC_4_28_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_170_LC_4_28_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_170_LC_4_28_1 (
            .in0(N__27487),
            .in1(N__30310),
            .in2(N__30528),
            .in3(N__27474),
            .lcout(),
            .ltout(n14742_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_171_LC_4_28_2.C_ON=1'b0;
    defparam i1_4_lut_adj_171_LC_4_28_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_171_LC_4_28_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_171_LC_4_28_2 (
            .in0(N__30238),
            .in1(N__27457),
            .in2(N__27435),
            .in3(N__27574),
            .lcout(),
            .ltout(n14748_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_172_LC_4_28_3.C_ON=1'b0;
    defparam i1_4_lut_adj_172_LC_4_28_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_172_LC_4_28_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_172_LC_4_28_3 (
            .in0(N__27418),
            .in1(N__27394),
            .in2(N__27372),
            .in3(N__28196),
            .lcout(),
            .ltout(n14754_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12691_4_lut_LC_4_28_4.C_ON=1'b0;
    defparam i12691_4_lut_LC_4_28_4.SEQ_MODE=4'b0000;
    defparam i12691_4_lut_LC_4_28_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12691_4_lut_LC_4_28_4 (
            .in0(N__27365),
            .in1(N__27341),
            .in2(N__27327),
            .in3(N__27311),
            .lcout(n3039),
            .ltout(n3039_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2067_3_lut_LC_4_28_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2067_3_lut_LC_4_28_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2067_3_lut_LC_4_28_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2067_3_lut_LC_4_28_5 (
            .in0(_gnd_net_),
            .in1(N__27291),
            .in2(N__27285),
            .in3(N__30077),
            .lcout(n3131),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2053_3_lut_LC_4_29_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2053_3_lut_LC_4_29_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2053_3_lut_LC_4_29_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2053_3_lut_LC_4_29_0 (
            .in0(_gnd_net_),
            .in1(N__27277),
            .in2(N__27252),
            .in3(N__34604),
            .lcout(n3117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2066_3_lut_LC_4_29_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2066_3_lut_LC_4_29_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2066_3_lut_LC_4_29_1.LUT_INIT=16'b1101100011011000;
    LogicCell40 encoder0_position_31__I_0_i2066_3_lut_LC_4_29_1 (
            .in0(N__34612),
            .in1(N__29927),
            .in2(N__27633),
            .in3(_gnd_net_),
            .lcout(n3130),
            .ltout(n3130_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_177_LC_4_29_2.C_ON=1'b0;
    defparam i1_4_lut_adj_177_LC_4_29_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_177_LC_4_29_2.LUT_INIT=16'b1010000010000000;
    LogicCell40 i1_4_lut_adj_177_LC_4_29_2 (
            .in0(N__30484),
            .in1(N__30385),
            .in2(N__27624),
            .in3(N__27600),
            .lcout(n13831),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2069_3_lut_LC_4_29_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2069_3_lut_LC_4_29_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2069_3_lut_LC_4_29_3.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i2069_3_lut_LC_4_29_3 (
            .in0(N__27621),
            .in1(_gnd_net_),
            .in2(N__34657),
            .in3(N__41571),
            .lcout(n3133),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2065_3_lut_LC_4_29_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2065_3_lut_LC_4_29_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2065_3_lut_LC_4_29_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2065_3_lut_LC_4_29_4 (
            .in0(_gnd_net_),
            .in1(N__27615),
            .in2(N__29978),
            .in3(N__34611),
            .lcout(n3129),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2068_3_lut_LC_4_29_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2068_3_lut_LC_4_29_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2068_3_lut_LC_4_29_5.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i2068_3_lut_LC_4_29_5 (
            .in0(_gnd_net_),
            .in1(N__30095),
            .in2(N__34658),
            .in3(N__27609),
            .lcout(n3132),
            .ltout(n3132_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9968_3_lut_LC_4_29_6.C_ON=1'b0;
    defparam i9968_3_lut_LC_4_29_6.SEQ_MODE=4'b0000;
    defparam i9968_3_lut_LC_4_29_6.LUT_INIT=16'b1111000011000000;
    LogicCell40 i9968_3_lut_LC_4_29_6 (
            .in0(_gnd_net_),
            .in1(N__34166),
            .in2(N__27603),
            .in3(N__30421),
            .lcout(n11945),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2048_3_lut_LC_4_29_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2048_3_lut_LC_4_29_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2048_3_lut_LC_4_29_7.LUT_INIT=16'b1110010011100100;
    LogicCell40 encoder0_position_31__I_0_i2048_3_lut_LC_4_29_7 (
            .in0(N__34613),
            .in1(N__27594),
            .in2(N__27588),
            .in3(_gnd_net_),
            .lcout(n3112),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2195_3_lut_LC_4_30_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2195_3_lut_LC_4_30_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2195_3_lut_LC_4_30_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2195_3_lut_LC_4_30_0 (
            .in0(_gnd_net_),
            .in1(N__37152),
            .in2(N__37172),
            .in3(N__35041),
            .lcout(),
            .ltout(n23_adj_715_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_89_LC_4_30_1.C_ON=1'b0;
    defparam i1_4_lut_adj_89_LC_4_30_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_89_LC_4_30_1.LUT_INIT=16'b1111111011110100;
    LogicCell40 i1_4_lut_adj_89_LC_4_30_1 (
            .in0(N__35045),
            .in1(N__36999),
            .in2(N__27558),
            .in3(N__37019),
            .lcout(n14260),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2126_3_lut_LC_4_30_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2126_3_lut_LC_4_30_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2126_3_lut_LC_4_30_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2126_3_lut_LC_4_30_2 (
            .in0(_gnd_net_),
            .in1(N__27555),
            .in2(N__27825),
            .in3(N__34824),
            .lcout(n3222),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2124_3_lut_LC_4_30_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2124_3_lut_LC_4_30_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2124_3_lut_LC_4_30_3.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i2124_3_lut_LC_4_30_3 (
            .in0(_gnd_net_),
            .in1(N__27813),
            .in2(N__34881),
            .in3(N__27786),
            .lcout(n3220),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2128_3_lut_LC_4_30_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2128_3_lut_LC_4_30_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2128_3_lut_LC_4_30_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2128_3_lut_LC_4_30_4 (
            .in0(_gnd_net_),
            .in1(N__27777),
            .in2(N__27768),
            .in3(N__34823),
            .lcout(n3224),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_90_LC_4_30_5.C_ON=1'b0;
    defparam i1_4_lut_adj_90_LC_4_30_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_90_LC_4_30_5.LUT_INIT=16'b1111111110101100;
    LogicCell40 i1_4_lut_adj_90_LC_4_30_5 (
            .in0(N__36677),
            .in1(N__36663),
            .in2(N__35087),
            .in3(N__30756),
            .lcout(n14264),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2130_3_lut_LC_4_30_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2130_3_lut_LC_4_30_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2130_3_lut_LC_4_30_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2130_3_lut_LC_4_30_6 (
            .in0(_gnd_net_),
            .in1(N__27734),
            .in2(N__27705),
            .in3(N__34825),
            .lcout(n3226),
            .ltout(n3226_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_121_LC_4_30_7.C_ON=1'b0;
    defparam i1_4_lut_adj_121_LC_4_30_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_121_LC_4_30_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_121_LC_4_30_7 (
            .in0(N__36712),
            .in1(N__37165),
            .in2(N__27690),
            .in3(N__37090),
            .lcout(n14768),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2122_3_lut_LC_4_31_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2122_3_lut_LC_4_31_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2122_3_lut_LC_4_31_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2122_3_lut_LC_4_31_0 (
            .in0(_gnd_net_),
            .in1(N__27687),
            .in2(N__27663),
            .in3(N__34876),
            .lcout(n3218),
            .ltout(n3218_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_128_LC_4_31_1.C_ON=1'b0;
    defparam i1_3_lut_adj_128_LC_4_31_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_128_LC_4_31_1.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_128_LC_4_31_1 (
            .in0(_gnd_net_),
            .in1(N__37015),
            .in2(N__27648),
            .in3(N__36976),
            .lcout(n14798),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2116_3_lut_LC_4_31_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2116_3_lut_LC_4_31_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2116_3_lut_LC_4_31_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2116_3_lut_LC_4_31_2 (
            .in0(_gnd_net_),
            .in1(N__27881),
            .in2(N__27645),
            .in3(N__34880),
            .lcout(n3212),
            .ltout(n3212_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_131_LC_4_31_3.C_ON=1'b0;
    defparam i1_4_lut_adj_131_LC_4_31_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_131_LC_4_31_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_131_LC_4_31_3 (
            .in0(N__37432),
            .in1(N__37550),
            .in2(N__28086),
            .in3(N__28083),
            .lcout(n14804),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12725_4_lut_LC_4_31_4.C_ON=1'b0;
    defparam i12725_4_lut_LC_4_31_4.SEQ_MODE=4'b0000;
    defparam i12725_4_lut_LC_4_31_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12725_4_lut_LC_4_31_4 (
            .in0(N__28075),
            .in1(N__28057),
            .in2(N__28041),
            .in3(N__27831),
            .lcout(n3138),
            .ltout(n3138_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2131_3_lut_LC_4_31_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2131_3_lut_LC_4_31_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2131_3_lut_LC_4_31_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2131_3_lut_LC_4_31_5 (
            .in0(_gnd_net_),
            .in1(N__28026),
            .in2(N__28014),
            .in3(N__28011),
            .lcout(n3227),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2117_3_lut_LC_4_31_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2117_3_lut_LC_4_31_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2117_3_lut_LC_4_31_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2117_3_lut_LC_4_31_6 (
            .in0(_gnd_net_),
            .in1(N__27915),
            .in2(N__27990),
            .in3(N__34875),
            .lcout(n3213),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2120_3_lut_LC_4_31_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2120_3_lut_LC_4_31_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2120_3_lut_LC_4_31_7.LUT_INIT=16'b1100101011001010;
    LogicCell40 encoder0_position_31__I_0_i2120_3_lut_LC_4_31_7 (
            .in0(N__27978),
            .in1(N__27967),
            .in2(N__34910),
            .in3(_gnd_net_),
            .lcout(n3216),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2051_3_lut_LC_4_32_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2051_3_lut_LC_4_32_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2051_3_lut_LC_4_32_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2051_3_lut_LC_4_32_0 (
            .in0(_gnd_net_),
            .in1(N__30324),
            .in2(N__27939),
            .in3(N__34704),
            .lcout(n3115),
            .ltout(n3115_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_178_LC_4_32_1.C_ON=1'b0;
    defparam i1_4_lut_adj_178_LC_4_32_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_178_LC_4_32_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_178_LC_4_32_1 (
            .in0(N__27924),
            .in1(N__27913),
            .in2(N__27897),
            .in3(N__27894),
            .lcout(),
            .ltout(n14162_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_179_LC_4_32_2.C_ON=1'b0;
    defparam i1_4_lut_adj_179_LC_4_32_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_179_LC_4_32_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_179_LC_4_32_2 (
            .in0(N__30737),
            .in1(N__27877),
            .in2(N__27849),
            .in3(N__31063),
            .lcout(),
            .ltout(n14168_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_180_LC_4_32_3.C_ON=1'b0;
    defparam i1_4_lut_adj_180_LC_4_32_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_180_LC_4_32_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_180_LC_4_32_3 (
            .in0(N__30847),
            .in1(N__31027),
            .in2(N__27846),
            .in3(N__27842),
            .lcout(n14174),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2045_3_lut_LC_4_32_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2045_3_lut_LC_4_32_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2045_3_lut_LC_4_32_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2045_3_lut_LC_4_32_4 (
            .in0(_gnd_net_),
            .in1(N__28209),
            .in2(N__28185),
            .in3(N__34703),
            .lcout(n3109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_95_LC_4_32_6.C_ON=1'b0;
    defparam i1_4_lut_adj_95_LC_4_32_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_95_LC_4_32_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_95_LC_4_32_6 (
            .in0(N__30867),
            .in1(N__28176),
            .in2(N__28167),
            .in3(N__33000),
            .lcout(n14282),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1386_3_lut_LC_5_16_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1386_3_lut_LC_5_16_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1386_3_lut_LC_5_16_0.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1386_3_lut_LC_5_16_0 (
            .in0(_gnd_net_),
            .in1(N__30912),
            .in2(N__35302),
            .in3(N__33345),
            .lcout(n2130),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_30_LC_5_17_0.C_ON=1'b0;
    defparam i1_4_lut_adj_30_LC_5_17_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_30_LC_5_17_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_30_LC_5_17_0 (
            .in0(N__28581),
            .in1(N__33103),
            .in2(N__31312),
            .in3(N__28107),
            .lcout(),
            .ltout(n14324_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_35_LC_5_17_1.C_ON=1'b0;
    defparam i1_4_lut_adj_35_LC_5_17_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_35_LC_5_17_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_35_LC_5_17_1 (
            .in0(N__28895),
            .in1(N__33220),
            .in2(N__28137),
            .in3(N__28134),
            .lcout(n14330),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1383_3_lut_LC_5_17_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1383_3_lut_LC_5_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1383_3_lut_LC_5_17_2.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1383_3_lut_LC_5_17_2 (
            .in0(_gnd_net_),
            .in1(N__31143),
            .in2(N__35303),
            .in3(N__33447),
            .lcout(n2127),
            .ltout(n2127_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_5_17_3.C_ON=1'b0;
    defparam i1_3_lut_LC_5_17_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_5_17_3.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_LC_5_17_3 (
            .in0(_gnd_net_),
            .in1(N__28450),
            .in2(N__28110),
            .in3(N__28573),
            .lcout(n14318),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1387_3_lut_LC_5_17_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1387_3_lut_LC_5_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1387_3_lut_LC_5_17_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1387_3_lut_LC_5_17_5 (
            .in0(_gnd_net_),
            .in1(N__33369),
            .in2(N__30924),
            .in3(N__35292),
            .lcout(n2131),
            .ltout(n2131_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1454_3_lut_LC_5_17_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1454_3_lut_LC_5_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1454_3_lut_LC_5_17_6.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1454_3_lut_LC_5_17_6 (
            .in0(N__28395),
            .in1(_gnd_net_),
            .in2(N__28389),
            .in3(N__35399),
            .lcout(n2230),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_36_LC_5_17_7.C_ON=1'b0;
    defparam i1_2_lut_adj_36_LC_5_17_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_36_LC_5_17_7.LUT_INIT=16'b1111111111110000;
    LogicCell40 i1_2_lut_adj_36_LC_5_17_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28247),
            .in3(N__28288),
            .lcout(n14584),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1447_3_lut_LC_5_18_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1447_3_lut_LC_5_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1447_3_lut_LC_5_18_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1447_3_lut_LC_5_18_0 (
            .in0(_gnd_net_),
            .in1(N__28421),
            .in2(N__28350),
            .in3(N__35379),
            .lcout(n2223),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1382_3_lut_LC_5_18_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1382_3_lut_LC_5_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1382_3_lut_LC_5_18_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1382_3_lut_LC_5_18_1 (
            .in0(_gnd_net_),
            .in1(N__33393),
            .in2(N__31134),
            .in3(N__35258),
            .lcout(n2126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1448_3_lut_LC_5_18_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1448_3_lut_LC_5_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1448_3_lut_LC_5_18_2.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1448_3_lut_LC_5_18_2 (
            .in0(N__28311),
            .in1(_gnd_net_),
            .in2(N__28575),
            .in3(N__35378),
            .lcout(n2224),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1372_3_lut_LC_5_18_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1372_3_lut_LC_5_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1372_3_lut_LC_5_18_3.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1372_3_lut_LC_5_18_3 (
            .in0(N__33180),
            .in1(_gnd_net_),
            .in2(N__31239),
            .in3(N__35262),
            .lcout(n2116),
            .ltout(n2116_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12995_4_lut_LC_5_18_4.C_ON=1'b0;
    defparam i12995_4_lut_LC_5_18_4.SEQ_MODE=4'b0000;
    defparam i12995_4_lut_LC_5_18_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12995_4_lut_LC_5_18_4 (
            .in0(N__31356),
            .in1(N__28272),
            .in2(N__28266),
            .in3(N__31217),
            .lcout(n2148),
            .ltout(n2148_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1451_3_lut_LC_5_18_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1451_3_lut_LC_5_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1451_3_lut_LC_5_18_5.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1451_3_lut_LC_5_18_5 (
            .in0(_gnd_net_),
            .in1(N__28223),
            .in2(N__28263),
            .in3(N__28260),
            .lcout(n2227),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1384_3_lut_LC_5_18_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1384_3_lut_LC_5_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1384_3_lut_LC_5_18_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1384_3_lut_LC_5_18_6 (
            .in0(_gnd_net_),
            .in1(N__31152),
            .in2(N__35288),
            .in3(N__33810),
            .lcout(n2128),
            .ltout(n2128_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_5_18_7.C_ON=1'b0;
    defparam i1_4_lut_LC_5_18_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_5_18_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_LC_5_18_7 (
            .in0(N__28420),
            .in1(N__28600),
            .in2(N__28584),
            .in3(N__31181),
            .lcout(n14316),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1381_3_lut_LC_5_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1381_3_lut_LC_5_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1381_3_lut_LC_5_19_0.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1381_3_lut_LC_5_19_0 (
            .in0(N__31122),
            .in1(_gnd_net_),
            .in2(N__35280),
            .in3(N__33420),
            .lcout(n2125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1441_3_lut_LC_5_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1441_3_lut_LC_5_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1441_3_lut_LC_5_19_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1441_3_lut_LC_5_19_1 (
            .in0(_gnd_net_),
            .in1(N__28548),
            .in2(N__28896),
            .in3(N__35409),
            .lcout(n2217),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1439_3_lut_LC_5_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1439_3_lut_LC_5_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1439_3_lut_LC_5_19_2.LUT_INIT=16'b1100101011001010;
    LogicCell40 encoder0_position_31__I_0_i1439_3_lut_LC_5_19_2 (
            .in0(N__28506),
            .in1(N__28500),
            .in2(N__35441),
            .in3(_gnd_net_),
            .lcout(n2215),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12992_1_lut_LC_5_19_3.C_ON=1'b0;
    defparam i12992_1_lut_LC_5_19_3.SEQ_MODE=4'b0000;
    defparam i12992_1_lut_LC_5_19_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12992_1_lut_LC_5_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35408),
            .lcout(n15722),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1440_3_lut_LC_5_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1440_3_lut_LC_5_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1440_3_lut_LC_5_19_4.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1440_3_lut_LC_5_19_4 (
            .in0(N__28461),
            .in1(_gnd_net_),
            .in2(N__35442),
            .in3(N__31345),
            .lcout(n2216),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1378_3_lut_LC_5_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1378_3_lut_LC_5_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1378_3_lut_LC_5_19_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1378_3_lut_LC_5_19_5 (
            .in0(_gnd_net_),
            .in1(N__31101),
            .in2(N__33270),
            .in3(N__35244),
            .lcout(n2122),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1380_3_lut_LC_5_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1380_3_lut_LC_5_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1380_3_lut_LC_5_19_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1380_3_lut_LC_5_19_6 (
            .in0(_gnd_net_),
            .in1(N__31113),
            .in2(N__35281),
            .in3(N__33465),
            .lcout(n2124),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1593_3_lut_LC_5_20_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1593_3_lut_LC_5_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1593_3_lut_LC_5_20_0.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1593_3_lut_LC_5_20_0 (
            .in0(N__28407),
            .in1(_gnd_net_),
            .in2(N__35738),
            .in3(N__38344),
            .lcout(n2433),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1582_3_lut_LC_5_20_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1582_3_lut_LC_5_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1582_3_lut_LC_5_20_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1582_3_lut_LC_5_20_1 (
            .in0(_gnd_net_),
            .in1(N__28932),
            .in2(N__28923),
            .in3(N__35702),
            .lcout(n2422),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1374_3_lut_LC_5_20_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1374_3_lut_LC_5_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1374_3_lut_LC_5_20_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1374_3_lut_LC_5_20_2 (
            .in0(_gnd_net_),
            .in1(N__31254),
            .in2(N__41272),
            .in3(N__35279),
            .lcout(n2118),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1585_3_lut_LC_5_20_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1585_3_lut_LC_5_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1585_3_lut_LC_5_20_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1585_3_lut_LC_5_20_3 (
            .in0(_gnd_net_),
            .in1(N__28872),
            .in2(N__28859),
            .in3(N__35695),
            .lcout(n2425),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1589_3_lut_LC_5_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1589_3_lut_LC_5_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1589_3_lut_LC_5_20_4.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1589_3_lut_LC_5_20_4 (
            .in0(N__28833),
            .in1(_gnd_net_),
            .in2(N__35739),
            .in3(N__28803),
            .lcout(n2429),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1581_3_lut_LC_5_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1581_3_lut_LC_5_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1581_3_lut_LC_5_20_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1581_3_lut_LC_5_20_7 (
            .in0(_gnd_net_),
            .in1(N__28790),
            .in2(N__28761),
            .in3(N__35703),
            .lcout(n2421),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1591_3_lut_LC_5_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1591_3_lut_LC_5_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1591_3_lut_LC_5_21_0.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1591_3_lut_LC_5_21_0 (
            .in0(_gnd_net_),
            .in1(N__28749),
            .in2(N__35743),
            .in3(N__28736),
            .lcout(n2431),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1580_3_lut_LC_5_21_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1580_3_lut_LC_5_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1580_3_lut_LC_5_21_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1580_3_lut_LC_5_21_1 (
            .in0(_gnd_net_),
            .in1(N__28704),
            .in2(N__28692),
            .in3(N__35723),
            .lcout(n2420),
            .ltout(n2420_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_81_LC_5_21_2.C_ON=1'b0;
    defparam i1_4_lut_adj_81_LC_5_21_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_81_LC_5_21_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_81_LC_5_21_2 (
            .in0(N__31753),
            .in1(N__34030),
            .in2(N__28659),
            .in3(N__28656),
            .lcout(n14628),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1590_3_lut_LC_5_21_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1590_3_lut_LC_5_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1590_3_lut_LC_5_21_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1590_3_lut_LC_5_21_3 (
            .in0(_gnd_net_),
            .in1(N__28650),
            .in2(N__28638),
            .in3(N__35722),
            .lcout(n2430),
            .ltout(n2430_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_82_LC_5_21_4.C_ON=1'b0;
    defparam i1_4_lut_adj_82_LC_5_21_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_82_LC_5_21_4.LUT_INIT=16'b1010000010000000;
    LogicCell40 i1_4_lut_adj_82_LC_5_21_4 (
            .in0(N__31531),
            .in1(N__31606),
            .in2(N__29139),
            .in3(N__29085),
            .lcout(n13828),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1592_3_lut_LC_5_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1592_3_lut_LC_5_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1592_3_lut_LC_5_21_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1592_3_lut_LC_5_21_5 (
            .in0(_gnd_net_),
            .in1(N__29136),
            .in2(N__29124),
            .in3(N__35718),
            .lcout(n2432),
            .ltout(n2432_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9990_3_lut_LC_5_21_6.C_ON=1'b0;
    defparam i9990_3_lut_LC_5_21_6.SEQ_MODE=4'b0000;
    defparam i9990_3_lut_LC_5_21_6.LUT_INIT=16'b1111000010100000;
    LogicCell40 i9990_3_lut_LC_5_21_6 (
            .in0(N__33605),
            .in1(_gnd_net_),
            .in2(N__29088),
            .in3(N__31909),
            .lcout(n11967),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1656_3_lut_LC_5_22_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1656_3_lut_LC_5_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1656_3_lut_LC_5_22_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1656_3_lut_LC_5_22_1 (
            .in0(_gnd_net_),
            .in1(N__31515),
            .in2(N__31542),
            .in3(N__35867),
            .lcout(n2528),
            .ltout(n2528_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1723_3_lut_LC_5_22_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1723_3_lut_LC_5_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1723_3_lut_LC_5_22_2.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1723_3_lut_LC_5_22_2 (
            .in0(N__32178),
            .in1(_gnd_net_),
            .in2(N__29079),
            .in3(N__36057),
            .lcout(n2627),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1576_3_lut_LC_5_22_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1576_3_lut_LC_5_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1576_3_lut_LC_5_22_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1576_3_lut_LC_5_22_3 (
            .in0(_gnd_net_),
            .in1(N__29040),
            .in2(N__29028),
            .in3(N__35746),
            .lcout(n2416),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_149_LC_5_22_4.C_ON=1'b0;
    defparam i1_4_lut_adj_149_LC_5_22_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_149_LC_5_22_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_149_LC_5_22_4 (
            .in0(N__32695),
            .in1(N__28992),
            .in2(N__33871),
            .in3(N__28986),
            .lcout(n14634),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1577_3_lut_LC_5_22_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1577_3_lut_LC_5_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1577_3_lut_LC_5_22_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1577_3_lut_LC_5_22_5 (
            .in0(_gnd_net_),
            .in1(N__28980),
            .in2(N__28947),
            .in3(N__35747),
            .lcout(n2417),
            .ltout(n2417_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1644_3_lut_LC_5_22_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1644_3_lut_LC_5_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1644_3_lut_LC_5_22_6.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1644_3_lut_LC_5_22_6 (
            .in0(N__35868),
            .in1(_gnd_net_),
            .in2(N__29163),
            .in3(N__31680),
            .lcout(n2516),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1659_3_lut_LC_5_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1659_3_lut_LC_5_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1659_3_lut_LC_5_22_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1659_3_lut_LC_5_22_7 (
            .in0(_gnd_net_),
            .in1(N__31623),
            .in2(N__31641),
            .in3(N__35866),
            .lcout(n2531),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_160_LC_5_23_0.C_ON=1'b0;
    defparam i1_4_lut_adj_160_LC_5_23_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_160_LC_5_23_0.LUT_INIT=16'b1111111111101100;
    LogicCell40 i1_4_lut_adj_160_LC_5_23_0 (
            .in0(N__29145),
            .in1(N__32330),
            .in2(N__29268),
            .in3(N__34134),
            .lcout(n14188),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1642_3_lut_LC_5_23_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1642_3_lut_LC_5_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1642_3_lut_LC_5_23_1.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i1642_3_lut_LC_5_23_1 (
            .in0(N__32053),
            .in1(N__32031),
            .in2(N__35897),
            .in3(_gnd_net_),
            .lcout(n2514),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1648_3_lut_LC_5_23_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1648_3_lut_LC_5_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1648_3_lut_LC_5_23_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1648_3_lut_LC_5_23_2 (
            .in0(_gnd_net_),
            .in1(N__31737),
            .in2(N__31764),
            .in3(N__35855),
            .lcout(n2520),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_150_LC_5_23_3.C_ON=1'b0;
    defparam i1_4_lut_adj_150_LC_5_23_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_150_LC_5_23_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_150_LC_5_23_3 (
            .in0(N__31666),
            .in1(N__31691),
            .in2(N__32055),
            .in3(N__29160),
            .lcout(),
            .ltout(n14640_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13075_4_lut_LC_5_23_4.C_ON=1'b0;
    defparam i13075_4_lut_LC_5_23_4.SEQ_MODE=4'b0000;
    defparam i13075_4_lut_LC_5_23_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 i13075_4_lut_LC_5_23_4 (
            .in0(N__31972),
            .in1(N__32008),
            .in2(N__29154),
            .in3(N__31940),
            .lcout(n2445),
            .ltout(n2445_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1657_3_lut_LC_5_23_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1657_3_lut_LC_5_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1657_3_lut_LC_5_23_5.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1657_3_lut_LC_5_23_5 (
            .in0(N__31554),
            .in1(_gnd_net_),
            .in2(N__29151),
            .in3(N__31572),
            .lcout(n2529),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1658_3_lut_LC_5_23_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1658_3_lut_LC_5_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1658_3_lut_LC_5_23_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1658_3_lut_LC_5_23_6 (
            .in0(_gnd_net_),
            .in1(N__31611),
            .in2(N__31587),
            .in3(N__35856),
            .lcout(n2530),
            .ltout(n2530_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_158_LC_5_23_7.C_ON=1'b0;
    defparam i1_2_lut_adj_158_LC_5_23_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_158_LC_5_23_7.LUT_INIT=16'b1111000000000000;
    LogicCell40 i1_2_lut_adj_158_LC_5_23_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29148),
            .in3(N__32233),
            .lcout(n14646),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1661_3_lut_LC_5_24_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1661_3_lut_LC_5_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1661_3_lut_LC_5_24_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1661_3_lut_LC_5_24_0 (
            .in0(N__31278),
            .in1(N__33609),
            .in2(_gnd_net_),
            .in3(N__35870),
            .lcout(n2533),
            .ltout(n2533_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10086_4_lut_LC_5_24_1.C_ON=1'b0;
    defparam i10086_4_lut_LC_5_24_1.SEQ_MODE=4'b0000;
    defparam i10086_4_lut_LC_5_24_1.LUT_INIT=16'b1111111110101000;
    LogicCell40 i10086_4_lut_LC_5_24_1 (
            .in0(N__31834),
            .in1(N__35141),
            .in2(N__29271),
            .in3(N__32305),
            .lcout(n12063),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1728_3_lut_LC_5_24_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1728_3_lut_LC_5_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1728_3_lut_LC_5_24_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1728_3_lut_LC_5_24_2 (
            .in0(_gnd_net_),
            .in1(N__31865),
            .in2(N__31851),
            .in3(N__36011),
            .lcout(n2632),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1640_3_lut_LC_5_24_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1640_3_lut_LC_5_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1640_3_lut_LC_5_24_3.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1640_3_lut_LC_5_24_3 (
            .in0(_gnd_net_),
            .in1(N__31953),
            .in2(N__35899),
            .in3(N__31980),
            .lcout(n2512),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1643_3_lut_LC_5_24_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1643_3_lut_LC_5_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1643_3_lut_LC_5_24_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1643_3_lut_LC_5_24_4 (
            .in0(_gnd_net_),
            .in1(N__31671),
            .in2(N__31650),
            .in3(N__35874),
            .lcout(n2515),
            .ltout(n2515_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_27_LC_5_24_5.C_ON=1'b0;
    defparam i1_4_lut_adj_27_LC_5_24_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_27_LC_5_24_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_27_LC_5_24_5 (
            .in0(N__29220),
            .in1(N__32818),
            .in2(N__29214),
            .in3(N__29211),
            .lcout(),
            .ltout(n14194_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13103_4_lut_LC_5_24_6.C_ON=1'b0;
    defparam i13103_4_lut_LC_5_24_6.SEQ_MODE=4'b0000;
    defparam i13103_4_lut_LC_5_24_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 i13103_4_lut_LC_5_24_6 (
            .in0(N__32780),
            .in1(N__32579),
            .in2(N__29202),
            .in3(N__32750),
            .lcout(n2544),
            .ltout(n2544_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1727_3_lut_LC_5_24_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1727_3_lut_LC_5_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1727_3_lut_LC_5_24_7.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1727_3_lut_LC_5_24_7 (
            .in0(N__31835),
            .in1(_gnd_net_),
            .in2(N__29199),
            .in3(N__31821),
            .lcout(n2631),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1641_3_lut_LC_5_25_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1641_3_lut_LC_5_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1641_3_lut_LC_5_25_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1641_3_lut_LC_5_25_0 (
            .in0(_gnd_net_),
            .in1(N__31992),
            .in2(N__32022),
            .in3(N__35896),
            .lcout(n2513),
            .ltout(n2513_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1708_3_lut_LC_5_25_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1708_3_lut_LC_5_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1708_3_lut_LC_5_25_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1708_3_lut_LC_5_25_1 (
            .in0(N__36031),
            .in1(_gnd_net_),
            .in2(N__29547),
            .in3(N__32769),
            .lcout(n2612),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1725_3_lut_LC_5_25_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1725_3_lut_LC_5_25_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1725_3_lut_LC_5_25_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1725_3_lut_LC_5_25_2 (
            .in0(_gnd_net_),
            .in1(N__32253),
            .in2(N__32274),
            .in3(N__36023),
            .lcout(n2629),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13100_1_lut_LC_5_25_3.C_ON=1'b0;
    defparam i13100_1_lut_LC_5_25_3.SEQ_MODE=4'b0000;
    defparam i13100_1_lut_LC_5_25_3.LUT_INIT=16'b0000111100001111;
    LogicCell40 i13100_1_lut_LC_5_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36070),
            .in3(_gnd_net_),
            .lcout(n15830),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1931_3_lut_LC_5_25_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1931_3_lut_LC_5_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1931_3_lut_LC_5_25_4.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1931_3_lut_LC_5_25_4 (
            .in0(_gnd_net_),
            .in1(N__29472),
            .in2(N__34321),
            .in3(N__29453),
            .lcout(n2931),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1726_3_lut_LC_5_25_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1726_3_lut_LC_5_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1726_3_lut_LC_5_25_5.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1726_3_lut_LC_5_25_5 (
            .in0(N__32283),
            .in1(_gnd_net_),
            .in2(N__36069),
            .in3(N__32306),
            .lcout(n2630),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1716_3_lut_LC_5_25_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1716_3_lut_LC_5_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1716_3_lut_LC_5_25_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1716_3_lut_LC_5_25_6 (
            .in0(_gnd_net_),
            .in1(N__32466),
            .in2(N__34014),
            .in3(N__36030),
            .lcout(n2620),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1933_3_lut_LC_5_25_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1933_3_lut_LC_5_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1933_3_lut_LC_5_25_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i1933_3_lut_LC_5_25_7 (
            .in0(N__33500),
            .in1(N__29352),
            .in2(_gnd_net_),
            .in3(N__34282),
            .lcout(n2933),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1923_3_lut_LC_5_26_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1923_3_lut_LC_5_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1923_3_lut_LC_5_26_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1923_3_lut_LC_5_26_0 (
            .in0(_gnd_net_),
            .in1(N__29340),
            .in2(N__34315),
            .in3(N__29313),
            .lcout(n2923),
            .ltout(n2923_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_68_LC_5_26_1.C_ON=1'b0;
    defparam i1_4_lut_adj_68_LC_5_26_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_68_LC_5_26_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_68_LC_5_26_1 (
            .in0(N__29848),
            .in1(N__29701),
            .in2(N__29280),
            .in3(N__30172),
            .lcout(n14214),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1928_3_lut_LC_5_26_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1928_3_lut_LC_5_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1928_3_lut_LC_5_26_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1928_3_lut_LC_5_26_3 (
            .in0(_gnd_net_),
            .in1(N__29907),
            .in2(N__29895),
            .in3(N__34263),
            .lcout(n2928),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1920_3_lut_LC_5_26_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1920_3_lut_LC_5_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1920_3_lut_LC_5_26_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1920_3_lut_LC_5_26_4 (
            .in0(_gnd_net_),
            .in1(N__29832),
            .in2(N__34314),
            .in3(N__29805),
            .lcout(n2920),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12688_1_lut_LC_5_26_5.C_ON=1'b0;
    defparam i12688_1_lut_LC_5_26_5.SEQ_MODE=4'b0000;
    defparam i12688_1_lut_LC_5_26_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12688_1_lut_LC_5_26_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34660),
            .lcout(n15418),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1913_3_lut_LC_5_26_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1913_3_lut_LC_5_26_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1913_3_lut_LC_5_26_6.LUT_INIT=16'b1110010011100100;
    LogicCell40 encoder0_position_31__I_0_i1913_3_lut_LC_5_26_6 (
            .in0(N__34271),
            .in1(N__29793),
            .in2(N__29781),
            .in3(_gnd_net_),
            .lcout(n2913),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1925_3_lut_LC_5_26_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1925_3_lut_LC_5_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1925_3_lut_LC_5_26_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1925_3_lut_LC_5_26_7 (
            .in0(_gnd_net_),
            .in1(N__29751),
            .in2(N__29739),
            .in3(N__34267),
            .lcout(n2925),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1711_3_lut_LC_5_27_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1711_3_lut_LC_5_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1711_3_lut_LC_5_27_0.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1711_3_lut_LC_5_27_0 (
            .in0(_gnd_net_),
            .in1(N__32319),
            .in2(N__36100),
            .in3(N__32349),
            .lcout(n2615),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1930_3_lut_LC_5_27_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1930_3_lut_LC_5_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1930_3_lut_LC_5_27_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1930_3_lut_LC_5_27_2 (
            .in0(_gnd_net_),
            .in1(N__29648),
            .in2(N__29616),
            .in3(N__34322),
            .lcout(n2930),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1991_3_lut_LC_5_27_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1991_3_lut_LC_5_27_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1991_3_lut_LC_5_27_3.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1991_3_lut_LC_5_27_3 (
            .in0(_gnd_net_),
            .in1(N__29574),
            .in2(N__34504),
            .in3(N__29561),
            .lcout(n3023),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1980_3_lut_LC_5_27_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1980_3_lut_LC_5_27_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1980_3_lut_LC_5_27_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1980_3_lut_LC_5_27_4 (
            .in0(_gnd_net_),
            .in1(N__30290),
            .in2(N__30270),
            .in3(N__34472),
            .lcout(n3012),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10076_4_lut_LC_5_27_5.C_ON=1'b0;
    defparam i10076_4_lut_LC_5_27_5.SEQ_MODE=4'b0000;
    defparam i10076_4_lut_LC_5_27_5.LUT_INIT=16'b1111111011110000;
    LogicCell40 i10076_4_lut_LC_5_27_5 (
            .in0(N__35177),
            .in1(N__30220),
            .in2(N__30008),
            .in3(N__30140),
            .lcout(n12053),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1987_3_lut_LC_5_27_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1987_3_lut_LC_5_27_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1987_3_lut_LC_5_27_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1987_3_lut_LC_5_27_6 (
            .in0(_gnd_net_),
            .in1(N__30192),
            .in2(N__30180),
            .in3(N__34468),
            .lcout(n3019),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1999_3_lut_LC_5_28_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1999_3_lut_LC_5_28_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1999_3_lut_LC_5_28_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1999_3_lut_LC_5_28_0 (
            .in0(_gnd_net_),
            .in1(N__30156),
            .in2(N__30144),
            .in3(N__34466),
            .lcout(n3031),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2001_3_lut_LC_5_28_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2001_3_lut_LC_5_28_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2001_3_lut_LC_5_28_1.LUT_INIT=16'b1100101011001010;
    LogicCell40 encoder0_position_31__I_0_i2001_3_lut_LC_5_28_1 (
            .in0(N__30111),
            .in1(N__35176),
            .in2(N__34503),
            .in3(_gnd_net_),
            .lcout(n3033),
            .ltout(n3033_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9970_3_lut_LC_5_28_2.C_ON=1'b0;
    defparam i9970_3_lut_LC_5_28_2.SEQ_MODE=4'b0000;
    defparam i9970_3_lut_LC_5_28_2.LUT_INIT=16'b1111110000000000;
    LogicCell40 i9970_3_lut_LC_5_28_2 (
            .in0(_gnd_net_),
            .in1(N__41563),
            .in2(N__30081),
            .in3(N__30073),
            .lcout(n11947),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2118_3_lut_LC_5_28_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2118_3_lut_LC_5_28_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2118_3_lut_LC_5_28_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2118_3_lut_LC_5_28_3 (
            .in0(_gnd_net_),
            .in1(N__30057),
            .in2(N__30045),
            .in3(N__34889),
            .lcout(n3214),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1998_3_lut_LC_5_28_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1998_3_lut_LC_5_28_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1998_3_lut_LC_5_28_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1998_3_lut_LC_5_28_4 (
            .in0(_gnd_net_),
            .in1(N__30021),
            .in2(N__30009),
            .in3(N__34467),
            .lcout(n3030),
            .ltout(n3030_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_167_LC_5_28_5.C_ON=1'b0;
    defparam i1_4_lut_adj_167_LC_5_28_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_167_LC_5_28_5.LUT_INIT=16'b1010000010000000;
    LogicCell40 i1_4_lut_adj_167_LC_5_28_5 (
            .in0(N__29947),
            .in1(N__29926),
            .in2(N__30633),
            .in3(N__30630),
            .lcout(),
            .ltout(n13871_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_169_LC_5_28_6.C_ON=1'b0;
    defparam i1_4_lut_adj_169_LC_5_28_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_169_LC_5_28_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_169_LC_5_28_6 (
            .in0(N__30608),
            .in1(N__30580),
            .in2(N__30564),
            .in3(N__30544),
            .lcout(n14078),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2135_3_lut_LC_5_29_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2135_3_lut_LC_5_29_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2135_3_lut_LC_5_29_0.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2135_3_lut_LC_5_29_0 (
            .in0(_gnd_net_),
            .in1(N__30519),
            .in2(N__34915),
            .in3(N__30506),
            .lcout(n3231),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2132_3_lut_LC_5_29_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2132_3_lut_LC_5_29_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2132_3_lut_LC_5_29_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2132_3_lut_LC_5_29_1 (
            .in0(_gnd_net_),
            .in1(N__30488),
            .in2(N__30468),
            .in3(N__34890),
            .lcout(n3228),
            .ltout(n3228_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_125_LC_5_29_2.C_ON=1'b0;
    defparam i1_3_lut_adj_125_LC_5_29_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_125_LC_5_29_2.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_125_LC_5_29_2 (
            .in0(_gnd_net_),
            .in1(N__37129),
            .in2(N__30453),
            .in3(N__30450),
            .lcout(n14770),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2136_3_lut_LC_5_29_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2136_3_lut_LC_5_29_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2136_3_lut_LC_5_29_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2136_3_lut_LC_5_29_3 (
            .in0(_gnd_net_),
            .in1(N__30444),
            .in2(N__30431),
            .in3(N__34891),
            .lcout(n3232),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2134_3_lut_LC_5_29_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2134_3_lut_LC_5_29_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2134_3_lut_LC_5_29_4.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2134_3_lut_LC_5_29_4 (
            .in0(_gnd_net_),
            .in1(N__30405),
            .in2(N__34916),
            .in3(N__30389),
            .lcout(n3230),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1984_3_lut_LC_5_29_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1984_3_lut_LC_5_29_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1984_3_lut_LC_5_29_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1984_3_lut_LC_5_29_5 (
            .in0(_gnd_net_),
            .in1(N__30369),
            .in2(N__30339),
            .in3(N__34505),
            .lcout(n3016),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_129_LC_5_29_7.C_ON=1'b0;
    defparam i1_4_lut_adj_129_LC_5_29_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_129_LC_5_29_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_129_LC_5_29_7 (
            .in0(N__37048),
            .in1(N__37598),
            .in2(N__37211),
            .in3(N__32868),
            .lcout(n14025),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2127_3_lut_LC_5_30_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2127_3_lut_LC_5_30_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2127_3_lut_LC_5_30_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2127_3_lut_LC_5_30_0 (
            .in0(_gnd_net_),
            .in1(N__30816),
            .in2(N__30786),
            .in3(N__34835),
            .lcout(n3223),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12759_4_lut_LC_5_30_1.C_ON=1'b0;
    defparam i12759_4_lut_LC_5_30_1.SEQ_MODE=4'b0000;
    defparam i12759_4_lut_LC_5_30_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12759_4_lut_LC_5_30_1 (
            .in0(N__37639),
            .in1(N__30774),
            .in2(N__30768),
            .in3(N__32973),
            .lcout(n3237),
            .ltout(n3237_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2200_3_lut_LC_5_30_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2200_3_lut_LC_5_30_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2200_3_lut_LC_5_30_2.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2200_3_lut_LC_5_30_2 (
            .in0(_gnd_net_),
            .in1(N__36774),
            .in2(N__30759),
            .in3(N__36801),
            .lcout(n13_adj_713),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2115_3_lut_LC_5_30_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2115_3_lut_LC_5_30_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2115_3_lut_LC_5_30_3.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i2115_3_lut_LC_5_30_3 (
            .in0(N__30750),
            .in1(_gnd_net_),
            .in2(N__34888),
            .in3(N__30730),
            .lcout(n3211),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_126_LC_5_30_4.C_ON=1'b0;
    defparam i1_4_lut_adj_126_LC_5_30_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_126_LC_5_30_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_126_LC_5_30_4 (
            .in0(N__37399),
            .in1(N__37366),
            .in2(N__37472),
            .in3(N__30711),
            .lcout(),
            .ltout(n14776_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_127_LC_5_30_5.C_ON=1'b0;
    defparam i1_4_lut_adj_127_LC_5_30_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_127_LC_5_30_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_127_LC_5_30_5 (
            .in0(N__37273),
            .in1(N__37333),
            .in2(N__30705),
            .in3(N__37247),
            .lcout(n14782),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2125_3_lut_LC_5_30_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2125_3_lut_LC_5_30_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2125_3_lut_LC_5_30_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2125_3_lut_LC_5_30_6 (
            .in0(_gnd_net_),
            .in1(N__30702),
            .in2(N__30681),
            .in3(N__34839),
            .lcout(n3221),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2119_3_lut_LC_5_31_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2119_3_lut_LC_5_31_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2119_3_lut_LC_5_31_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2119_3_lut_LC_5_31_0 (
            .in0(_gnd_net_),
            .in1(N__30669),
            .in2(N__30645),
            .in3(N__34866),
            .lcout(n3215),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2121_3_lut_LC_5_31_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2121_3_lut_LC_5_31_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2121_3_lut_LC_5_31_1.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i2121_3_lut_LC_5_31_1 (
            .in0(N__30903),
            .in1(_gnd_net_),
            .in2(N__34908),
            .in3(N__30894),
            .lcout(n3217),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2193_3_lut_LC_5_31_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2193_3_lut_LC_5_31_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2193_3_lut_LC_5_31_2.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i2193_3_lut_LC_5_31_2 (
            .in0(_gnd_net_),
            .in1(N__37094),
            .in2(N__35088),
            .in3(N__37074),
            .lcout(),
            .ltout(n27_adj_716_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_87_LC_5_31_3.C_ON=1'b0;
    defparam i1_4_lut_adj_87_LC_5_31_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_87_LC_5_31_3.LUT_INIT=16'b1111101011111100;
    LogicCell40 i1_4_lut_adj_87_LC_5_31_3 (
            .in0(N__37471),
            .in1(N__37449),
            .in2(N__30870),
            .in3(N__35050),
            .lcout(n14266),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_91_LC_5_31_4.C_ON=1'b0;
    defparam i1_4_lut_adj_91_LC_5_31_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_91_LC_5_31_4.LUT_INIT=16'b1111111111001010;
    LogicCell40 i1_4_lut_adj_91_LC_5_31_4 (
            .in0(N__36738),
            .in1(N__36758),
            .in2(N__35090),
            .in3(N__30861),
            .lcout(n14268),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2189_3_lut_LC_5_31_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2189_3_lut_LC_5_31_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2189_3_lut_LC_5_31_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2189_3_lut_LC_5_31_5 (
            .in0(_gnd_net_),
            .in1(N__36932),
            .in2(N__36918),
            .in3(N__35049),
            .lcout(n35_adj_719),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2198_3_lut_LC_5_31_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2198_3_lut_LC_5_31_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2198_3_lut_LC_5_31_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2198_3_lut_LC_5_31_6 (
            .in0(_gnd_net_),
            .in1(N__36696),
            .in2(N__35089),
            .in3(N__36716),
            .lcout(),
            .ltout(n17_adj_714_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_93_LC_5_31_7.C_ON=1'b0;
    defparam i1_4_lut_adj_93_LC_5_31_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_93_LC_5_31_7.LUT_INIT=16'b1111110011111010;
    LogicCell40 i1_4_lut_adj_93_LC_5_31_7 (
            .in0(N__37416),
            .in1(N__37436),
            .in2(N__30855),
            .in3(N__35057),
            .lcout(n14272),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2112_3_lut_LC_5_32_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2112_3_lut_LC_5_32_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2112_3_lut_LC_5_32_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2112_3_lut_LC_5_32_0 (
            .in0(_gnd_net_),
            .in1(N__30851),
            .in2(N__30831),
            .in3(N__34874),
            .lcout(n3208),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2190_3_lut_LC_5_32_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2190_3_lut_LC_5_32_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2190_3_lut_LC_5_32_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2190_3_lut_LC_5_32_3 (
            .in0(_gnd_net_),
            .in1(N__36986),
            .in2(N__36954),
            .in3(N__35091),
            .lcout(),
            .ltout(n33_adj_718_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_94_LC_5_32_4.C_ON=1'b0;
    defparam i1_4_lut_adj_94_LC_5_32_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_94_LC_5_32_4.LUT_INIT=16'b1111111011110100;
    LogicCell40 i1_4_lut_adj_94_LC_5_32_4 (
            .in0(N__35092),
            .in1(N__37113),
            .in2(N__30819),
            .in3(N__37139),
            .lcout(),
            .ltout(n14262_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_97_LC_5_32_5.C_ON=1'b0;
    defparam i1_4_lut_adj_97_LC_5_32_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_97_LC_5_32_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_97_LC_5_32_5 (
            .in0(N__31089),
            .in1(N__31083),
            .in2(N__31077),
            .in3(N__31074),
            .lcout(n14284),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2114_3_lut_LC_5_32_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2114_3_lut_LC_5_32_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2114_3_lut_LC_5_32_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2114_3_lut_LC_5_32_6 (
            .in0(_gnd_net_),
            .in1(N__31068),
            .in2(N__31047),
            .in3(N__34870),
            .lcout(n3210),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2113_3_lut_LC_5_32_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2113_3_lut_LC_5_32_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2113_3_lut_LC_5_32_7.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i2113_3_lut_LC_5_32_7 (
            .in0(_gnd_net_),
            .in1(N__31032),
            .in2(N__34909),
            .in3(N__31011),
            .lcout(n3209),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1507_3_lut_LC_6_16_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1507_3_lut_LC_6_16_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1507_3_lut_LC_6_16_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1507_3_lut_LC_6_16_1 (
            .in0(_gnd_net_),
            .in1(N__31002),
            .in2(N__30993),
            .in3(N__35597),
            .lcout(n2315),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_2_lut_LC_6_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_2_lut_LC_6_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_2_lut_LC_6_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_2_lut_LC_6_17_0 (
            .in0(_gnd_net_),
            .in1(N__38087),
            .in2(_gnd_net_),
            .in3(N__30930),
            .lcout(n2101),
            .ltout(),
            .carryin(bfn_6_17_0_),
            .carryout(n12639),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_3_lut_LC_6_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_3_lut_LC_6_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_3_lut_LC_6_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_3_lut_LC_6_17_1 (
            .in0(_gnd_net_),
            .in1(N__55346),
            .in2(N__33732),
            .in3(N__30927),
            .lcout(n2100),
            .ltout(),
            .carryin(n12639),
            .carryout(n12640),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_4_lut_LC_6_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_4_lut_LC_6_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_4_lut_LC_6_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_4_lut_LC_6_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33368),
            .in3(N__30915),
            .lcout(n2099),
            .ltout(),
            .carryin(n12640),
            .carryout(n12641),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_5_lut_LC_6_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_5_lut_LC_6_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_5_lut_LC_6_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_5_lut_LC_6_17_3 (
            .in0(_gnd_net_),
            .in1(N__55347),
            .in2(N__33341),
            .in3(N__30906),
            .lcout(n2098),
            .ltout(),
            .carryin(n12641),
            .carryout(n12642),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_6_lut_LC_6_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_6_lut_LC_6_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_6_lut_LC_6_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_6_lut_LC_6_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33776),
            .in3(N__31155),
            .lcout(n2097),
            .ltout(),
            .carryin(n12642),
            .carryout(n12643),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_7_lut_LC_6_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_7_lut_LC_6_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_7_lut_LC_6_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_7_lut_LC_6_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33806),
            .in3(N__31146),
            .lcout(n2096),
            .ltout(),
            .carryin(n12643),
            .carryout(n12644),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_8_lut_LC_6_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_8_lut_LC_6_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_8_lut_LC_6_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_8_lut_LC_6_17_6 (
            .in0(_gnd_net_),
            .in1(N__55045),
            .in2(N__33443),
            .in3(N__31137),
            .lcout(n2095),
            .ltout(),
            .carryin(n12644),
            .carryout(n12645),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_9_lut_LC_6_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_9_lut_LC_6_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_9_lut_LC_6_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_9_lut_LC_6_17_7 (
            .in0(_gnd_net_),
            .in1(N__55348),
            .in2(N__33392),
            .in3(N__31125),
            .lcout(n2094),
            .ltout(),
            .carryin(n12645),
            .carryout(n12646),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_10_lut_LC_6_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_10_lut_LC_6_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_10_lut_LC_6_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_10_lut_LC_6_18_0 (
            .in0(_gnd_net_),
            .in1(N__55157),
            .in2(N__33419),
            .in3(N__31116),
            .lcout(n2093),
            .ltout(),
            .carryin(bfn_6_18_0_),
            .carryout(n12647),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_11_lut_LC_6_18_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_11_lut_LC_6_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_11_lut_LC_6_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_11_lut_LC_6_18_1 (
            .in0(_gnd_net_),
            .in1(N__55160),
            .in2(N__33464),
            .in3(N__31107),
            .lcout(n2092),
            .ltout(),
            .carryin(n12647),
            .carryout(n12648),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_12_lut_LC_6_18_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_12_lut_LC_6_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_12_lut_LC_6_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_12_lut_LC_6_18_2 (
            .in0(_gnd_net_),
            .in1(N__33287),
            .in2(N__55345),
            .in3(N__31104),
            .lcout(n2091),
            .ltout(),
            .carryin(n12648),
            .carryout(n12649),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_13_lut_LC_6_18_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_13_lut_LC_6_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_13_lut_LC_6_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_13_lut_LC_6_18_3 (
            .in0(_gnd_net_),
            .in1(N__55164),
            .in2(N__33269),
            .in3(N__31095),
            .lcout(n2090),
            .ltout(),
            .carryin(n12649),
            .carryout(n12650),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_14_lut_LC_6_18_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_14_lut_LC_6_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_14_lut_LC_6_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_14_lut_LC_6_18_4 (
            .in0(_gnd_net_),
            .in1(N__55158),
            .in2(N__33314),
            .in3(N__31092),
            .lcout(n2089),
            .ltout(),
            .carryin(n12650),
            .carryout(n12651),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_15_lut_LC_6_18_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_15_lut_LC_6_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_15_lut_LC_6_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_15_lut_LC_6_18_5 (
            .in0(_gnd_net_),
            .in1(N__55165),
            .in2(N__33141),
            .in3(N__31260),
            .lcout(n2088),
            .ltout(),
            .carryin(n12651),
            .carryout(n12652),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_16_lut_LC_6_18_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_16_lut_LC_6_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_16_lut_LC_6_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_16_lut_LC_6_18_6 (
            .in0(_gnd_net_),
            .in1(N__55159),
            .in2(N__33084),
            .in3(N__31257),
            .lcout(n2087),
            .ltout(),
            .carryin(n12652),
            .carryout(n12653),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_17_lut_LC_6_18_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_17_lut_LC_6_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_17_lut_LC_6_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_17_lut_LC_6_18_7 (
            .in0(_gnd_net_),
            .in1(N__55166),
            .in2(N__41274),
            .in3(N__31245),
            .lcout(n2086),
            .ltout(),
            .carryin(n12653),
            .carryout(n12654),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_18_lut_LC_6_19_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_18_lut_LC_6_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_18_lut_LC_6_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_18_lut_LC_6_19_0 (
            .in0(_gnd_net_),
            .in1(N__31377),
            .in2(N__55490),
            .in3(N__31242),
            .lcout(n2085),
            .ltout(),
            .carryin(bfn_6_19_0_),
            .carryout(n12655),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_19_lut_LC_6_19_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1369_19_lut_LC_6_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_19_lut_LC_6_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1369_19_lut_LC_6_19_1 (
            .in0(_gnd_net_),
            .in1(N__33176),
            .in2(N__55240),
            .in3(N__31230),
            .lcout(n2084),
            .ltout(),
            .carryin(n12655),
            .carryout(n12656),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1369_20_lut_LC_6_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1369_20_lut_LC_6_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1369_20_lut_LC_6_19_2.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1369_20_lut_LC_6_19_2 (
            .in0(N__55344),
            .in1(N__35315),
            .in2(N__37929),
            .in3(N__31227),
            .lcout(n2115),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1379_3_lut_LC_6_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1379_3_lut_LC_6_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1379_3_lut_LC_6_19_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1379_3_lut_LC_6_19_3 (
            .in0(_gnd_net_),
            .in1(N__31206),
            .in2(N__33291),
            .in3(N__35257),
            .lcout(n2123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_148_LC_6_19_4.C_ON=1'b0;
    defparam i1_4_lut_adj_148_LC_6_19_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_148_LC_6_19_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_148_LC_6_19_4 (
            .in0(N__33140),
            .in1(N__33083),
            .in2(N__41273),
            .in3(N__33750),
            .lcout(),
            .ltout(n14558_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12970_4_lut_LC_6_19_5.C_ON=1'b0;
    defparam i12970_4_lut_LC_6_19_5.SEQ_MODE=4'b0000;
    defparam i12970_4_lut_LC_6_19_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12970_4_lut_LC_6_19_5 (
            .in0(N__31376),
            .in1(N__33175),
            .in2(N__31392),
            .in3(N__37925),
            .lcout(n2049),
            .ltout(n2049_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1389_3_lut_LC_6_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1389_3_lut_LC_6_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1389_3_lut_LC_6_19_6.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1389_3_lut_LC_6_19_6 (
            .in0(N__31389),
            .in1(_gnd_net_),
            .in2(N__31380),
            .in3(N__38088),
            .lcout(n2133),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1311_3_lut_LC_6_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1311_3_lut_LC_6_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1311_3_lut_LC_6_19_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1311_3_lut_LC_6_19_7 (
            .in0(_gnd_net_),
            .in1(N__38064),
            .in2(N__41132),
            .in3(N__41359),
            .lcout(n2023),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12967_1_lut_LC_6_20_0.C_ON=1'b0;
    defparam i12967_1_lut_LC_6_20_0.SEQ_MODE=4'b0000;
    defparam i12967_1_lut_LC_6_20_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12967_1_lut_LC_6_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35277),
            .lcout(n15697),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1306_3_lut_LC_6_20_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1306_3_lut_LC_6_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1306_3_lut_LC_6_20_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1306_3_lut_LC_6_20_2 (
            .in0(_gnd_net_),
            .in1(N__38142),
            .in2(N__37986),
            .in3(N__41374),
            .lcout(n2018),
            .ltout(n2018_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1373_3_lut_LC_6_20_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1373_3_lut_LC_6_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1373_3_lut_LC_6_20_3.LUT_INIT=16'b1110010011100100;
    LogicCell40 encoder0_position_31__I_0_i1373_3_lut_LC_6_20_3 (
            .in0(N__35278),
            .in1(N__31365),
            .in2(N__31359),
            .in3(_gnd_net_),
            .lcout(n2117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1377_3_lut_LC_6_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1377_3_lut_LC_6_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1377_3_lut_LC_6_20_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1377_3_lut_LC_6_20_4 (
            .in0(_gnd_net_),
            .in1(N__31323),
            .in2(N__33315),
            .in3(N__35276),
            .lcout(n2121),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_2_lut_LC_6_21_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_2_lut_LC_6_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_2_lut_LC_6_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_2_lut_LC_6_21_0 (
            .in0(_gnd_net_),
            .in1(N__33601),
            .in2(_gnd_net_),
            .in3(N__31266),
            .lcout(n2501),
            .ltout(),
            .carryin(bfn_6_21_0_),
            .carryout(n12717),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_3_lut_LC_6_21_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_3_lut_LC_6_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_3_lut_LC_6_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_3_lut_LC_6_21_1 (
            .in0(_gnd_net_),
            .in1(N__54787),
            .in2(N__31916),
            .in3(N__31263),
            .lcout(n2500),
            .ltout(),
            .carryin(n12717),
            .carryout(n12718),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_4_lut_LC_6_21_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_4_lut_LC_6_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_4_lut_LC_6_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_4_lut_LC_6_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31640),
            .in3(N__31614),
            .lcout(n2499),
            .ltout(),
            .carryin(n12718),
            .carryout(n12719),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_5_lut_LC_6_21_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_5_lut_LC_6_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_5_lut_LC_6_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_5_lut_LC_6_21_3 (
            .in0(_gnd_net_),
            .in1(N__54788),
            .in2(N__31610),
            .in3(N__31575),
            .lcout(n2498),
            .ltout(),
            .carryin(n12719),
            .carryout(n12720),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_6_lut_LC_6_21_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_6_lut_LC_6_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_6_lut_LC_6_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_6_lut_LC_6_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31571),
            .in3(N__31545),
            .lcout(n2497),
            .ltout(),
            .carryin(n12720),
            .carryout(n12721),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_7_lut_LC_6_21_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_7_lut_LC_6_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_7_lut_LC_6_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_7_lut_LC_6_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31538),
            .in3(N__31509),
            .lcout(n2496),
            .ltout(),
            .carryin(n12721),
            .carryout(n12722),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_8_lut_LC_6_21_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_8_lut_LC_6_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_8_lut_LC_6_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_8_lut_LC_6_21_6 (
            .in0(_gnd_net_),
            .in1(N__54763),
            .in2(N__31506),
            .in3(N__31467),
            .lcout(n2495),
            .ltout(),
            .carryin(n12722),
            .carryout(n12723),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_9_lut_LC_6_21_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_9_lut_LC_6_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_9_lut_LC_6_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_9_lut_LC_6_21_7 (
            .in0(_gnd_net_),
            .in1(N__31463),
            .in2(N__55041),
            .in3(N__31437),
            .lcout(n2494),
            .ltout(),
            .carryin(n12723),
            .carryout(n12724),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_10_lut_LC_6_22_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_10_lut_LC_6_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_10_lut_LC_6_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_10_lut_LC_6_22_0 (
            .in0(_gnd_net_),
            .in1(N__54756),
            .in2(N__33984),
            .in3(N__31434),
            .lcout(n2493),
            .ltout(),
            .carryin(bfn_6_22_0_),
            .carryout(n12725),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_11_lut_LC_6_22_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_11_lut_LC_6_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_11_lut_LC_6_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_11_lut_LC_6_22_1 (
            .in0(_gnd_net_),
            .in1(N__54784),
            .in2(N__31431),
            .in3(N__31395),
            .lcout(n2492),
            .ltout(),
            .carryin(n12725),
            .carryout(n12726),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_12_lut_LC_6_22_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_12_lut_LC_6_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_12_lut_LC_6_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_12_lut_LC_6_22_2 (
            .in0(_gnd_net_),
            .in1(N__54757),
            .in2(N__31812),
            .in3(N__31773),
            .lcout(n2491),
            .ltout(),
            .carryin(n12726),
            .carryout(n12727),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_13_lut_LC_6_22_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_13_lut_LC_6_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_13_lut_LC_6_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_13_lut_LC_6_22_3 (
            .in0(_gnd_net_),
            .in1(N__54785),
            .in2(N__34119),
            .in3(N__31770),
            .lcout(n2490),
            .ltout(),
            .carryin(n12727),
            .carryout(n12728),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_14_lut_LC_6_22_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_14_lut_LC_6_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_14_lut_LC_6_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_14_lut_LC_6_22_4 (
            .in0(_gnd_net_),
            .in1(N__54758),
            .in2(N__34043),
            .in3(N__31767),
            .lcout(n2489),
            .ltout(),
            .carryin(n12728),
            .carryout(n12729),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_15_lut_LC_6_22_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_15_lut_LC_6_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_15_lut_LC_6_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_15_lut_LC_6_22_5 (
            .in0(_gnd_net_),
            .in1(N__31760),
            .in2(N__55040),
            .in3(N__31731),
            .lcout(n2488),
            .ltout(),
            .carryin(n12729),
            .carryout(n12730),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_16_lut_LC_6_22_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_16_lut_LC_6_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_16_lut_LC_6_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_16_lut_LC_6_22_6 (
            .in0(_gnd_net_),
            .in1(N__54762),
            .in2(N__31727),
            .in3(N__31701),
            .lcout(n2487),
            .ltout(),
            .carryin(n12730),
            .carryout(n12731),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_17_lut_LC_6_22_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_17_lut_LC_6_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_17_lut_LC_6_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_17_lut_LC_6_22_7 (
            .in0(_gnd_net_),
            .in1(N__54786),
            .in2(N__33878),
            .in3(N__31698),
            .lcout(n2486),
            .ltout(),
            .carryin(n12731),
            .carryout(n12732),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_18_lut_LC_6_23_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_18_lut_LC_6_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_18_lut_LC_6_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_18_lut_LC_6_23_0 (
            .in0(_gnd_net_),
            .in1(N__54746),
            .in2(N__32702),
            .in3(N__31695),
            .lcout(n2485),
            .ltout(),
            .carryin(bfn_6_23_0_),
            .carryout(n12733),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_19_lut_LC_6_23_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_19_lut_LC_6_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_19_lut_LC_6_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_19_lut_LC_6_23_1 (
            .in0(_gnd_net_),
            .in1(N__31692),
            .in2(N__55037),
            .in3(N__31674),
            .lcout(n2484),
            .ltout(),
            .carryin(n12733),
            .carryout(n12734),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_20_lut_LC_6_23_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_20_lut_LC_6_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_20_lut_LC_6_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_20_lut_LC_6_23_2 (
            .in0(_gnd_net_),
            .in1(N__31667),
            .in2(N__55055),
            .in3(N__32058),
            .lcout(n2483),
            .ltout(),
            .carryin(n12734),
            .carryout(n12735),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_21_lut_LC_6_23_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_21_lut_LC_6_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_21_lut_LC_6_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_21_lut_LC_6_23_3 (
            .in0(_gnd_net_),
            .in1(N__32054),
            .in2(N__55038),
            .in3(N__32025),
            .lcout(n2482),
            .ltout(),
            .carryin(n12735),
            .carryout(n12736),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_22_lut_LC_6_23_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_22_lut_LC_6_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_22_lut_LC_6_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_22_lut_LC_6_23_4 (
            .in0(_gnd_net_),
            .in1(N__32015),
            .in2(N__55056),
            .in3(N__31983),
            .lcout(n2481),
            .ltout(),
            .carryin(n12736),
            .carryout(n12737),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_23_lut_LC_6_23_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1637_23_lut_LC_6_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_23_lut_LC_6_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1637_23_lut_LC_6_23_5 (
            .in0(_gnd_net_),
            .in1(N__31979),
            .in2(N__55039),
            .in3(N__31947),
            .lcout(n2480),
            .ltout(),
            .carryin(n12737),
            .carryout(n12738),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1637_24_lut_LC_6_23_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1637_24_lut_LC_6_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1637_24_lut_LC_6_23_6.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1637_24_lut_LC_6_23_6 (
            .in0(N__54783),
            .in1(N__31944),
            .in2(N__35948),
            .in3(N__31923),
            .lcout(n2511),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1660_3_lut_LC_6_23_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1660_3_lut_LC_6_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1660_3_lut_LC_6_23_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1660_3_lut_LC_6_23_7 (
            .in0(_gnd_net_),
            .in1(N__31920),
            .in2(N__31893),
            .in3(N__35869),
            .lcout(n2532),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_2_lut_LC_6_24_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_2_lut_LC_6_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_2_lut_LC_6_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_2_lut_LC_6_24_0 (
            .in0(_gnd_net_),
            .in1(N__35137),
            .in2(_gnd_net_),
            .in3(N__31869),
            .lcout(n2601),
            .ltout(),
            .carryin(bfn_6_24_0_),
            .carryout(n12739),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_3_lut_LC_6_24_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_3_lut_LC_6_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_3_lut_LC_6_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_3_lut_LC_6_24_1 (
            .in0(_gnd_net_),
            .in1(N__53816),
            .in2(N__31866),
            .in3(N__31842),
            .lcout(n2600),
            .ltout(),
            .carryin(n12739),
            .carryout(n12740),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_4_lut_LC_6_24_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_4_lut_LC_6_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_4_lut_LC_6_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_4_lut_LC_6_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31839),
            .in3(N__31815),
            .lcout(n2599),
            .ltout(),
            .carryin(n12740),
            .carryout(n12741),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_5_lut_LC_6_24_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_5_lut_LC_6_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_5_lut_LC_6_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_5_lut_LC_6_24_3 (
            .in0(_gnd_net_),
            .in1(N__53817),
            .in2(N__32310),
            .in3(N__32277),
            .lcout(n2598),
            .ltout(),
            .carryin(n12741),
            .carryout(n12742),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_6_lut_LC_6_24_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_6_lut_LC_6_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_6_lut_LC_6_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_6_lut_LC_6_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32270),
            .in3(N__32247),
            .lcout(n2597),
            .ltout(),
            .carryin(n12742),
            .carryout(n12743),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_7_lut_LC_6_24_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_7_lut_LC_6_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_7_lut_LC_6_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_7_lut_LC_6_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32240),
            .in3(N__32202),
            .lcout(n2596),
            .ltout(),
            .carryin(n12743),
            .carryout(n12744),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_8_lut_LC_6_24_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_8_lut_LC_6_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_8_lut_LC_6_24_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_8_lut_LC_6_24_6 (
            .in0(_gnd_net_),
            .in1(N__53819),
            .in2(N__32199),
            .in3(N__32169),
            .lcout(n2595),
            .ltout(),
            .carryin(n12744),
            .carryout(n12745),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_9_lut_LC_6_24_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_9_lut_LC_6_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_9_lut_LC_6_24_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_9_lut_LC_6_24_7 (
            .in0(_gnd_net_),
            .in1(N__53818),
            .in2(N__32166),
            .in3(N__32133),
            .lcout(n2594),
            .ltout(),
            .carryin(n12745),
            .carryout(n12746),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_10_lut_LC_6_25_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_10_lut_LC_6_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_10_lut_LC_6_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_10_lut_LC_6_25_0 (
            .in0(_gnd_net_),
            .in1(N__54506),
            .in2(N__32130),
            .in3(N__32097),
            .lcout(n2593),
            .ltout(),
            .carryin(bfn_6_25_0_),
            .carryout(n12747),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_11_lut_LC_6_25_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_11_lut_LC_6_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_11_lut_LC_6_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_11_lut_LC_6_25_1 (
            .in0(_gnd_net_),
            .in1(N__54417),
            .in2(N__33951),
            .in3(N__32094),
            .lcout(n2592),
            .ltout(),
            .carryin(n12747),
            .carryout(n12748),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_12_lut_LC_6_25_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_12_lut_LC_6_25_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_12_lut_LC_6_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_12_lut_LC_6_25_2 (
            .in0(_gnd_net_),
            .in1(N__32091),
            .in2(N__54776),
            .in3(N__32523),
            .lcout(n2591),
            .ltout(),
            .carryin(n12748),
            .carryout(n12749),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_13_lut_LC_6_25_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_13_lut_LC_6_25_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_13_lut_LC_6_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_13_lut_LC_6_25_3 (
            .in0(_gnd_net_),
            .in1(N__54421),
            .in2(N__32520),
            .in3(N__32487),
            .lcout(n2590),
            .ltout(),
            .carryin(n12749),
            .carryout(n12750),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_14_lut_LC_6_25_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_14_lut_LC_6_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_14_lut_LC_6_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_14_lut_LC_6_25_4 (
            .in0(_gnd_net_),
            .in1(N__54507),
            .in2(N__34082),
            .in3(N__32469),
            .lcout(n2589),
            .ltout(),
            .carryin(n12750),
            .carryout(n12751),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_15_lut_LC_6_25_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_15_lut_LC_6_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_15_lut_LC_6_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_15_lut_LC_6_25_5 (
            .in0(_gnd_net_),
            .in1(N__54422),
            .in2(N__34010),
            .in3(N__32457),
            .lcout(n2588),
            .ltout(),
            .carryin(n12751),
            .carryout(n12752),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_16_lut_LC_6_25_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_16_lut_LC_6_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_16_lut_LC_6_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_16_lut_LC_6_25_6 (
            .in0(_gnd_net_),
            .in1(N__54508),
            .in2(N__32454),
            .in3(N__32418),
            .lcout(n2587),
            .ltout(),
            .carryin(n12752),
            .carryout(n12753),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_17_lut_LC_6_25_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_17_lut_LC_6_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_17_lut_LC_6_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_17_lut_LC_6_25_7 (
            .in0(_gnd_net_),
            .in1(N__54423),
            .in2(N__32415),
            .in3(N__32373),
            .lcout(n2586),
            .ltout(),
            .carryin(n12753),
            .carryout(n12754),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_18_lut_LC_6_26_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_18_lut_LC_6_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_18_lut_LC_6_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_18_lut_LC_6_26_0 (
            .in0(_gnd_net_),
            .in1(N__33839),
            .in2(N__54744),
            .in3(N__32355),
            .lcout(n2585),
            .ltout(),
            .carryin(bfn_6_26_0_),
            .carryout(n12755),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_19_lut_LC_6_26_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_19_lut_LC_6_26_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_19_lut_LC_6_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_19_lut_LC_6_26_1 (
            .in0(_gnd_net_),
            .in1(N__54373),
            .in2(N__32657),
            .in3(N__32352),
            .lcout(n2584),
            .ltout(),
            .carryin(n12755),
            .carryout(n12756),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_20_lut_LC_6_26_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_20_lut_LC_6_26_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_20_lut_LC_6_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_20_lut_LC_6_26_2 (
            .in0(_gnd_net_),
            .in1(N__54379),
            .in2(N__32348),
            .in3(N__32313),
            .lcout(n2583),
            .ltout(),
            .carryin(n12756),
            .carryout(n12757),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_21_lut_LC_6_26_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_21_lut_LC_6_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_21_lut_LC_6_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_21_lut_LC_6_26_3 (
            .in0(_gnd_net_),
            .in1(N__54374),
            .in2(N__32862),
            .in3(N__32832),
            .lcout(n2582),
            .ltout(),
            .carryin(n12757),
            .carryout(n12758),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_22_lut_LC_6_26_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_22_lut_LC_6_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_22_lut_LC_6_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_22_lut_LC_6_26_4 (
            .in0(_gnd_net_),
            .in1(N__54380),
            .in2(N__32829),
            .in3(N__32787),
            .lcout(n2581),
            .ltout(),
            .carryin(n12758),
            .carryout(n12759),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_23_lut_LC_6_26_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_23_lut_LC_6_26_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_23_lut_LC_6_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_23_lut_LC_6_26_5 (
            .in0(_gnd_net_),
            .in1(N__54375),
            .in2(N__32784),
            .in3(N__32763),
            .lcout(n2580),
            .ltout(),
            .carryin(n12759),
            .carryout(n12760),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_24_lut_LC_6_26_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1704_24_lut_LC_6_26_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_24_lut_LC_6_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1704_24_lut_LC_6_26_6 (
            .in0(_gnd_net_),
            .in1(N__32591),
            .in2(N__54745),
            .in3(N__32760),
            .lcout(n2579),
            .ltout(),
            .carryin(n12760),
            .carryout(n12761),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1704_25_lut_LC_6_26_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1704_25_lut_LC_6_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1704_25_lut_LC_6_26_7.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1704_25_lut_LC_6_26_7 (
            .in0(N__54381),
            .in1(N__36113),
            .in2(N__32757),
            .in3(N__32739),
            .lcout(n2610),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1645_3_lut_LC_6_27_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1645_3_lut_LC_6_27_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1645_3_lut_LC_6_27_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1645_3_lut_LC_6_27_0 (
            .in0(_gnd_net_),
            .in1(N__32703),
            .in2(N__32673),
            .in3(N__35900),
            .lcout(n2517),
            .ltout(n2517_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1712_3_lut_LC_6_27_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1712_3_lut_LC_6_27_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1712_3_lut_LC_6_27_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1712_3_lut_LC_6_27_1 (
            .in0(_gnd_net_),
            .in1(N__32637),
            .in2(N__32631),
            .in3(N__36098),
            .lcout(n2616),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1707_3_lut_LC_6_27_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1707_3_lut_LC_6_27_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1707_3_lut_LC_6_27_3.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1707_3_lut_LC_6_27_3 (
            .in0(N__32592),
            .in1(_gnd_net_),
            .in2(N__32568),
            .in3(N__36099),
            .lcout(n2611),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12755_1_lut_LC_6_27_4.C_ON=1'b0;
    defparam i12755_1_lut_LC_6_27_4.SEQ_MODE=4'b0000;
    defparam i12755_1_lut_LC_6_27_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12755_1_lut_LC_6_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35099),
            .lcout(n15485),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2133_3_lut_LC_6_27_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2133_3_lut_LC_6_27_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2133_3_lut_LC_6_27_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2133_3_lut_LC_6_27_5 (
            .in0(_gnd_net_),
            .in1(N__32961),
            .in2(N__32943),
            .in3(N__34917),
            .lcout(n3229),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2129_3_lut_LC_6_28_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2129_3_lut_LC_6_28_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2129_3_lut_LC_6_28_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i2129_3_lut_LC_6_28_1 (
            .in0(_gnd_net_),
            .in1(N__32928),
            .in2(N__34923),
            .in3(N__32915),
            .lcout(n3225),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12562_1_lut_LC_6_28_2.C_ON=1'b0;
    defparam i12562_1_lut_LC_6_28_2.SEQ_MODE=4'b0000;
    defparam i12562_1_lut_LC_6_28_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12562_1_lut_LC_6_28_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36297),
            .lcout(n15292),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i8_1_lut_LC_6_28_3.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i8_1_lut_LC_6_28_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i8_1_lut_LC_6_28_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i8_1_lut_LC_6_28_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36135),
            .lcout(n18_adj_558),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2137_3_lut_LC_6_28_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2137_3_lut_LC_6_28_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2137_3_lut_LC_6_28_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i2137_3_lut_LC_6_28_4 (
            .in0(N__32889),
            .in1(N__34165),
            .in2(_gnd_net_),
            .in3(N__34918),
            .lcout(n3233),
            .ltout(n3233_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9966_3_lut_LC_6_28_5.C_ON=1'b0;
    defparam i9966_3_lut_LC_6_28_5.SEQ_MODE=4'b0000;
    defparam i9966_3_lut_LC_6_28_5.LUT_INIT=16'b1111101000000000;
    LogicCell40 i9966_3_lut_LC_6_28_5 (
            .in0(N__36592),
            .in1(_gnd_net_),
            .in2(N__32874),
            .in3(N__36895),
            .lcout(),
            .ltout(n11943_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_120_LC_6_28_6.C_ON=1'b0;
    defparam i1_4_lut_adj_120_LC_6_28_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_120_LC_6_28_6.LUT_INIT=16'b1000100010000000;
    LogicCell40 i1_4_lut_adj_120_LC_6_28_6 (
            .in0(N__36793),
            .in1(N__36832),
            .in2(N__32871),
            .in3(N__36865),
            .lcout(n13875),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2192_3_lut_LC_6_29_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2192_3_lut_LC_6_29_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2192_3_lut_LC_6_29_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i2192_3_lut_LC_6_29_1 (
            .in0(_gnd_net_),
            .in1(N__37032),
            .in2(N__37058),
            .in3(N__35035),
            .lcout(),
            .ltout(n29_adj_717_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_88_LC_6_29_2.C_ON=1'b0;
    defparam i1_4_lut_adj_88_LC_6_29_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_88_LC_6_29_2.LUT_INIT=16'b1111110111111000;
    LogicCell40 i1_4_lut_adj_88_LC_6_29_2 (
            .in0(N__35036),
            .in1(N__37207),
            .in2(N__33003),
            .in3(N__37185),
            .lcout(n14270),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9964_4_lut_LC_6_29_3.C_ON=1'b0;
    defparam i9964_4_lut_LC_6_29_3.SEQ_MODE=4'b0000;
    defparam i9964_4_lut_LC_6_29_3.LUT_INIT=16'b1010000010001000;
    LogicCell40 i9964_4_lut_LC_6_29_3 (
            .in0(N__32985),
            .in1(N__36540),
            .in2(N__36558),
            .in3(N__35038),
            .lcout(),
            .ltout(n11941_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10062_4_lut_LC_6_29_4.C_ON=1'b0;
    defparam i10062_4_lut_LC_6_29_4.SEQ_MODE=4'b0000;
    defparam i10062_4_lut_LC_6_29_4.LUT_INIT=16'b1111111011110100;
    LogicCell40 i10062_4_lut_LC_6_29_4 (
            .in0(N__35039),
            .in1(N__36879),
            .in2(N__32988),
            .in3(N__36899),
            .lcout(n12039),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9902_4_lut_LC_6_29_5.C_ON=1'b0;
    defparam i9902_4_lut_LC_6_29_5.SEQ_MODE=4'b0000;
    defparam i9902_4_lut_LC_6_29_5.LUT_INIT=16'b1110111011111100;
    LogicCell40 i9902_4_lut_LC_6_29_5 (
            .in0(N__36594),
            .in1(N__36618),
            .in2(N__36570),
            .in3(N__35037),
            .lcout(n11878),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12763_4_lut_LC_6_29_6.C_ON=1'b0;
    defparam i12763_4_lut_LC_6_29_6.SEQ_MODE=4'b0000;
    defparam i12763_4_lut_LC_6_29_6.LUT_INIT=16'b0000000000100111;
    LogicCell40 i12763_4_lut_LC_6_29_6 (
            .in0(N__35040),
            .in1(N__37554),
            .in2(N__37521),
            .in3(N__33060),
            .lcout(n12051),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_130_LC_6_30_0.C_ON=1'b0;
    defparam i1_4_lut_adj_130_LC_6_30_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_130_LC_6_30_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_130_LC_6_30_0 (
            .in0(N__37753),
            .in1(N__37672),
            .in2(N__37716),
            .in3(N__32979),
            .lcout(n14788),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_113_LC_6_30_1.C_ON=1'b0;
    defparam i1_4_lut_adj_113_LC_6_30_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_113_LC_6_30_1.LUT_INIT=16'b1111111110111000;
    LogicCell40 i1_4_lut_adj_113_LC_6_30_1 (
            .in0(N__37754),
            .in1(N__35076),
            .in2(N__37731),
            .in3(N__33009),
            .lcout(),
            .ltout(n14300_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_114_LC_6_30_2.C_ON=1'b0;
    defparam i1_4_lut_adj_114_LC_6_30_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_114_LC_6_30_2.LUT_INIT=16'b1111110111111000;
    LogicCell40 i1_4_lut_adj_114_LC_6_30_2 (
            .in0(N__35077),
            .in1(N__37714),
            .in2(N__32967),
            .in3(N__37689),
            .lcout(),
            .ltout(n14302_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_115_LC_6_30_3.C_ON=1'b0;
    defparam i1_4_lut_adj_115_LC_6_30_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_115_LC_6_30_3.LUT_INIT=16'b1111101011111100;
    LogicCell40 i1_4_lut_adj_115_LC_6_30_3 (
            .in0(N__37673),
            .in1(N__37653),
            .in2(N__32964),
            .in3(N__35078),
            .lcout(),
            .ltout(n14304_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_116_LC_6_30_4.C_ON=1'b0;
    defparam i1_4_lut_adj_116_LC_6_30_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_116_LC_6_30_4.LUT_INIT=16'b1111111011110100;
    LogicCell40 i1_4_lut_adj_116_LC_6_30_4 (
            .in0(N__35079),
            .in1(N__37611),
            .in2(N__33066),
            .in3(N__37641),
            .lcout(),
            .ltout(n14306_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_117_LC_6_30_5.C_ON=1'b0;
    defparam i1_4_lut_adj_117_LC_6_30_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_117_LC_6_30_5.LUT_INIT=16'b1111101011111100;
    LogicCell40 i1_4_lut_adj_117_LC_6_30_5 (
            .in0(N__37599),
            .in1(N__37566),
            .in2(N__33063),
            .in3(N__35080),
            .lcout(n14308),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i16_4_lut_LC_6_30_6.C_ON=1'b0;
    defparam i16_4_lut_LC_6_30_6.SEQ_MODE=4'b0000;
    defparam i16_4_lut_LC_6_30_6.LUT_INIT=16'b1100101000001010;
    LogicCell40 i16_4_lut_LC_6_30_6 (
            .in0(N__36813),
            .in1(N__36866),
            .in2(N__35095),
            .in3(N__36833),
            .lcout(n5_adj_704),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_103_LC_6_31_0.C_ON=1'b0;
    defparam i1_4_lut_adj_103_LC_6_31_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_103_LC_6_31_0.LUT_INIT=16'b1111111111101010;
    LogicCell40 i1_4_lut_adj_103_LC_6_31_0 (
            .in0(N__33162),
            .in1(N__33054),
            .in2(N__33048),
            .in3(N__33024),
            .lcout(),
            .ltout(n14292_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_104_LC_6_31_1.C_ON=1'b0;
    defparam i1_4_lut_adj_104_LC_6_31_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_104_LC_6_31_1.LUT_INIT=16'b1111101011111100;
    LogicCell40 i1_4_lut_adj_104_LC_6_31_1 (
            .in0(N__37307),
            .in1(N__37290),
            .in2(N__33036),
            .in3(N__35068),
            .lcout(n14294),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_98_LC_6_31_2.C_ON=1'b0;
    defparam i1_4_lut_adj_98_LC_6_31_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_98_LC_6_31_2.LUT_INIT=16'b1111111111001010;
    LogicCell40 i1_4_lut_adj_98_LC_6_31_2 (
            .in0(N__37383),
            .in1(N__37403),
            .in2(N__35093),
            .in3(N__33033),
            .lcout(),
            .ltout(n14286_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_102_LC_6_31_3.C_ON=1'b0;
    defparam i1_4_lut_adj_102_LC_6_31_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_102_LC_6_31_3.LUT_INIT=16'b1111101011111100;
    LogicCell40 i1_4_lut_adj_102_LC_6_31_3 (
            .in0(N__37374),
            .in1(N__37350),
            .in2(N__33027),
            .in3(N__35067),
            .lcout(n14288),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_109_LC_6_31_4.C_ON=1'b0;
    defparam i1_4_lut_adj_109_LC_6_31_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_109_LC_6_31_4.LUT_INIT=16'b1111111111001010;
    LogicCell40 i1_4_lut_adj_109_LC_6_31_4 (
            .in0(N__37257),
            .in1(N__37277),
            .in2(N__35094),
            .in3(N__33018),
            .lcout(),
            .ltout(n14296_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_111_LC_6_31_5.C_ON=1'b0;
    defparam i1_4_lut_adj_111_LC_6_31_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_111_LC_6_31_5.LUT_INIT=16'b1111110011111010;
    LogicCell40 i1_4_lut_adj_111_LC_6_31_5 (
            .in0(N__37224),
            .in1(N__37246),
            .in2(N__33012),
            .in3(N__35072),
            .lcout(n14298),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i2184_3_lut_LC_6_31_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i2184_3_lut_LC_6_31_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i2184_3_lut_LC_6_31_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i2184_3_lut_LC_6_31_7 (
            .in0(_gnd_net_),
            .in1(N__37341),
            .in2(N__37320),
            .in3(N__35066),
            .lcout(n45_adj_720),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.a_new_i0_LC_6_32_1 .C_ON=1'b0;
    defparam \quad_counter0.a_new_i0_LC_6_32_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_new_i0_LC_6_32_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \quad_counter0.a_new_i0_LC_6_32_1  (
            .in0(N__33156),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\quad_counter0.a_new_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56222),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1318_3_lut_LC_7_16_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1318_3_lut_LC_7_16_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1318_3_lut_LC_7_16_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1318_3_lut_LC_7_16_5 (
            .in0(_gnd_net_),
            .in1(N__37866),
            .in2(N__39354),
            .in3(N__41370),
            .lcout(n2030),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1242_3_lut_LC_7_17_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1242_3_lut_LC_7_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1242_3_lut_LC_7_17_0.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1242_3_lut_LC_7_17_0 (
            .in0(N__41007),
            .in1(_gnd_net_),
            .in2(N__43035),
            .in3(N__41515),
            .lcout(n1922),
            .ltout(n1922_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1309_3_lut_LC_7_17_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1309_3_lut_LC_7_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1309_3_lut_LC_7_17_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1309_3_lut_LC_7_17_1 (
            .in0(_gnd_net_),
            .in1(N__38016),
            .in2(N__33144),
            .in3(N__41357),
            .lcout(n2021),
            .ltout(n2021_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1376_3_lut_LC_7_17_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1376_3_lut_LC_7_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1376_3_lut_LC_7_17_2.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1376_3_lut_LC_7_17_2 (
            .in0(N__33123),
            .in1(_gnd_net_),
            .in2(N__33117),
            .in3(N__35296),
            .lcout(n2120),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1317_3_lut_LC_7_17_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1317_3_lut_LC_7_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1317_3_lut_LC_7_17_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1317_3_lut_LC_7_17_3 (
            .in0(_gnd_net_),
            .in1(N__39123),
            .in2(N__37854),
            .in3(N__41356),
            .lcout(n2029),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10008_4_lut_LC_7_17_4.C_ON=1'b0;
    defparam i10008_4_lut_LC_7_17_4.SEQ_MODE=4'b0000;
    defparam i10008_4_lut_LC_7_17_4.LUT_INIT=16'b1111111111001000;
    LogicCell40 i10008_4_lut_LC_7_17_4 (
            .in0(N__38118),
            .in1(N__39536),
            .in2(N__39321),
            .in3(N__39353),
            .lcout(n11985),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1308_3_lut_LC_7_17_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1308_3_lut_LC_7_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1308_3_lut_LC_7_17_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1308_3_lut_LC_7_17_5 (
            .in0(_gnd_net_),
            .in1(N__37911),
            .in2(N__38004),
            .in3(N__41358),
            .lcout(n2020),
            .ltout(n2020_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1375_3_lut_LC_7_17_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1375_3_lut_LC_7_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1375_3_lut_LC_7_17_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1375_3_lut_LC_7_17_6 (
            .in0(_gnd_net_),
            .in1(N__33237),
            .in2(N__33231),
            .in3(N__35297),
            .lcout(n2119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1316_3_lut_LC_7_18_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1316_3_lut_LC_7_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1316_3_lut_LC_7_18_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1316_3_lut_LC_7_18_0 (
            .in0(_gnd_net_),
            .in1(N__39285),
            .in2(N__37836),
            .in3(N__41332),
            .lcout(n2028),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12944_1_lut_LC_7_18_1.C_ON=1'b0;
    defparam i12944_1_lut_LC_7_18_1.SEQ_MODE=4'b0000;
    defparam i12944_1_lut_LC_7_18_1.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12944_1_lut_LC_7_18_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41367),
            .in3(_gnd_net_),
            .lcout(n15674),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1315_3_lut_LC_7_18_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1315_3_lut_LC_7_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1315_3_lut_LC_7_18_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1315_3_lut_LC_7_18_2 (
            .in0(_gnd_net_),
            .in1(N__39246),
            .in2(N__37818),
            .in3(N__41333),
            .lcout(n2027),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_142_LC_7_18_3.C_ON=1'b0;
    defparam i1_4_lut_adj_142_LC_7_18_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_142_LC_7_18_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_142_LC_7_18_3 (
            .in0(N__38027),
            .in1(N__37906),
            .in2(N__39555),
            .in3(N__41103),
            .lcout(),
            .ltout(n14446_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_144_LC_7_18_4.C_ON=1'b0;
    defparam i1_4_lut_adj_144_LC_7_18_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_144_LC_7_18_4.LUT_INIT=16'b1111111011111100;
    LogicCell40 i1_4_lut_adj_144_LC_7_18_4 (
            .in0(N__38169),
            .in1(N__41420),
            .in2(N__33195),
            .in3(N__33192),
            .lcout(),
            .ltout(n14450_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12947_4_lut_LC_7_18_5.C_ON=1'b0;
    defparam i12947_4_lut_LC_7_18_5.SEQ_MODE=4'b0000;
    defparam i12947_4_lut_LC_7_18_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12947_4_lut_LC_7_18_5 (
            .in0(N__38138),
            .in1(N__41636),
            .in2(N__33186),
            .in3(N__38159),
            .lcout(n1950),
            .ltout(n1950_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1305_3_lut_LC_7_18_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1305_3_lut_LC_7_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1305_3_lut_LC_7_18_6.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1305_3_lut_LC_7_18_6 (
            .in0(N__38160),
            .in1(_gnd_net_),
            .in2(N__33183),
            .in3(N__37968),
            .lcout(n2017),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1319_3_lut_LC_7_18_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1319_3_lut_LC_7_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1319_3_lut_LC_7_18_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1319_3_lut_LC_7_18_7 (
            .in0(N__37881),
            .in1(_gnd_net_),
            .in2(N__41366),
            .in3(N__39540),
            .lcout(n2031),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1314_3_lut_LC_7_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1314_3_lut_LC_7_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1314_3_lut_LC_7_19_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1314_3_lut_LC_7_19_0 (
            .in0(_gnd_net_),
            .in1(N__37800),
            .in2(N__41745),
            .in3(N__41340),
            .lcout(n2026),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1312_3_lut_LC_7_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1312_3_lut_LC_7_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1312_3_lut_LC_7_19_1.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1312_3_lut_LC_7_19_1 (
            .in0(_gnd_net_),
            .in1(N__39612),
            .in2(N__41368),
            .in3(N__37770),
            .lcout(n2024),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1313_3_lut_LC_7_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1313_3_lut_LC_7_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1313_3_lut_LC_7_19_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1313_3_lut_LC_7_19_2 (
            .in0(_gnd_net_),
            .in1(N__37785),
            .in2(N__41703),
            .in3(N__41342),
            .lcout(n2025),
            .ltout(n2025_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_145_LC_7_19_3.C_ON=1'b0;
    defparam i1_4_lut_adj_145_LC_7_19_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_145_LC_7_19_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_145_LC_7_19_3 (
            .in0(N__33436),
            .in1(N__33412),
            .in2(N__33396),
            .in3(N__33385),
            .lcout(n14544),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1321_3_lut_LC_7_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1321_3_lut_LC_7_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1321_3_lut_LC_7_19_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i1321_3_lut_LC_7_19_4 (
            .in0(N__38117),
            .in1(N__37506),
            .in2(_gnd_net_),
            .in3(N__41341),
            .lcout(n2033),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1310_3_lut_LC_7_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1310_3_lut_LC_7_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1310_3_lut_LC_7_19_5.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1310_3_lut_LC_7_19_5 (
            .in0(_gnd_net_),
            .in1(N__39582),
            .in2(N__41369),
            .in3(N__38049),
            .lcout(n2022),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1320_3_lut_LC_7_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1320_3_lut_LC_7_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1320_3_lut_LC_7_19_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1320_3_lut_LC_7_19_6 (
            .in0(_gnd_net_),
            .in1(N__39320),
            .in2(N__37491),
            .in3(N__41343),
            .lcout(n2032),
            .ltout(n2032_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10004_4_lut_LC_7_19_7.C_ON=1'b0;
    defparam i10004_4_lut_LC_7_19_7.SEQ_MODE=4'b0000;
    defparam i10004_4_lut_LC_7_19_7.LUT_INIT=16'b1111110011101100;
    LogicCell40 i10004_4_lut_LC_7_19_7 (
            .in0(N__38080),
            .in1(N__33334),
            .in2(N__33318),
            .in3(N__33721),
            .lcout(n11981),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12922_1_lut_LC_7_20_0.C_ON=1'b0;
    defparam i12922_1_lut_LC_7_20_0.SEQ_MODE=4'b0000;
    defparam i12922_1_lut_LC_7_20_0.LUT_INIT=16'b0011001100110011;
    LogicCell40 i12922_1_lut_LC_7_20_0 (
            .in0(_gnd_net_),
            .in1(N__41519),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n15652),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_146_LC_7_20_1.C_ON=1'b0;
    defparam i1_4_lut_adj_146_LC_7_20_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_146_LC_7_20_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_146_LC_7_20_1 (
            .in0(N__33307),
            .in1(N__33286),
            .in2(N__33268),
            .in3(N__33243),
            .lcout(),
            .ltout(n14550_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_147_LC_7_20_2.C_ON=1'b0;
    defparam i1_4_lut_adj_147_LC_7_20_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_147_LC_7_20_2.LUT_INIT=16'b1111100011110000;
    LogicCell40 i1_4_lut_adj_147_LC_7_20_2 (
            .in0(N__33816),
            .in1(N__33805),
            .in2(N__33780),
            .in3(N__33775),
            .lcout(n14552),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1388_3_lut_LC_7_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1388_3_lut_LC_7_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1388_3_lut_LC_7_20_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1388_3_lut_LC_7_20_4 (
            .in0(_gnd_net_),
            .in1(N__33744),
            .in2(N__33731),
            .in3(N__35243),
            .lcout(n2132),
            .ltout(n2132_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9933_3_lut_LC_7_20_5.C_ON=1'b0;
    defparam i9933_3_lut_LC_7_20_5.SEQ_MODE=4'b0000;
    defparam i9933_3_lut_LC_7_20_5.LUT_INIT=16'b1111000011000000;
    LogicCell40 i9933_3_lut_LC_7_20_5 (
            .in0(_gnd_net_),
            .in1(N__33620),
            .in2(N__33681),
            .in3(N__33661),
            .lcout(n11909),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i13_3_lut_LC_7_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i13_3_lut_LC_7_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i13_3_lut_LC_7_21_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i13_3_lut_LC_7_21_0 (
            .in0(N__38364),
            .in1(N__49591),
            .in2(_gnd_net_),
            .in3(N__39972),
            .lcout(n307),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i10_3_lut_LC_7_21_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i10_3_lut_LC_7_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i10_3_lut_LC_7_21_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i10_3_lut_LC_7_21_2 (
            .in0(N__38415),
            .in1(N__49592),
            .in2(_gnd_net_),
            .in3(N__39699),
            .lcout(n310),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i8_3_lut_LC_7_21_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i8_3_lut_LC_7_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i8_3_lut_LC_7_21_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i8_3_lut_LC_7_21_3 (
            .in0(N__49593),
            .in1(N__38469),
            .in2(_gnd_net_),
            .in3(N__39765),
            .lcout(n312),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i7_3_lut_LC_7_22_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i7_3_lut_LC_7_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i7_3_lut_LC_7_22_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i7_3_lut_LC_7_22_0 (
            .in0(N__38490),
            .in1(N__49623),
            .in2(_gnd_net_),
            .in3(N__39384),
            .lcout(n313),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i6_3_lut_LC_7_22_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i6_3_lut_LC_7_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i6_3_lut_LC_7_22_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i6_3_lut_LC_7_22_1 (
            .in0(N__49624),
            .in1(N__38511),
            .in2(_gnd_net_),
            .in3(N__39414),
            .lcout(n314),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i3_3_lut_LC_7_22_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i3_3_lut_LC_7_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i3_3_lut_LC_7_22_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i3_3_lut_LC_7_22_2 (
            .in0(N__38262),
            .in1(N__49625),
            .in2(_gnd_net_),
            .in3(N__39477),
            .lcout(n317),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i2_3_lut_LC_7_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i2_3_lut_LC_7_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i2_3_lut_LC_7_22_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i2_3_lut_LC_7_22_7 (
            .in0(N__49626),
            .in1(N__38286),
            .in2(_gnd_net_),
            .in3(N__45804),
            .lcout(n318),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_157_LC_7_23_0.C_ON=1'b0;
    defparam i1_4_lut_adj_157_LC_7_23_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_157_LC_7_23_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_157_LC_7_23_0 (
            .in0(N__33944),
            .in1(N__33997),
            .in2(N__34075),
            .in3(N__33832),
            .lcout(n14184),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i1_3_lut_LC_7_23_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i1_3_lut_LC_7_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i1_3_lut_LC_7_23_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i1_3_lut_LC_7_23_2 (
            .in0(N__49621),
            .in1(N__38301),
            .in2(_gnd_net_),
            .in3(N__39513),
            .lcout(n319),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1650_3_lut_LC_7_23_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1650_3_lut_LC_7_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1650_3_lut_LC_7_23_3.LUT_INIT=16'b1110111001000100;
    LogicCell40 encoder0_position_31__I_0_i1650_3_lut_LC_7_23_3 (
            .in0(N__35903),
            .in1(N__34125),
            .in2(_gnd_net_),
            .in3(N__34118),
            .lcout(n2522),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1649_3_lut_LC_7_23_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1649_3_lut_LC_7_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1649_3_lut_LC_7_23_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1649_3_lut_LC_7_23_4 (
            .in0(_gnd_net_),
            .in1(N__34053),
            .in2(N__34047),
            .in3(N__35902),
            .lcout(n2521),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12486_3_lut_LC_7_23_5.C_ON=1'b0;
    defparam i12486_3_lut_LC_7_23_5.SEQ_MODE=4'b0000;
    defparam i12486_3_lut_LC_7_23_5.LUT_INIT=16'b1100111111000000;
    LogicCell40 i12486_3_lut_LC_7_23_5 (
            .in0(_gnd_net_),
            .in1(N__33983),
            .in2(N__35912),
            .in3(N__33957),
            .lcout(n2525),
            .ltout(n2525_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1720_3_lut_LC_7_23_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1720_3_lut_LC_7_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1720_3_lut_LC_7_23_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1720_3_lut_LC_7_23_6 (
            .in0(_gnd_net_),
            .in1(N__33933),
            .in2(N__33924),
            .in3(N__36096),
            .lcout(n2624),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1646_3_lut_LC_7_23_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1646_3_lut_LC_7_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1646_3_lut_LC_7_23_7.LUT_INIT=16'b1110010011100100;
    LogicCell40 encoder0_position_31__I_0_i1646_3_lut_LC_7_23_7 (
            .in0(N__35904),
            .in1(N__33885),
            .in2(N__33879),
            .in3(_gnd_net_),
            .lcout(n2518),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i5_3_lut_LC_7_24_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i5_3_lut_LC_7_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i5_3_lut_LC_7_24_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i5_3_lut_LC_7_24_1 (
            .in0(N__49605),
            .in1(N__38226),
            .in2(_gnd_net_),
            .in3(N__39447),
            .lcout(n315),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i9_3_lut_LC_7_24_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i9_3_lut_LC_7_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i9_3_lut_LC_7_24_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i9_3_lut_LC_7_24_6 (
            .in0(N__38442),
            .in1(N__49604),
            .in2(_gnd_net_),
            .in3(N__39735),
            .lcout(n311),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i0_LC_7_25_0.C_ON=1'b1;
    defparam encoder0_position_scaled_i0_LC_7_25_0.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i0_LC_7_25_0.LUT_INIT=16'b1000101110111000;
    LogicCell40 encoder0_position_scaled_i0_LC_7_25_0 (
            .in0(N__36627),
            .in1(N__40111),
            .in2(N__36648),
            .in3(N__35118),
            .lcout(encoder0_position_scaled_0),
            .ltout(),
            .carryin(bfn_7_25_0_),
            .carryout(n12952),
            .clk(N__56209),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i1_LC_7_25_1.C_ON=1'b1;
    defparam encoder0_position_scaled_i1_LC_7_25_1.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i1_LC_7_25_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i1_LC_7_25_1 (
            .in0(N__35115),
            .in1(N__35103),
            .in2(N__40169),
            .in3(N__34950),
            .lcout(encoder0_position_scaled_1),
            .ltout(),
            .carryin(n12952),
            .carryout(n12953),
            .clk(N__56209),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i2_LC_7_25_2.C_ON=1'b1;
    defparam encoder0_position_scaled_i2_LC_7_25_2.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i2_LC_7_25_2.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i2_LC_7_25_2 (
            .in0(N__34947),
            .in1(N__34922),
            .in2(N__40173),
            .in3(N__34743),
            .lcout(encoder0_position_scaled_2),
            .ltout(),
            .carryin(n12953),
            .carryout(n12954),
            .clk(N__56209),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i3_LC_7_25_3.C_ON=1'b1;
    defparam encoder0_position_scaled_i3_LC_7_25_3.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i3_LC_7_25_3.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i3_LC_7_25_3 (
            .in0(N__34740),
            .in1(N__34715),
            .in2(N__40170),
            .in3(N__34542),
            .lcout(encoder0_position_scaled_3),
            .ltout(),
            .carryin(n12954),
            .carryout(n12955),
            .clk(N__56209),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i4_LC_7_25_4.C_ON=1'b1;
    defparam encoder0_position_scaled_i4_LC_7_25_4.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i4_LC_7_25_4.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i4_LC_7_25_4 (
            .in0(N__34539),
            .in1(N__34515),
            .in2(N__40174),
            .in3(N__34359),
            .lcout(encoder0_position_scaled_4),
            .ltout(),
            .carryin(n12955),
            .carryout(n12956),
            .clk(N__56209),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i5_LC_7_25_5.C_ON=1'b1;
    defparam encoder0_position_scaled_i5_LC_7_25_5.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i5_LC_7_25_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i5_LC_7_25_5 (
            .in0(N__34356),
            .in1(N__34334),
            .in2(N__40171),
            .in3(N__34173),
            .lcout(encoder0_position_scaled_5),
            .ltout(),
            .carryin(n12956),
            .carryout(n12957),
            .clk(N__56209),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i6_LC_7_25_6.C_ON=1'b1;
    defparam encoder0_position_scaled_i6_LC_7_25_6.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i6_LC_7_25_6.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i6_LC_7_25_6 (
            .in0(N__36492),
            .in1(N__36465),
            .in2(N__40175),
            .in3(N__36312),
            .lcout(encoder0_position_scaled_6),
            .ltout(),
            .carryin(n12957),
            .carryout(n12958),
            .clk(N__56209),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i7_LC_7_25_7.C_ON=1'b1;
    defparam encoder0_position_scaled_i7_LC_7_25_7.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i7_LC_7_25_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i7_LC_7_25_7 (
            .in0(N__36309),
            .in1(N__36296),
            .in2(N__40172),
            .in3(N__36123),
            .lcout(encoder0_position_scaled_7),
            .ltout(),
            .carryin(n12958),
            .carryout(n12959),
            .clk(N__56209),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i8_LC_7_26_0.C_ON=1'b1;
    defparam encoder0_position_scaled_i8_LC_7_26_0.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i8_LC_7_26_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i8_LC_7_26_0 (
            .in0(N__36120),
            .in1(N__36101),
            .in2(N__40220),
            .in3(N__35952),
            .lcout(encoder0_position_scaled_8),
            .ltout(),
            .carryin(bfn_7_26_0_),
            .carryout(n12960),
            .clk(N__56211),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i9_LC_7_26_1.C_ON=1'b1;
    defparam encoder0_position_scaled_i9_LC_7_26_1.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i9_LC_7_26_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i9_LC_7_26_1 (
            .in0(N__35949),
            .in1(N__35901),
            .in2(N__40224),
            .in3(N__35781),
            .lcout(encoder0_position_scaled_9),
            .ltout(),
            .carryin(n12960),
            .carryout(n12961),
            .clk(N__56211),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i10_LC_7_26_2.C_ON=1'b1;
    defparam encoder0_position_scaled_i10_LC_7_26_2.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i10_LC_7_26_2.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i10_LC_7_26_2 (
            .in0(N__35778),
            .in1(N__35754),
            .in2(N__40221),
            .in3(N__35628),
            .lcout(encoder0_position_scaled_10),
            .ltout(),
            .carryin(n12961),
            .carryout(n12962),
            .clk(N__56211),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i11_LC_7_26_3.C_ON=1'b1;
    defparam encoder0_position_scaled_i11_LC_7_26_3.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i11_LC_7_26_3.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i11_LC_7_26_3 (
            .in0(N__35625),
            .in1(N__35601),
            .in2(N__40225),
            .in3(N__35475),
            .lcout(encoder0_position_scaled_11),
            .ltout(),
            .carryin(n12962),
            .carryout(n12963),
            .clk(N__56211),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i12_LC_7_26_4.C_ON=1'b1;
    defparam encoder0_position_scaled_i12_LC_7_26_4.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i12_LC_7_26_4.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i12_LC_7_26_4 (
            .in0(N__35472),
            .in1(N__35451),
            .in2(N__40222),
            .in3(N__35328),
            .lcout(encoder0_position_scaled_12),
            .ltout(),
            .carryin(n12963),
            .carryout(n12964),
            .clk(N__56211),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i13_LC_7_26_5.C_ON=1'b1;
    defparam encoder0_position_scaled_i13_LC_7_26_5.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i13_LC_7_26_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i13_LC_7_26_5 (
            .in0(N__35325),
            .in1(N__35304),
            .in2(N__40226),
            .in3(N__35181),
            .lcout(encoder0_position_scaled_13),
            .ltout(),
            .carryin(n12964),
            .carryout(n12965),
            .clk(N__56211),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i14_LC_7_26_6.C_ON=1'b1;
    defparam encoder0_position_scaled_i14_LC_7_26_6.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i14_LC_7_26_6.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i14_LC_7_26_6 (
            .in0(N__37952),
            .in1(N__41382),
            .in2(N__40223),
            .in3(N__36531),
            .lcout(encoder0_position_scaled_14),
            .ltout(),
            .carryin(n12965),
            .carryout(n12966),
            .clk(N__56211),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i15_LC_7_26_7.C_ON=1'b1;
    defparam encoder0_position_scaled_i15_LC_7_26_7.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i15_LC_7_26_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i15_LC_7_26_7 (
            .in0(N__36528),
            .in1(N__41523),
            .in2(N__40227),
            .in3(N__36516),
            .lcout(encoder0_position_scaled_15),
            .ltout(),
            .carryin(n12966),
            .carryout(n12967),
            .clk(N__56211),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i16_LC_7_27_0.C_ON=1'b1;
    defparam encoder0_position_scaled_i16_LC_7_27_0.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i16_LC_7_27_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i16_LC_7_27_0 (
            .in0(N__45399),
            .in1(N__45510),
            .in2(N__40228),
            .in3(N__36513),
            .lcout(encoder0_position_scaled_16),
            .ltout(),
            .carryin(bfn_7_27_0_),
            .carryout(n12968),
            .clk(N__56214),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i17_LC_7_27_1.C_ON=1'b1;
    defparam encoder0_position_scaled_i17_LC_7_27_1.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i17_LC_7_27_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i17_LC_7_27_1 (
            .in0(N__45180),
            .in1(N__45621),
            .in2(N__40232),
            .in3(N__36510),
            .lcout(encoder0_position_scaled_17),
            .ltout(),
            .carryin(n12968),
            .carryout(n12969),
            .clk(N__56214),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i18_LC_7_27_2.C_ON=1'b1;
    defparam encoder0_position_scaled_i18_LC_7_27_2.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i18_LC_7_27_2.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i18_LC_7_27_2 (
            .in0(N__52479),
            .in1(N__48900),
            .in2(N__40229),
            .in3(N__36507),
            .lcout(encoder0_position_scaled_18),
            .ltout(),
            .carryin(n12969),
            .carryout(n12970),
            .clk(N__56214),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i19_LC_7_27_3.C_ON=1'b1;
    defparam encoder0_position_scaled_i19_LC_7_27_3.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i19_LC_7_27_3.LUT_INIT=16'b1000101110111000;
    LogicCell40 encoder0_position_scaled_i19_LC_7_27_3 (
            .in0(N__51753),
            .in1(N__40206),
            .in2(N__49014),
            .in3(N__36504),
            .lcout(encoder0_position_scaled_19),
            .ltout(),
            .carryin(n12970),
            .carryout(n12971),
            .clk(N__56214),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i20_LC_7_27_4.C_ON=1'b1;
    defparam encoder0_position_scaled_i20_LC_7_27_4.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i20_LC_7_27_4.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i20_LC_7_27_4 (
            .in0(N__47502),
            .in1(N__52359),
            .in2(N__40230),
            .in3(N__36501),
            .lcout(encoder0_position_scaled_20),
            .ltout(),
            .carryin(n12971),
            .carryout(n12972),
            .clk(N__56214),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i21_LC_7_27_5.C_ON=1'b1;
    defparam encoder0_position_scaled_i21_LC_7_27_5.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i21_LC_7_27_5.LUT_INIT=16'b1000101110111000;
    LogicCell40 encoder0_position_scaled_i21_LC_7_27_5 (
            .in0(N__52632),
            .in1(N__40210),
            .in2(N__53193),
            .in3(N__36498),
            .lcout(encoder0_position_scaled_21),
            .ltout(),
            .carryin(n12972),
            .carryout(n12973),
            .clk(N__56214),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i22_LC_7_27_6.C_ON=1'b1;
    defparam encoder0_position_scaled_i22_LC_7_27_6.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i22_LC_7_27_6.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i22_LC_7_27_6 (
            .in0(N__47745),
            .in1(N__49953),
            .in2(N__40231),
            .in3(N__36495),
            .lcout(encoder0_position_scaled_22),
            .ltout(),
            .carryin(n12973),
            .carryout(n12974),
            .clk(N__56214),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_scaled_i23_LC_7_27_7.C_ON=1'b0;
    defparam encoder0_position_scaled_i23_LC_7_27_7.SEQ_MODE=4'b1000;
    defparam encoder0_position_scaled_i23_LC_7_27_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 encoder0_position_scaled_i23_LC_7_27_7 (
            .in0(N__38673),
            .in1(N__49881),
            .in2(N__40233),
            .in3(N__36651),
            .lcout(encoder0_position_scaled_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56214),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i15_1_lut_LC_7_28_1.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i15_1_lut_LC_7_28_1.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i15_1_lut_LC_7_28_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i15_1_lut_LC_7_28_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44121),
            .lcout(n11_adj_583),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12760_1_lut_LC_7_28_2.C_ON=1'b0;
    defparam i12760_1_lut_LC_7_28_2.SEQ_MODE=4'b0000;
    defparam i12760_1_lut_LC_7_28_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12760_1_lut_LC_7_28_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36641),
            .lcout(n15490),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i10_1_lut_LC_7_28_3.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i10_1_lut_LC_7_28_3.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i10_1_lut_LC_7_28_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i10_1_lut_LC_7_28_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44270),
            .lcout(n16_adj_588),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i12_1_lut_LC_7_28_4.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i12_1_lut_LC_7_28_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i12_1_lut_LC_7_28_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i12_1_lut_LC_7_28_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44202),
            .lcout(n14_adj_586),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i9_1_lut_LC_7_28_5.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i9_1_lut_LC_7_28_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i9_1_lut_LC_7_28_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i9_1_lut_LC_7_28_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44310),
            .lcout(n17_adj_589),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_2_LC_7_29_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_2_LC_7_29_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_2_LC_7_29_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 encoder0_position_31__I_0_add_2173_2_LC_7_29_0 (
            .in0(_gnd_net_),
            .in1(N__36617),
            .in2(N__54369),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_29_0_),
            .carryout(n12921),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_3_lut_LC_7_29_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_3_lut_LC_7_29_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_3_lut_LC_7_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_3_lut_LC_7_29_1 (
            .in0(_gnd_net_),
            .in1(N__36593),
            .in2(_gnd_net_),
            .in3(N__36561),
            .lcout(n3301),
            .ltout(),
            .carryin(n12921),
            .carryout(n12922),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_4_lut_LC_7_29_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_4_lut_LC_7_29_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_4_lut_LC_7_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_4_lut_LC_7_29_2 (
            .in0(_gnd_net_),
            .in1(N__54074),
            .in2(N__36557),
            .in3(N__36534),
            .lcout(n3300),
            .ltout(),
            .carryin(n12922),
            .carryout(n12923),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_5_lut_LC_7_29_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_5_lut_LC_7_29_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_5_lut_LC_7_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_5_lut_LC_7_29_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36903),
            .in3(N__36873),
            .lcout(n3299),
            .ltout(),
            .carryin(n12923),
            .carryout(n12924),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_6_lut_LC_7_29_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_6_lut_LC_7_29_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_6_lut_LC_7_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_6_lut_LC_7_29_4 (
            .in0(_gnd_net_),
            .in1(N__54075),
            .in2(N__36870),
            .in3(N__36846),
            .lcout(n3298),
            .ltout(),
            .carryin(n12924),
            .carryout(n12925),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_7_lut_LC_7_29_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_7_lut_LC_7_29_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_7_lut_LC_7_29_5.LUT_INIT=16'b1000001000101000;
    LogicCell40 encoder0_position_31__I_0_add_2173_7_lut_LC_7_29_5 (
            .in0(N__36843),
            .in1(_gnd_net_),
            .in2(N__36837),
            .in3(N__36804),
            .lcout(n15079),
            .ltout(),
            .carryin(n12925),
            .carryout(n12926),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_8_lut_LC_7_29_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_8_lut_LC_7_29_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_8_lut_LC_7_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_8_lut_LC_7_29_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36800),
            .in3(N__36762),
            .lcout(n3296),
            .ltout(),
            .carryin(n12926),
            .carryout(n12927),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_9_lut_LC_7_29_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_9_lut_LC_7_29_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_9_lut_LC_7_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_9_lut_LC_7_29_7 (
            .in0(_gnd_net_),
            .in1(N__53982),
            .in2(N__36759),
            .in3(N__36726),
            .lcout(n3295),
            .ltout(),
            .carryin(n12927),
            .carryout(n12928),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_10_lut_LC_7_30_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_10_lut_LC_7_30_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_10_lut_LC_7_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_10_lut_LC_7_30_0 (
            .in0(_gnd_net_),
            .in1(N__53975),
            .in2(N__36723),
            .in3(N__36684),
            .lcout(n3294),
            .ltout(),
            .carryin(bfn_7_30_0_),
            .carryout(n12929),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_11_lut_LC_7_30_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_11_lut_LC_7_30_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_11_lut_LC_7_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_11_lut_LC_7_30_1 (
            .in0(_gnd_net_),
            .in1(N__54021),
            .in2(N__36681),
            .in3(N__36654),
            .lcout(n3293),
            .ltout(),
            .carryin(n12929),
            .carryout(n12930),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_12_lut_LC_7_30_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_12_lut_LC_7_30_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_12_lut_LC_7_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_12_lut_LC_7_30_2 (
            .in0(_gnd_net_),
            .in1(N__53976),
            .in2(N__37212),
            .in3(N__37179),
            .lcout(n3292),
            .ltout(),
            .carryin(n12930),
            .carryout(n12931),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_13_lut_LC_7_30_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_13_lut_LC_7_30_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_13_lut_LC_7_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_13_lut_LC_7_30_3 (
            .in0(_gnd_net_),
            .in1(N__54022),
            .in2(N__37176),
            .in3(N__37143),
            .lcout(n3291),
            .ltout(),
            .carryin(n12931),
            .carryout(n12932),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_14_lut_LC_7_30_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_14_lut_LC_7_30_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_14_lut_LC_7_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_14_lut_LC_7_30_4 (
            .in0(_gnd_net_),
            .in1(N__53977),
            .in2(N__37140),
            .in3(N__37101),
            .lcout(n3290),
            .ltout(),
            .carryin(n12932),
            .carryout(n12933),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_15_lut_LC_7_30_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_15_lut_LC_7_30_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_15_lut_LC_7_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_15_lut_LC_7_30_5 (
            .in0(_gnd_net_),
            .in1(N__54023),
            .in2(N__37098),
            .in3(N__37062),
            .lcout(n3289),
            .ltout(),
            .carryin(n12933),
            .carryout(n12934),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_16_lut_LC_7_30_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_16_lut_LC_7_30_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_16_lut_LC_7_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_16_lut_LC_7_30_6 (
            .in0(_gnd_net_),
            .in1(N__53978),
            .in2(N__37059),
            .in3(N__37026),
            .lcout(n3288),
            .ltout(),
            .carryin(n12934),
            .carryout(n12935),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_17_lut_LC_7_30_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_17_lut_LC_7_30_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_17_lut_LC_7_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_17_lut_LC_7_30_7 (
            .in0(_gnd_net_),
            .in1(N__54024),
            .in2(N__37023),
            .in3(N__36990),
            .lcout(n3287),
            .ltout(),
            .carryin(n12935),
            .carryout(n12936),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_18_lut_LC_7_31_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_18_lut_LC_7_31_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_18_lut_LC_7_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_18_lut_LC_7_31_0 (
            .in0(_gnd_net_),
            .in1(N__53968),
            .in2(N__36987),
            .in3(N__36939),
            .lcout(n3286),
            .ltout(),
            .carryin(bfn_7_31_0_),
            .carryout(n12937),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_19_lut_LC_7_31_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_19_lut_LC_7_31_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_19_lut_LC_7_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_19_lut_LC_7_31_1 (
            .in0(_gnd_net_),
            .in1(N__54010),
            .in2(N__36936),
            .in3(N__36906),
            .lcout(n3285),
            .ltout(),
            .carryin(n12937),
            .carryout(n12938),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_20_lut_LC_7_31_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_20_lut_LC_7_31_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_20_lut_LC_7_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_20_lut_LC_7_31_2 (
            .in0(_gnd_net_),
            .in1(N__37473),
            .in2(N__54414),
            .in3(N__37440),
            .lcout(n3284),
            .ltout(),
            .carryin(n12938),
            .carryout(n12939),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_21_lut_LC_7_31_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_21_lut_LC_7_31_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_21_lut_LC_7_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_21_lut_LC_7_31_3 (
            .in0(_gnd_net_),
            .in1(N__37437),
            .in2(N__54367),
            .in3(N__37407),
            .lcout(n3283),
            .ltout(),
            .carryin(n12939),
            .carryout(n12940),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_22_lut_LC_7_31_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_22_lut_LC_7_31_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_22_lut_LC_7_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_22_lut_LC_7_31_4 (
            .in0(_gnd_net_),
            .in1(N__37404),
            .in2(N__54415),
            .in3(N__37377),
            .lcout(n3282),
            .ltout(),
            .carryin(n12940),
            .carryout(n12941),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_23_lut_LC_7_31_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_23_lut_LC_7_31_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_23_lut_LC_7_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_23_lut_LC_7_31_5 (
            .in0(_gnd_net_),
            .in1(N__37373),
            .in2(N__54368),
            .in3(N__37344),
            .lcout(n3281),
            .ltout(),
            .carryin(n12941),
            .carryout(n12942),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_24_lut_LC_7_31_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_24_lut_LC_7_31_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_24_lut_LC_7_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_24_lut_LC_7_31_6 (
            .in0(_gnd_net_),
            .in1(N__37340),
            .in2(N__54416),
            .in3(N__37311),
            .lcout(n3280),
            .ltout(),
            .carryin(n12942),
            .carryout(n12943),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_25_lut_LC_7_31_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_25_lut_LC_7_31_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_25_lut_LC_7_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_25_lut_LC_7_31_7 (
            .in0(_gnd_net_),
            .in1(N__54020),
            .in2(N__37308),
            .in3(N__37284),
            .lcout(n3279),
            .ltout(),
            .carryin(n12943),
            .carryout(n12944),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_26_lut_LC_7_32_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_26_lut_LC_7_32_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_26_lut_LC_7_32_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_26_lut_LC_7_32_0 (
            .in0(_gnd_net_),
            .in1(N__37281),
            .in2(N__53646),
            .in3(N__37251),
            .lcout(n3278),
            .ltout(),
            .carryin(bfn_7_32_0_),
            .carryout(n12945),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_27_lut_LC_7_32_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_27_lut_LC_7_32_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_27_lut_LC_7_32_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_27_lut_LC_7_32_1 (
            .in0(_gnd_net_),
            .in1(N__37248),
            .in2(N__53917),
            .in3(N__37215),
            .lcout(n3277),
            .ltout(),
            .carryin(n12945),
            .carryout(n12946),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_28_lut_LC_7_32_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_28_lut_LC_7_32_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_28_lut_LC_7_32_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_28_lut_LC_7_32_2 (
            .in0(_gnd_net_),
            .in1(N__37755),
            .in2(N__53647),
            .in3(N__37719),
            .lcout(n3276),
            .ltout(),
            .carryin(n12946),
            .carryout(n12947),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_29_lut_LC_7_32_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_29_lut_LC_7_32_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_29_lut_LC_7_32_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_29_lut_LC_7_32_3 (
            .in0(_gnd_net_),
            .in1(N__37715),
            .in2(N__53918),
            .in3(N__37680),
            .lcout(n3275),
            .ltout(),
            .carryin(n12947),
            .carryout(n12948),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_30_lut_LC_7_32_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_30_lut_LC_7_32_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_30_lut_LC_7_32_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_30_lut_LC_7_32_4 (
            .in0(_gnd_net_),
            .in1(N__37677),
            .in2(N__53648),
            .in3(N__37644),
            .lcout(n3274),
            .ltout(),
            .carryin(n12948),
            .carryout(n12949),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_31_lut_LC_7_32_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_31_lut_LC_7_32_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_31_lut_LC_7_32_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_31_lut_LC_7_32_5 (
            .in0(_gnd_net_),
            .in1(N__37640),
            .in2(N__53919),
            .in3(N__37602),
            .lcout(n3273),
            .ltout(),
            .carryin(n12949),
            .carryout(n12950),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_32_lut_LC_7_32_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_2173_32_lut_LC_7_32_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_32_lut_LC_7_32_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_2173_32_lut_LC_7_32_6 (
            .in0(_gnd_net_),
            .in1(N__37594),
            .in2(N__53649),
            .in3(N__37557),
            .lcout(n3272),
            .ltout(),
            .carryin(n12950),
            .carryout(n12951),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_2173_33_lut_LC_7_32_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_2173_33_lut_LC_7_32_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_2173_33_lut_LC_7_32_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 encoder0_position_31__I_0_add_2173_33_lut_LC_7_32_7 (
            .in0(N__53659),
            .in1(N__37549),
            .in2(_gnd_net_),
            .in3(N__37524),
            .lcout(n3271),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_2_lut_LC_9_16_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_2_lut_LC_9_16_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_2_lut_LC_9_16_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_2_lut_LC_9_16_0 (
            .in0(_gnd_net_),
            .in1(N__38107),
            .in2(_gnd_net_),
            .in3(N__37494),
            .lcout(n2001),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(n12622),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_3_lut_LC_9_16_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_3_lut_LC_9_16_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_3_lut_LC_9_16_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_3_lut_LC_9_16_1 (
            .in0(_gnd_net_),
            .in1(N__55209),
            .in2(N__39313),
            .in3(N__37476),
            .lcout(n2000),
            .ltout(),
            .carryin(n12622),
            .carryout(n12623),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_4_lut_LC_9_16_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_4_lut_LC_9_16_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_4_lut_LC_9_16_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_4_lut_LC_9_16_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39535),
            .in3(N__37869),
            .lcout(n1999),
            .ltout(),
            .carryin(n12623),
            .carryout(n12624),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_5_lut_LC_9_16_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_5_lut_LC_9_16_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_5_lut_LC_9_16_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_5_lut_LC_9_16_3 (
            .in0(_gnd_net_),
            .in1(N__55210),
            .in2(N__39349),
            .in3(N__37857),
            .lcout(n1998),
            .ltout(),
            .carryin(n12624),
            .carryout(n12625),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_6_lut_LC_9_16_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_6_lut_LC_9_16_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_6_lut_LC_9_16_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_6_lut_LC_9_16_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39118),
            .in3(N__37839),
            .lcout(n1997),
            .ltout(),
            .carryin(n12625),
            .carryout(n12626),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_7_lut_LC_9_16_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_7_lut_LC_9_16_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_7_lut_LC_9_16_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_7_lut_LC_9_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39281),
            .in3(N__37821),
            .lcout(n1996),
            .ltout(),
            .carryin(n12626),
            .carryout(n12627),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_8_lut_LC_9_16_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_8_lut_LC_9_16_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_8_lut_LC_9_16_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_8_lut_LC_9_16_6 (
            .in0(_gnd_net_),
            .in1(N__55218),
            .in2(N__39242),
            .in3(N__37803),
            .lcout(n1995),
            .ltout(),
            .carryin(n12627),
            .carryout(n12628),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_9_lut_LC_9_16_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_9_lut_LC_9_16_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_9_lut_LC_9_16_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_9_lut_LC_9_16_7 (
            .in0(_gnd_net_),
            .in1(N__55211),
            .in2(N__41744),
            .in3(N__37788),
            .lcout(n1994),
            .ltout(),
            .carryin(n12628),
            .carryout(n12629),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_10_lut_LC_9_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_10_lut_LC_9_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_10_lut_LC_9_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_10_lut_LC_9_17_0 (
            .in0(_gnd_net_),
            .in1(N__55203),
            .in2(N__41702),
            .in3(N__37773),
            .lcout(n1993),
            .ltout(),
            .carryin(bfn_9_17_0_),
            .carryout(n12630),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_11_lut_LC_9_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_11_lut_LC_9_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_11_lut_LC_9_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_11_lut_LC_9_17_1 (
            .in0(_gnd_net_),
            .in1(N__55212),
            .in2(N__39608),
            .in3(N__37758),
            .lcout(n1992),
            .ltout(),
            .carryin(n12630),
            .carryout(n12631),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_12_lut_LC_9_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_12_lut_LC_9_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_12_lut_LC_9_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_12_lut_LC_9_17_2 (
            .in0(_gnd_net_),
            .in1(N__55204),
            .in2(N__41133),
            .in3(N__38052),
            .lcout(n1991),
            .ltout(),
            .carryin(n12631),
            .carryout(n12632),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_13_lut_LC_9_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_13_lut_LC_9_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_13_lut_LC_9_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_13_lut_LC_9_17_3 (
            .in0(_gnd_net_),
            .in1(N__55213),
            .in2(N__39578),
            .in3(N__38037),
            .lcout(n1990),
            .ltout(),
            .carryin(n12632),
            .carryout(n12633),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_14_lut_LC_9_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_14_lut_LC_9_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_14_lut_LC_9_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_14_lut_LC_9_17_4 (
            .in0(_gnd_net_),
            .in1(N__55205),
            .in2(N__38034),
            .in3(N__38007),
            .lcout(n1989),
            .ltout(),
            .carryin(n12633),
            .carryout(n12634),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_15_lut_LC_9_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_15_lut_LC_9_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_15_lut_LC_9_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_15_lut_LC_9_17_5 (
            .in0(_gnd_net_),
            .in1(N__55214),
            .in2(N__37907),
            .in3(N__37992),
            .lcout(n1988),
            .ltout(),
            .carryin(n12634),
            .carryout(n12635),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_16_lut_LC_9_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_16_lut_LC_9_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_16_lut_LC_9_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_16_lut_LC_9_17_6 (
            .in0(_gnd_net_),
            .in1(N__41421),
            .in2(N__55393),
            .in3(N__37989),
            .lcout(n1987),
            .ltout(),
            .carryin(n12635),
            .carryout(n12636),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_17_lut_LC_9_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_17_lut_LC_9_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_17_lut_LC_9_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_17_lut_LC_9_17_7 (
            .in0(_gnd_net_),
            .in1(N__38137),
            .in2(N__55392),
            .in3(N__37971),
            .lcout(n1986),
            .ltout(),
            .carryin(n12636),
            .carryout(n12637),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_18_lut_LC_9_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1302_18_lut_LC_9_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_18_lut_LC_9_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1302_18_lut_LC_9_18_0 (
            .in0(_gnd_net_),
            .in1(N__38158),
            .in2(N__55340),
            .in3(N__37956),
            .lcout(n1985),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(n12638),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1302_19_lut_LC_9_18_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1302_19_lut_LC_9_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1302_19_lut_LC_9_18_1.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1302_19_lut_LC_9_18_1 (
            .in0(N__41637),
            .in1(N__55151),
            .in2(N__37953),
            .in3(N__37932),
            .lcout(n2016),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1241_3_lut_LC_9_18_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1241_3_lut_LC_9_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1241_3_lut_LC_9_18_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1241_3_lut_LC_9_18_3 (
            .in0(_gnd_net_),
            .in1(N__41091),
            .in2(N__41193),
            .in3(N__41495),
            .lcout(n1921),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_143_LC_9_18_4.C_ON=1'b0;
    defparam i1_2_lut_adj_143_LC_9_18_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_143_LC_9_18_4.LUT_INIT=16'b1111000000000000;
    LogicCell40 i1_2_lut_adj_143_LC_9_18_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39122),
            .in3(N__39280),
            .lcout(n14530),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1238_3_lut_LC_9_18_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1238_3_lut_LC_9_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1238_3_lut_LC_9_18_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1238_3_lut_LC_9_18_5 (
            .in0(_gnd_net_),
            .in1(N__41229),
            .in2(N__41160),
            .in3(N__41497),
            .lcout(n1918),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1239_3_lut_LC_9_18_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1239_3_lut_LC_9_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1239_3_lut_LC_9_18_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1239_3_lut_LC_9_18_7 (
            .in0(_gnd_net_),
            .in1(N__43194),
            .in2(N__41175),
            .in3(N__41496),
            .lcout(n1919),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut_LC_9_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut_LC_9_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut_LC_9_19_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut_LC_9_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39469),
            .lcout(n31_adj_649),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut_LC_9_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut_LC_9_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut_LC_9_19_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut_LC_9_19_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39403),
            .lcout(n28_adj_646),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i15_3_lut_LC_9_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i15_3_lut_LC_9_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i15_3_lut_LC_9_19_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i15_3_lut_LC_9_19_2 (
            .in0(N__49589),
            .in1(N__38598),
            .in2(_gnd_net_),
            .in3(N__39632),
            .lcout(n305),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut_LC_9_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut_LC_9_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut_LC_9_19_3.LUT_INIT=16'b0000111100001111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut_LC_9_19_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39506),
            .in3(_gnd_net_),
            .lcout(n33_adj_651),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i14_3_lut_LC_9_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i14_3_lut_LC_9_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i14_3_lut_LC_9_19_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i14_3_lut_LC_9_19_7 (
            .in0(N__38625),
            .in1(N__49590),
            .in2(_gnd_net_),
            .in3(N__39928),
            .lcout(n306),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i16_3_lut_LC_9_20_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i16_3_lut_LC_9_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i16_3_lut_LC_9_20_0.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_mux_3_i16_3_lut_LC_9_20_0 (
            .in0(N__39827),
            .in1(_gnd_net_),
            .in2(N__49580),
            .in3(N__38574),
            .lcout(n304),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i20_3_lut_LC_9_20_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i20_3_lut_LC_9_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i20_3_lut_LC_9_20_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i20_3_lut_LC_9_20_1 (
            .in0(N__38538),
            .in1(N__49513),
            .in2(_gnd_net_),
            .in3(N__39799),
            .lcout(n300),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut_LC_9_20_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut_LC_9_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut_LC_9_20_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut_LC_9_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39631),
            .lcout(n19_adj_637),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut_LC_9_20_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut_LC_9_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut_LC_9_20_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut_LC_9_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39826),
            .lcout(n18_adj_636),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut_LC_9_20_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut_LC_9_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut_LC_9_20_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut_LC_9_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39664),
            .lcout(n23_adj_641),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut_LC_9_20_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut_LC_9_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut_LC_9_20_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut_LC_9_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39727),
            .in3(_gnd_net_),
            .lcout(n25_adj_643),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i12_3_lut_LC_9_20_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i12_3_lut_LC_9_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i12_3_lut_LC_9_20_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i12_3_lut_LC_9_20_6 (
            .in0(N__49517),
            .in1(N__38376),
            .in2(_gnd_net_),
            .in3(N__40000),
            .lcout(n308),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut_LC_9_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut_LC_9_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut_LC_9_20_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut_LC_9_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39691),
            .lcout(n24_adj_642),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut_LC_9_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut_LC_9_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut_LC_9_21_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut_LC_9_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39760),
            .lcout(n26_adj_644),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut_LC_9_21_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut_LC_9_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut_LC_9_21_1.LUT_INIT=16'b0000111100001111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut_LC_9_21_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39801),
            .in3(_gnd_net_),
            .lcout(n14_adj_632),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut_LC_9_21_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut_LC_9_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut_LC_9_21_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut_LC_9_21_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41596),
            .lcout(n30_adj_648),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut_LC_9_21_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut_LC_9_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut_LC_9_21_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut_LC_9_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39380),
            .lcout(n27_adj_645),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i11_3_lut_LC_9_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i11_3_lut_LC_9_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i11_3_lut_LC_9_21_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i11_3_lut_LC_9_21_5 (
            .in0(N__38388),
            .in1(N__49538),
            .in2(_gnd_net_),
            .in3(N__39671),
            .lcout(n309),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut_LC_9_21_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut_LC_9_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut_LC_9_21_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut_LC_9_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41949),
            .lcout(n4_adj_622),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut_LC_9_21_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut_LC_9_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut_LC_9_21_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut_LC_9_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39440),
            .lcout(n29_adj_647),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_2_lut_LC_9_22_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_2_lut_LC_9_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_2_lut_LC_9_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_2_lut_LC_9_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38313),
            .in3(N__38289),
            .lcout(n33),
            .ltout(),
            .carryin(bfn_9_22_0_),
            .carryout(n12975),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_3_lut_LC_9_22_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_3_lut_LC_9_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_3_lut_LC_9_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_3_lut_LC_9_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45771),
            .in3(N__38277),
            .lcout(n32),
            .ltout(),
            .carryin(n12975),
            .carryout(n12976),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_4_lut_LC_9_22_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_4_lut_LC_9_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_4_lut_LC_9_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_4_lut_LC_9_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38274),
            .in3(N__38250),
            .lcout(n31),
            .ltout(),
            .carryin(n12976),
            .carryout(n12977),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_5_lut_LC_9_22_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_5_lut_LC_9_22_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_5_lut_LC_9_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_5_lut_LC_9_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38247),
            .in3(N__38238),
            .lcout(n30),
            .ltout(),
            .carryin(n12977),
            .carryout(n12978),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_6_lut_LC_9_22_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_6_lut_LC_9_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_6_lut_LC_9_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_6_lut_LC_9_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38235),
            .in3(N__38214),
            .lcout(n29),
            .ltout(),
            .carryin(n12978),
            .carryout(n12979),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_7_lut_LC_9_22_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_7_lut_LC_9_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_7_lut_LC_9_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_7_lut_LC_9_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38523),
            .in3(N__38502),
            .lcout(n28),
            .ltout(),
            .carryin(n12979),
            .carryout(n12980),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_8_lut_LC_9_22_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_8_lut_LC_9_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_8_lut_LC_9_22_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_8_lut_LC_9_22_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38499),
            .in3(N__38481),
            .lcout(n27),
            .ltout(),
            .carryin(n12980),
            .carryout(n12981),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_9_lut_LC_9_22_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_9_lut_LC_9_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_9_lut_LC_9_22_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_9_lut_LC_9_22_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38478),
            .in3(N__38457),
            .lcout(n26),
            .ltout(),
            .carryin(n12981),
            .carryout(n12982),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_10_lut_LC_9_23_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_10_lut_LC_9_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_10_lut_LC_9_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_10_lut_LC_9_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38454),
            .in3(N__38430),
            .lcout(n25),
            .ltout(),
            .carryin(bfn_9_23_0_),
            .carryout(n12983),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_11_lut_LC_9_23_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_11_lut_LC_9_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_11_lut_LC_9_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_11_lut_LC_9_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38427),
            .in3(N__38403),
            .lcout(n24),
            .ltout(),
            .carryin(n12983),
            .carryout(n12984),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_12_lut_LC_9_23_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_12_lut_LC_9_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_12_lut_LC_9_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_12_lut_LC_9_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38400),
            .in3(N__38379),
            .lcout(n23),
            .ltout(),
            .carryin(n12984),
            .carryout(n12985),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_13_lut_LC_9_23_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_13_lut_LC_9_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_13_lut_LC_9_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_13_lut_LC_9_23_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39981),
            .in3(N__38367),
            .lcout(n22),
            .ltout(),
            .carryin(n12985),
            .carryout(n12986),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_14_lut_LC_9_23_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_14_lut_LC_9_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_14_lut_LC_9_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_14_lut_LC_9_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39939),
            .in3(N__38352),
            .lcout(n21),
            .ltout(),
            .carryin(n12986),
            .carryout(n12987),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_15_lut_LC_9_23_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_15_lut_LC_9_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_15_lut_LC_9_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_15_lut_LC_9_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39909),
            .in3(N__38613),
            .lcout(n20),
            .ltout(),
            .carryin(n12987),
            .carryout(n12988),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_16_lut_LC_9_23_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_16_lut_LC_9_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_16_lut_LC_9_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_16_lut_LC_9_23_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38610),
            .in3(N__38589),
            .lcout(n19),
            .ltout(),
            .carryin(n12988),
            .carryout(n12989),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_17_lut_LC_9_23_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_17_lut_LC_9_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_17_lut_LC_9_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_17_lut_LC_9_23_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38586),
            .in3(N__38562),
            .lcout(n18),
            .ltout(),
            .carryin(n12989),
            .carryout(n12990),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_18_lut_LC_9_24_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_18_lut_LC_9_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_18_lut_LC_9_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_18_lut_LC_9_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45732),
            .in3(N__38559),
            .lcout(n17),
            .ltout(),
            .carryin(bfn_9_24_0_),
            .carryout(n12991),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_19_lut_LC_9_24_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_19_lut_LC_9_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_19_lut_LC_9_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_19_lut_LC_9_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41904),
            .in3(N__38556),
            .lcout(n16),
            .ltout(),
            .carryin(n12991),
            .carryout(n12992),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_20_lut_LC_9_24_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_20_lut_LC_9_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_20_lut_LC_9_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_20_lut_LC_9_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40326),
            .in3(N__38553),
            .lcout(n15),
            .ltout(),
            .carryin(n12992),
            .carryout(n12993),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_21_lut_LC_9_24_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_21_lut_LC_9_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_21_lut_LC_9_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_21_lut_LC_9_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38550),
            .in3(N__38529),
            .lcout(n14),
            .ltout(),
            .carryin(n12993),
            .carryout(n12994),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_22_lut_LC_9_24_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_22_lut_LC_9_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_22_lut_LC_9_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_22_lut_LC_9_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39864),
            .in3(N__38526),
            .lcout(n13),
            .ltout(),
            .carryin(n12994),
            .carryout(n12995),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_23_lut_LC_9_24_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_23_lut_LC_9_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_23_lut_LC_9_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_23_lut_LC_9_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__52389),
            .in3(N__38664),
            .lcout(n12),
            .ltout(),
            .carryin(n12995),
            .carryout(n12996),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_24_lut_LC_9_24_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_24_lut_LC_9_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_24_lut_LC_9_24_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_24_lut_LC_9_24_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45645),
            .in3(N__38661),
            .lcout(n11),
            .ltout(),
            .carryin(n12996),
            .carryout(n12997),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_25_lut_LC_9_24_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_25_lut_LC_9_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_25_lut_LC_9_24_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_25_lut_LC_9_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43719),
            .in3(N__38658),
            .lcout(n10),
            .ltout(),
            .carryin(n12997),
            .carryout(n12998),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_26_lut_LC_9_25_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_26_lut_LC_9_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_26_lut_LC_9_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_26_lut_LC_9_25_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40065),
            .in3(N__38655),
            .lcout(n9),
            .ltout(),
            .carryin(bfn_9_25_0_),
            .carryout(n12999),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_27_lut_LC_9_25_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_27_lut_LC_9_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_27_lut_LC_9_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_27_lut_LC_9_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40251),
            .in3(N__38652),
            .lcout(n8),
            .ltout(),
            .carryin(n12999),
            .carryout(n13000),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_28_lut_LC_9_25_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_28_lut_LC_9_25_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_28_lut_LC_9_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_28_lut_LC_9_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41889),
            .in3(N__38649),
            .lcout(n7),
            .ltout(),
            .carryin(n13000),
            .carryout(n13001),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_29_lut_LC_9_25_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_29_lut_LC_9_25_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_29_lut_LC_9_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_29_lut_LC_9_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40317),
            .in3(N__38646),
            .lcout(n6),
            .ltout(),
            .carryin(n13001),
            .carryout(n13002),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_30_lut_LC_9_25_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_30_lut_LC_9_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_30_lut_LC_9_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_30_lut_LC_9_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40242),
            .in3(N__38643),
            .lcout(n5),
            .ltout(),
            .carryin(n13002),
            .carryout(n13003),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_31_lut_LC_9_25_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_31_lut_LC_9_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_31_lut_LC_9_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_31_lut_LC_9_25_5 (
            .in0(_gnd_net_),
            .in1(N__38640),
            .in2(_gnd_net_),
            .in3(N__38628),
            .lcout(n4),
            .ltout(),
            .carryin(n13003),
            .carryout(n13004),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_32_lut_LC_9_25_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_32_lut_LC_9_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_32_lut_LC_9_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_32_lut_LC_9_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41874),
            .in3(N__38733),
            .lcout(n3),
            .ltout(),
            .carryin(n13004),
            .carryout(n13005),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_33_lut_LC_9_25_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_33_lut_LC_9_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_33_lut_LC_9_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_add_3_33_lut_LC_9_25_7 (
            .in0(_gnd_net_),
            .in1(N__40083),
            .in2(_gnd_net_),
            .in3(N__38730),
            .lcout(n2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i9_1_lut_LC_9_26_0.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i9_1_lut_LC_9_26_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i9_1_lut_LC_9_26_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i9_1_lut_LC_9_26_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38727),
            .lcout(n17_adj_559),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i11_1_lut_LC_9_26_1.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i11_1_lut_LC_9_26_1.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i11_1_lut_LC_9_26_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i11_1_lut_LC_9_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44231),
            .lcout(n15_adj_587),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i15_1_lut_LC_9_26_2.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i15_1_lut_LC_9_26_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i15_1_lut_LC_9_26_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i15_1_lut_LC_9_26_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38718),
            .lcout(n11_adj_565),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i11_1_lut_LC_9_26_3.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i11_1_lut_LC_9_26_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i11_1_lut_LC_9_26_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i11_1_lut_LC_9_26_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38709),
            .lcout(n15_adj_561),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i13_1_lut_LC_9_26_4.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i13_1_lut_LC_9_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i13_1_lut_LC_9_26_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i13_1_lut_LC_9_26_4 (
            .in0(N__38700),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n13_adj_563),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i14_1_lut_LC_9_26_6.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i14_1_lut_LC_9_26_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i14_1_lut_LC_9_26_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i14_1_lut_LC_9_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38691),
            .lcout(n12_adj_564),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i16_1_lut_LC_9_26_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i16_1_lut_LC_9_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i16_1_lut_LC_9_26_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i16_1_lut_LC_9_26_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38682),
            .lcout(n10_adj_566),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12778_1_lut_LC_9_27_1.C_ON=1'b0;
    defparam i12778_1_lut_LC_9_27_1.SEQ_MODE=4'b0000;
    defparam i12778_1_lut_LC_9_27_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12778_1_lut_LC_9_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49877),
            .lcout(n15508),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i19_1_lut_LC_9_27_2.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i19_1_lut_LC_9_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i19_1_lut_LC_9_27_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i19_1_lut_LC_9_27_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38763),
            .lcout(n7_adj_569),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9552_2_lut_LC_9_27_3.C_ON=1'b0;
    defparam i9552_2_lut_LC_9_27_3.SEQ_MODE=4'b0000;
    defparam i9552_2_lut_LC_9_27_3.LUT_INIT=16'b1010101000000000;
    LogicCell40 i9552_2_lut_LC_9_27_3 (
            .in0(N__46659),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46615),
            .lcout(n11526),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9553_1_lut_2_lut_LC_9_27_4.C_ON=1'b0;
    defparam i9553_1_lut_2_lut_LC_9_27_4.SEQ_MODE=4'b0000;
    defparam i9553_1_lut_2_lut_LC_9_27_4.LUT_INIT=16'b0011001111111111;
    LogicCell40 i9553_1_lut_2_lut_LC_9_27_4 (
            .in0(_gnd_net_),
            .in1(N__46614),
            .in2(_gnd_net_),
            .in3(N__46658),
            .lcout(n1377),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i24_1_lut_LC_9_27_5.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i24_1_lut_LC_9_27_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i24_1_lut_LC_9_27_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i24_1_lut_LC_9_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38754),
            .lcout(n2_adj_574),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i18_1_lut_LC_9_27_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i18_1_lut_LC_9_27_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i18_1_lut_LC_9_27_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i18_1_lut_LC_9_27_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38745),
            .lcout(n8_adj_568),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i17_1_lut_LC_9_28_0.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i17_1_lut_LC_9_28_0.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i17_1_lut_LC_9_28_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i17_1_lut_LC_9_28_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44450),
            .lcout(n9_adj_581),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12768_2_lut_LC_9_28_1.C_ON=1'b0;
    defparam i12768_2_lut_LC_9_28_1.SEQ_MODE=4'b0000;
    defparam i12768_2_lut_LC_9_28_1.LUT_INIT=16'b1111111100110011;
    LogicCell40 i12768_2_lut_LC_9_28_1 (
            .in0(_gnd_net_),
            .in1(N__46616),
            .in2(_gnd_net_),
            .in3(N__46660),
            .lcout(),
            .ltout(dti_N_333_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_LC_9_28_2.C_ON=1'b0;
    defparam i1_2_lut_4_lut_LC_9_28_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_LC_9_28_2.LUT_INIT=16'b1101111111101111;
    LogicCell40 i1_2_lut_4_lut_LC_9_28_2 (
            .in0(N__39188),
            .in1(N__46692),
            .in2(N__38736),
            .in3(N__56517),
            .lcout(n5187),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12403_2_lut_4_lut_LC_9_28_3.C_ON=1'b0;
    defparam i12403_2_lut_4_lut_LC_9_28_3.SEQ_MODE=4'b0000;
    defparam i12403_2_lut_4_lut_LC_9_28_3.LUT_INIT=16'b0100000000010000;
    LogicCell40 i12403_2_lut_4_lut_LC_9_28_3 (
            .in0(N__46693),
            .in1(N__56518),
            .in2(N__39077),
            .in3(N__39189),
            .lcout(n15072),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \debounce.reg_out_i0_i1_LC_9_28_5 .C_ON=1'b0;
    defparam \debounce.reg_out_i0_i1_LC_9_28_5 .SEQ_MODE=4'b1000;
    defparam \debounce.reg_out_i0_i1_LC_9_28_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \debounce.reg_out_i0_i1_LC_9_28_5  (
            .in0(N__46988),
            .in1(N__38895),
            .in2(_gnd_net_),
            .in3(N__38874),
            .lcout(h2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56219),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_662__i0_LC_9_29_0.C_ON=1'b1;
    defparam dti_counter_662__i0_LC_9_29_0.SEQ_MODE=4'b1000;
    defparam dti_counter_662__i0_LC_9_29_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 dti_counter_662__i0_LC_9_29_0 (
            .in0(N__38985),
            .in1(N__39002),
            .in2(N__38841),
            .in3(N__38829),
            .lcout(dti_counter_0),
            .ltout(),
            .carryin(bfn_9_29_0_),
            .carryout(n13006),
            .clk(N__56223),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_662__i1_LC_9_29_1.C_ON=1'b1;
    defparam dti_counter_662__i1_LC_9_29_1.SEQ_MODE=4'b1000;
    defparam dti_counter_662__i1_LC_9_29_1.LUT_INIT=16'b1110001000101110;
    LogicCell40 dti_counter_662__i1_LC_9_29_1 (
            .in0(N__39198),
            .in1(N__38787),
            .in2(N__39224),
            .in3(N__38826),
            .lcout(dti_counter_1),
            .ltout(),
            .carryin(n13006),
            .carryout(n13007),
            .clk(N__56223),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_662__i2_LC_9_29_2.C_ON=1'b1;
    defparam dti_counter_662__i2_LC_9_29_2.SEQ_MODE=4'b1000;
    defparam dti_counter_662__i2_LC_9_29_2.LUT_INIT=16'b1100101000111010;
    LogicCell40 dti_counter_662__i2_LC_9_29_2 (
            .in0(N__39090),
            .in1(N__39027),
            .in2(N__38800),
            .in3(N__38823),
            .lcout(dti_counter_2),
            .ltout(),
            .carryin(n13007),
            .carryout(n13008),
            .clk(N__56223),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_662__i3_LC_9_29_3.C_ON=1'b1;
    defparam dti_counter_662__i3_LC_9_29_3.SEQ_MODE=4'b1000;
    defparam dti_counter_662__i3_LC_9_29_3.LUT_INIT=16'b1110001000101110;
    LogicCell40 dti_counter_662__i3_LC_9_29_3 (
            .in0(N__38961),
            .in1(N__38791),
            .in2(N__38979),
            .in3(N__38820),
            .lcout(dti_counter_3),
            .ltout(),
            .carryin(n13008),
            .carryout(n13009),
            .clk(N__56223),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_662__i4_LC_9_29_4.C_ON=1'b1;
    defparam dti_counter_662__i4_LC_9_29_4.SEQ_MODE=4'b1000;
    defparam dti_counter_662__i4_LC_9_29_4.LUT_INIT=16'b1100101000111010;
    LogicCell40 dti_counter_662__i4_LC_9_29_4 (
            .in0(N__38937),
            .in1(N__38954),
            .in2(N__38801),
            .in3(N__38817),
            .lcout(dti_counter_4),
            .ltout(),
            .carryin(n13009),
            .carryout(n13010),
            .clk(N__56223),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_662__i5_LC_9_29_5.C_ON=1'b1;
    defparam dti_counter_662__i5_LC_9_29_5.SEQ_MODE=4'b1000;
    defparam dti_counter_662__i5_LC_9_29_5.LUT_INIT=16'b1110001000101110;
    LogicCell40 dti_counter_662__i5_LC_9_29_5 (
            .in0(N__38814),
            .in1(N__38795),
            .in2(N__39078),
            .in3(N__38808),
            .lcout(dti_counter_5),
            .ltout(),
            .carryin(n13010),
            .carryout(n13011),
            .clk(N__56223),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_662__i6_LC_9_29_6.C_ON=1'b1;
    defparam dti_counter_662__i6_LC_9_29_6.SEQ_MODE=4'b1000;
    defparam dti_counter_662__i6_LC_9_29_6.LUT_INIT=16'b1100101000111010;
    LogicCell40 dti_counter_662__i6_LC_9_29_6 (
            .in0(N__39084),
            .in1(N__39052),
            .in2(N__38802),
            .in3(N__38805),
            .lcout(dti_counter_6),
            .ltout(),
            .carryin(n13011),
            .carryout(n13012),
            .clk(N__56223),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_counter_662__i7_LC_9_29_7.C_ON=1'b0;
    defparam dti_counter_662__i7_LC_9_29_7.SEQ_MODE=4'b1000;
    defparam dti_counter_662__i7_LC_9_29_7.LUT_INIT=16'b1011100001110100;
    LogicCell40 dti_counter_662__i7_LC_9_29_7 (
            .in0(N__38927),
            .in1(N__38799),
            .in2(N__38907),
            .in3(N__38766),
            .lcout(dti_counter_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56223),
            .ce(),
            .sr(_gnd_net_));
    defparam i12406_2_lut_4_lut_LC_9_30_0.C_ON=1'b0;
    defparam i12406_2_lut_4_lut_LC_9_30_0.SEQ_MODE=4'b0000;
    defparam i12406_2_lut_4_lut_LC_9_30_0.LUT_INIT=16'b0000100100000000;
    LogicCell40 i12406_2_lut_4_lut_LC_9_30_0 (
            .in0(N__39184),
            .in1(N__56522),
            .in2(N__46722),
            .in3(N__39026),
            .lcout(n15075),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12390_2_lut_4_lut_LC_9_30_1.C_ON=1'b0;
    defparam i12390_2_lut_4_lut_LC_9_30_1.SEQ_MODE=4'b0000;
    defparam i12390_2_lut_4_lut_LC_9_30_1.LUT_INIT=16'b0000000010010000;
    LogicCell40 i12390_2_lut_4_lut_LC_9_30_1 (
            .in0(N__56519),
            .in1(N__39185),
            .in2(N__39054),
            .in3(N__46718),
            .lcout(n15071),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_79_LC_9_30_2.C_ON=1'b0;
    defparam i6_4_lut_adj_79_LC_9_30_2.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_79_LC_9_30_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_adj_79_LC_9_30_2 (
            .in0(N__39070),
            .in1(N__38950),
            .in2(N__39053),
            .in3(N__38923),
            .lcout(),
            .ltout(n14_adj_705_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_LC_9_30_3.C_ON=1'b0;
    defparam i7_4_lut_LC_9_30_3.SEQ_MODE=4'b0000;
    defparam i7_4_lut_LC_9_30_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i7_4_lut_LC_9_30_3 (
            .in0(N__38974),
            .in1(N__39001),
            .in2(N__39030),
            .in3(N__39012),
            .lcout(n5137),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_adj_78_LC_9_30_4.C_ON=1'b0;
    defparam i2_2_lut_adj_78_LC_9_30_4.SEQ_MODE=4'b0000;
    defparam i2_2_lut_adj_78_LC_9_30_4.LUT_INIT=16'b1111111111001100;
    LogicCell40 i2_2_lut_adj_78_LC_9_30_4 (
            .in0(_gnd_net_),
            .in1(N__39214),
            .in2(_gnd_net_),
            .in3(N__39025),
            .lcout(n10_adj_706),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12360_2_lut_4_lut_LC_9_30_5.C_ON=1'b0;
    defparam i12360_2_lut_4_lut_LC_9_30_5.SEQ_MODE=4'b0000;
    defparam i12360_2_lut_4_lut_LC_9_30_5.LUT_INIT=16'b0000000010010000;
    LogicCell40 i12360_2_lut_4_lut_LC_9_30_5 (
            .in0(N__56523),
            .in1(N__39187),
            .in2(N__39006),
            .in3(N__46720),
            .lcout(n15081),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12405_2_lut_4_lut_LC_9_30_6.C_ON=1'b0;
    defparam i12405_2_lut_4_lut_LC_9_30_6.SEQ_MODE=4'b0000;
    defparam i12405_2_lut_4_lut_LC_9_30_6.LUT_INIT=16'b0000100100000000;
    LogicCell40 i12405_2_lut_4_lut_LC_9_30_6 (
            .in0(N__39183),
            .in1(N__56521),
            .in2(N__46721),
            .in3(N__38975),
            .lcout(n15074),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12404_2_lut_4_lut_LC_9_30_7.C_ON=1'b0;
    defparam i12404_2_lut_4_lut_LC_9_30_7.SEQ_MODE=4'b0000;
    defparam i12404_2_lut_4_lut_LC_9_30_7.LUT_INIT=16'b0000000010010000;
    LogicCell40 i12404_2_lut_4_lut_LC_9_30_7 (
            .in0(N__56520),
            .in1(N__39186),
            .in2(N__38955),
            .in3(N__46719),
            .lcout(n15073),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12418_2_lut_4_lut_LC_9_31_0.C_ON=1'b0;
    defparam i12418_2_lut_4_lut_LC_9_31_0.SEQ_MODE=4'b0000;
    defparam i12418_2_lut_4_lut_LC_9_31_0.LUT_INIT=16'b0010000000010000;
    LogicCell40 i12418_2_lut_4_lut_LC_9_31_0 (
            .in0(N__56509),
            .in1(N__46711),
            .in2(N__38931),
            .in3(N__39182),
            .lcout(n15070),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_3_lut_LC_9_31_1.C_ON=1'b0;
    defparam i14_3_lut_LC_9_31_1.SEQ_MODE=4'b0000;
    defparam i14_3_lut_LC_9_31_1.LUT_INIT=16'b0111011111101110;
    LogicCell40 i14_3_lut_LC_9_31_1 (
            .in0(N__47000),
            .in1(N__46955),
            .in2(_gnd_net_),
            .in3(N__46892),
            .lcout(n6_adj_721),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12199_4_lut_LC_9_31_2.C_ON=1'b0;
    defparam i12199_4_lut_LC_9_31_2.SEQ_MODE=4'b0000;
    defparam i12199_4_lut_LC_9_31_2.LUT_INIT=16'b1111110011011000;
    LogicCell40 i12199_4_lut_LC_9_31_2 (
            .in0(N__40764),
            .in1(N__40784),
            .in2(N__40746),
            .in3(N__40992),
            .lcout(n14929),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12198_4_lut_LC_9_31_3.C_ON=1'b0;
    defparam i12198_4_lut_LC_9_31_3.SEQ_MODE=4'b0000;
    defparam i12198_4_lut_LC_9_31_3.LUT_INIT=16'b1101010011010000;
    LogicCell40 i12198_4_lut_LC_9_31_3 (
            .in0(N__40991),
            .in1(N__40763),
            .in2(N__40785),
            .in3(N__40742),
            .lcout(n14928),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12407_2_lut_4_lut_LC_9_31_4.C_ON=1'b0;
    defparam i12407_2_lut_4_lut_LC_9_31_4.SEQ_MODE=4'b0000;
    defparam i12407_2_lut_4_lut_LC_9_31_4.LUT_INIT=16'b0010000000010000;
    LogicCell40 i12407_2_lut_4_lut_LC_9_31_4 (
            .in0(N__56508),
            .in1(N__46710),
            .in2(N__39225),
            .in3(N__39181),
            .lcout(n15076),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam commutation_state_prev_i0_LC_9_31_7.C_ON=1'b0;
    defparam commutation_state_prev_i0_LC_9_31_7.SEQ_MODE=4'b1000;
    defparam commutation_state_prev_i0_LC_9_31_7.LUT_INIT=16'b1100110011001100;
    LogicCell40 commutation_state_prev_i0_LC_9_31_7 (
            .in0(_gnd_net_),
            .in1(N__56510),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(commutation_state_prev_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56235),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i18_LC_9_32_4.C_ON=1'b0;
    defparam pwm_setpoint_i18_LC_9_32_4.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i18_LC_9_32_4.LUT_INIT=16'b1110111001000100;
    LogicCell40 pwm_setpoint_i18_LC_9_32_4 (
            .in0(N__50899),
            .in1(N__44553),
            .in2(_gnd_net_),
            .in3(N__42669),
            .lcout(pwm_setpoint_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56241),
            .ce(),
            .sr(_gnd_net_));
    defparam i12200_3_lut_LC_9_32_6.C_ON=1'b0;
    defparam i12200_3_lut_LC_9_32_6.SEQ_MODE=4'b0000;
    defparam i12200_3_lut_LC_9_32_6.LUT_INIT=16'b0010001001110111;
    LogicCell40 i12200_3_lut_LC_9_32_6 (
            .in0(N__40971),
            .in1(N__39150),
            .in2(_gnd_net_),
            .in3(N__39144),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1183_3_lut_LC_10_16_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1183_3_lut_LC_10_16_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1183_3_lut_LC_10_16_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1183_3_lut_LC_10_16_0 (
            .in0(_gnd_net_),
            .in1(N__43287),
            .in2(N__43317),
            .in3(N__45500),
            .lcout(n1831),
            .ltout(n1831_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1250_3_lut_LC_10_16_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1250_3_lut_LC_10_16_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1250_3_lut_LC_10_16_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1250_3_lut_LC_10_16_1 (
            .in0(_gnd_net_),
            .in1(N__40836),
            .in2(N__39126),
            .in3(N__41490),
            .lcout(n1930),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1251_3_lut_LC_10_16_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1251_3_lut_LC_10_16_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1251_3_lut_LC_10_16_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1251_3_lut_LC_10_16_5 (
            .in0(_gnd_net_),
            .in1(N__40883),
            .in2(N__40863),
            .in3(N__41494),
            .lcout(n1931),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1253_3_lut_LC_10_16_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1253_3_lut_LC_10_16_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1253_3_lut_LC_10_16_6.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1253_3_lut_LC_10_16_6 (
            .in0(_gnd_net_),
            .in1(N__40950),
            .in2(N__41514),
            .in3(N__40920),
            .lcout(n1933),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1249_3_lut_LC_10_16_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1249_3_lut_LC_10_16_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1249_3_lut_LC_10_16_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1249_3_lut_LC_10_16_7 (
            .in0(_gnd_net_),
            .in1(N__41055),
            .in2(N__43119),
            .in3(N__41489),
            .lcout(n1929),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1243_3_lut_LC_10_17_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1243_3_lut_LC_10_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1243_3_lut_LC_10_17_0.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i1243_3_lut_LC_10_17_0 (
            .in0(N__43057),
            .in1(_gnd_net_),
            .in2(N__41019),
            .in3(N__41482),
            .lcout(n1923),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1245_3_lut_LC_10_17_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1245_3_lut_LC_10_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1245_3_lut_LC_10_17_1.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1245_3_lut_LC_10_17_1 (
            .in0(_gnd_net_),
            .in1(N__43083),
            .in2(N__41512),
            .in3(N__41031),
            .lcout(n1925),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_137_LC_10_17_2.C_ON=1'b0;
    defparam i1_3_lut_adj_137_LC_10_17_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_137_LC_10_17_2.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_137_LC_10_17_2 (
            .in0(_gnd_net_),
            .in1(N__43027),
            .in2(N__43059),
            .in3(N__42858),
            .lcout(),
            .ltout(n14524_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_138_LC_10_17_3.C_ON=1'b0;
    defparam i1_4_lut_adj_138_LC_10_17_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_138_LC_10_17_3.LUT_INIT=16'b1111100011110000;
    LogicCell40 i1_4_lut_adj_138_LC_10_17_3 (
            .in0(N__41665),
            .in1(N__43112),
            .in2(N__39255),
            .in3(N__40956),
            .lcout(),
            .ltout(n14526_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12925_4_lut_LC_10_17_4.C_ON=1'b0;
    defparam i12925_4_lut_LC_10_17_4.SEQ_MODE=4'b0000;
    defparam i12925_4_lut_LC_10_17_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12925_4_lut_LC_10_17_4 (
            .in0(N__41227),
            .in1(N__41067),
            .in2(N__39252),
            .in3(N__43748),
            .lcout(n1851),
            .ltout(n1851_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1248_3_lut_LC_10_17_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1248_3_lut_LC_10_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1248_3_lut_LC_10_17_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1248_3_lut_LC_10_17_5 (
            .in0(N__41666),
            .in1(_gnd_net_),
            .in2(N__39249),
            .in3(N__41046),
            .lcout(n1928),
            .ltout(n1928_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_141_LC_10_17_6.C_ON=1'b0;
    defparam i1_3_lut_adj_141_LC_10_17_6.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_141_LC_10_17_6.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_141_LC_10_17_6 (
            .in0(_gnd_net_),
            .in1(N__39601),
            .in2(N__39585),
            .in3(N__39571),
            .lcout(n14440),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1252_3_lut_LC_10_17_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1252_3_lut_LC_10_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1252_3_lut_LC_10_17_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1252_3_lut_LC_10_17_7 (
            .in0(_gnd_net_),
            .in1(N__40893),
            .in2(N__41513),
            .in3(N__40911),
            .lcout(n1932),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i0_LC_10_18_0 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i0_LC_10_18_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i0_LC_10_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i0_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(N__39505),
            .in2(_gnd_net_),
            .in3(N__39483),
            .lcout(encoder0_position_0),
            .ltout(),
            .carryin(bfn_10_18_0_),
            .carryout(\quad_counter0.n13095 ),
            .clk(N__56201),
            .ce(N__40308),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i1_LC_10_18_1 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i1_LC_10_18_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i1_LC_10_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i1_LC_10_18_1  (
            .in0(_gnd_net_),
            .in1(N__40455),
            .in2(N__45799),
            .in3(N__39480),
            .lcout(encoder0_position_1),
            .ltout(),
            .carryin(\quad_counter0.n13095 ),
            .carryout(\quad_counter0.n13096 ),
            .clk(N__56201),
            .ce(N__40308),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i2_LC_10_18_2 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i2_LC_10_18_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i2_LC_10_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i2_LC_10_18_2  (
            .in0(_gnd_net_),
            .in1(N__39473),
            .in2(N__40514),
            .in3(N__39453),
            .lcout(encoder0_position_2),
            .ltout(),
            .carryin(\quad_counter0.n13096 ),
            .carryout(\quad_counter0.n13097 ),
            .clk(N__56201),
            .ce(N__40308),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i3_LC_10_18_3 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i3_LC_10_18_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i3_LC_10_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i3_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(N__40459),
            .in2(N__41600),
            .in3(N__39450),
            .lcout(encoder0_position_3),
            .ltout(),
            .carryin(\quad_counter0.n13097 ),
            .carryout(\quad_counter0.n13098 ),
            .clk(N__56201),
            .ce(N__40308),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i4_LC_10_18_4 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i4_LC_10_18_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i4_LC_10_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i4_LC_10_18_4  (
            .in0(_gnd_net_),
            .in1(N__39439),
            .in2(N__40515),
            .in3(N__39417),
            .lcout(encoder0_position_4),
            .ltout(),
            .carryin(\quad_counter0.n13098 ),
            .carryout(\quad_counter0.n13099 ),
            .clk(N__56201),
            .ce(N__40308),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i5_LC_10_18_5 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i5_LC_10_18_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i5_LC_10_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i5_LC_10_18_5  (
            .in0(_gnd_net_),
            .in1(N__40463),
            .in2(N__39413),
            .in3(N__39387),
            .lcout(encoder0_position_5),
            .ltout(),
            .carryin(\quad_counter0.n13099 ),
            .carryout(\quad_counter0.n13100 ),
            .clk(N__56201),
            .ce(N__40308),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i6_LC_10_18_6 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i6_LC_10_18_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i6_LC_10_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i6_LC_10_18_6  (
            .in0(_gnd_net_),
            .in1(N__39379),
            .in2(N__40516),
            .in3(N__39357),
            .lcout(encoder0_position_6),
            .ltout(),
            .carryin(\quad_counter0.n13100 ),
            .carryout(\quad_counter0.n13101 ),
            .clk(N__56201),
            .ce(N__40308),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i7_LC_10_18_7 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i7_LC_10_18_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i7_LC_10_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i7_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(N__40467),
            .in2(N__39764),
            .in3(N__39738),
            .lcout(encoder0_position_7),
            .ltout(),
            .carryin(\quad_counter0.n13101 ),
            .carryout(\quad_counter0.n13102 ),
            .clk(N__56201),
            .ce(N__40308),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i8_LC_10_19_0 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i8_LC_10_19_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i8_LC_10_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i8_LC_10_19_0  (
            .in0(_gnd_net_),
            .in1(N__40468),
            .in2(N__39731),
            .in3(N__39702),
            .lcout(encoder0_position_8),
            .ltout(),
            .carryin(bfn_10_19_0_),
            .carryout(\quad_counter0.n13103 ),
            .clk(N__56202),
            .ce(N__40303),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i9_LC_10_19_1 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i9_LC_10_19_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i9_LC_10_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i9_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(N__39695),
            .in2(N__40517),
            .in3(N__39675),
            .lcout(encoder0_position_9),
            .ltout(),
            .carryin(\quad_counter0.n13103 ),
            .carryout(\quad_counter0.n13104 ),
            .clk(N__56202),
            .ce(N__40303),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i10_LC_10_19_2 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i10_LC_10_19_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i10_LC_10_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i10_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(N__40472),
            .in2(N__39672),
            .in3(N__39648),
            .lcout(encoder0_position_10),
            .ltout(),
            .carryin(\quad_counter0.n13104 ),
            .carryout(\quad_counter0.n13105 ),
            .clk(N__56202),
            .ce(N__40303),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i11_LC_10_19_3 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i11_LC_10_19_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i11_LC_10_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i11_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(N__40001),
            .in2(N__40518),
            .in3(N__39645),
            .lcout(encoder0_position_11),
            .ltout(),
            .carryin(\quad_counter0.n13105 ),
            .carryout(\quad_counter0.n13106 ),
            .clk(N__56202),
            .ce(N__40303),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i12_LC_10_19_4 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i12_LC_10_19_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i12_LC_10_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i12_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(N__40476),
            .in2(N__39970),
            .in3(N__39642),
            .lcout(encoder0_position_12),
            .ltout(),
            .carryin(\quad_counter0.n13106 ),
            .carryout(\quad_counter0.n13107 ),
            .clk(N__56202),
            .ce(N__40303),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i13_LC_10_19_5 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i13_LC_10_19_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i13_LC_10_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i13_LC_10_19_5  (
            .in0(_gnd_net_),
            .in1(N__39929),
            .in2(N__40519),
            .in3(N__39639),
            .lcout(encoder0_position_13),
            .ltout(),
            .carryin(\quad_counter0.n13107 ),
            .carryout(\quad_counter0.n13108 ),
            .clk(N__56202),
            .ce(N__40303),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i14_LC_10_19_6 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i14_LC_10_19_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i14_LC_10_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i14_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(N__40480),
            .in2(N__39636),
            .in3(N__39615),
            .lcout(encoder0_position_14),
            .ltout(),
            .carryin(\quad_counter0.n13108 ),
            .carryout(\quad_counter0.n13109 ),
            .clk(N__56202),
            .ce(N__40303),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i15_LC_10_19_7 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i15_LC_10_19_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i15_LC_10_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i15_LC_10_19_7  (
            .in0(_gnd_net_),
            .in1(N__39828),
            .in2(N__40520),
            .in3(N__39813),
            .lcout(encoder0_position_15),
            .ltout(),
            .carryin(\quad_counter0.n13109 ),
            .carryout(\quad_counter0.n13110 ),
            .clk(N__56202),
            .ce(N__40303),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i16_LC_10_20_0 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i16_LC_10_20_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i16_LC_10_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i16_LC_10_20_0  (
            .in0(_gnd_net_),
            .in1(N__40484),
            .in2(N__45757),
            .in3(N__39810),
            .lcout(encoder0_position_16),
            .ltout(),
            .carryin(bfn_10_20_0_),
            .carryout(\quad_counter0.n13111 ),
            .clk(N__56205),
            .ce(N__40304),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i17_LC_10_20_1 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i17_LC_10_20_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i17_LC_10_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i17_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(N__41919),
            .in2(N__40521),
            .in3(N__39807),
            .lcout(encoder0_position_17),
            .ltout(),
            .carryin(\quad_counter0.n13111 ),
            .carryout(\quad_counter0.n13112 ),
            .clk(N__56205),
            .ce(N__40304),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i18_LC_10_20_2 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i18_LC_10_20_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i18_LC_10_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i18_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(N__40488),
            .in2(N__43656),
            .in3(N__39804),
            .lcout(encoder0_position_18),
            .ltout(),
            .carryin(\quad_counter0.n13112 ),
            .carryout(\quad_counter0.n13113 ),
            .clk(N__56205),
            .ce(N__40304),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i19_LC_10_20_3 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i19_LC_10_20_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i19_LC_10_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i19_LC_10_20_3  (
            .in0(_gnd_net_),
            .in1(N__39800),
            .in2(N__40522),
            .in3(N__39780),
            .lcout(encoder0_position_19),
            .ltout(),
            .carryin(\quad_counter0.n13113 ),
            .carryout(\quad_counter0.n13114 ),
            .clk(N__56205),
            .ce(N__40304),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i20_LC_10_20_4 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i20_LC_10_20_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i20_LC_10_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i20_LC_10_20_4  (
            .in0(_gnd_net_),
            .in1(N__40492),
            .in2(N__47711),
            .in3(N__39777),
            .lcout(encoder0_position_20),
            .ltout(),
            .carryin(\quad_counter0.n13114 ),
            .carryout(\quad_counter0.n13115 ),
            .clk(N__56205),
            .ce(N__40304),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i21_LC_10_20_5 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i21_LC_10_20_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i21_LC_10_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i21_LC_10_20_5  (
            .in0(_gnd_net_),
            .in1(N__52408),
            .in2(N__40523),
            .in3(N__39774),
            .lcout(encoder0_position_21),
            .ltout(),
            .carryin(\quad_counter0.n13115 ),
            .carryout(\quad_counter0.n13116 ),
            .clk(N__56205),
            .ce(N__40304),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i22_LC_10_20_6 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i22_LC_10_20_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i22_LC_10_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i22_LC_10_20_6  (
            .in0(_gnd_net_),
            .in1(N__40496),
            .in2(N__47369),
            .in3(N__39771),
            .lcout(encoder0_position_22),
            .ltout(),
            .carryin(\quad_counter0.n13116 ),
            .carryout(\quad_counter0.n13117 ),
            .clk(N__56205),
            .ce(N__40304),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i23_LC_10_20_7 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i23_LC_10_20_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i23_LC_10_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i23_LC_10_20_7  (
            .in0(_gnd_net_),
            .in1(N__43837),
            .in2(N__40524),
            .in3(N__39768),
            .lcout(encoder0_position_23),
            .ltout(),
            .carryin(\quad_counter0.n13117 ),
            .carryout(\quad_counter0.n13118 ),
            .clk(N__56205),
            .ce(N__40304),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i24_LC_10_21_0 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i24_LC_10_21_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i24_LC_10_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i24_LC_10_21_0  (
            .in0(_gnd_net_),
            .in1(N__40500),
            .in2(N__43809),
            .in3(N__39855),
            .lcout(encoder0_position_24),
            .ltout(),
            .carryin(bfn_10_21_0_),
            .carryout(\quad_counter0.n13119 ),
            .clk(N__56206),
            .ce(N__40302),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i25_LC_10_21_1 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i25_LC_10_21_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i25_LC_10_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i25_LC_10_21_1  (
            .in0(_gnd_net_),
            .in1(N__43909),
            .in2(N__40525),
            .in3(N__39852),
            .lcout(encoder0_position_25),
            .ltout(),
            .carryin(\quad_counter0.n13119 ),
            .carryout(\quad_counter0.n13120 ),
            .clk(N__56206),
            .ce(N__40302),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i26_LC_10_21_2 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i26_LC_10_21_2 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i26_LC_10_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i26_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(N__40504),
            .in2(N__41828),
            .in3(N__39849),
            .lcout(encoder0_position_26),
            .ltout(),
            .carryin(\quad_counter0.n13120 ),
            .carryout(\quad_counter0.n13121 ),
            .clk(N__56206),
            .ce(N__40302),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i27_LC_10_21_3 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i27_LC_10_21_3 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i27_LC_10_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i27_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(N__41785),
            .in2(N__40526),
            .in3(N__39846),
            .lcout(encoder0_position_27),
            .ltout(),
            .carryin(\quad_counter0.n13121 ),
            .carryout(\quad_counter0.n13122 ),
            .clk(N__56206),
            .ce(N__40302),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i28_LC_10_21_4 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i28_LC_10_21_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i28_LC_10_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i28_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(N__40508),
            .in2(N__42073),
            .in3(N__39843),
            .lcout(encoder0_position_28),
            .ltout(),
            .carryin(\quad_counter0.n13122 ),
            .carryout(\quad_counter0.n13123 ),
            .clk(N__56206),
            .ce(N__40302),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i29_LC_10_21_5 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i29_LC_10_21_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i29_LC_10_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i29_LC_10_21_5  (
            .in0(_gnd_net_),
            .in1(N__41954),
            .in2(N__40527),
            .in3(N__39840),
            .lcout(encoder0_position_29),
            .ltout(),
            .carryin(\quad_counter0.n13123 ),
            .carryout(\quad_counter0.n13124 ),
            .clk(N__56206),
            .ce(N__40302),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i30_LC_10_21_6 .C_ON=1'b1;
    defparam \quad_counter0.position_659__i30_LC_10_21_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i30_LC_10_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \quad_counter0.position_659__i30_LC_10_21_6  (
            .in0(_gnd_net_),
            .in1(N__40512),
            .in2(N__42019),
            .in3(N__39837),
            .lcout(encoder0_position_30),
            .ltout(),
            .carryin(\quad_counter0.n13124 ),
            .carryout(\quad_counter0.n13125 ),
            .clk(N__56206),
            .ce(N__40302),
            .sr(_gnd_net_));
    defparam \quad_counter0.position_659__i31_LC_10_21_7 .C_ON=1'b0;
    defparam \quad_counter0.position_659__i31_LC_10_21_7 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.position_659__i31_LC_10_21_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \quad_counter0.position_659__i31_LC_10_21_7  (
            .in0(N__40513),
            .in1(N__49540),
            .in2(_gnd_net_),
            .in3(N__39834),
            .lcout(encoder0_position_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56206),
            .ce(N__40302),
            .sr(_gnd_net_));
    defparam add_741_2_lut_LC_10_22_0.C_ON=1'b1;
    defparam add_741_2_lut_LC_10_22_0.SEQ_MODE=4'b0000;
    defparam add_741_2_lut_LC_10_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_741_2_lut_LC_10_22_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42282),
            .in3(N__39831),
            .lcout(n2566),
            .ltout(),
            .carryin(bfn_10_22_0_),
            .carryout(n12496),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_741_3_lut_LC_10_22_1.C_ON=1'b1;
    defparam add_741_3_lut_LC_10_22_1.SEQ_MODE=4'b0000;
    defparam add_741_3_lut_LC_10_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_741_3_lut_LC_10_22_1 (
            .in0(_gnd_net_),
            .in1(N__54700),
            .in2(N__40029),
            .in3(N__39900),
            .lcout(n2565),
            .ltout(),
            .carryin(n12496),
            .carryout(n12497),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_741_4_lut_LC_10_22_2.C_ON=1'b1;
    defparam add_741_4_lut_LC_10_22_2.SEQ_MODE=4'b0000;
    defparam add_741_4_lut_LC_10_22_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_741_4_lut_LC_10_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40047),
            .in3(N__39897),
            .lcout(n2564),
            .ltout(),
            .carryin(n12497),
            .carryout(n12498),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_741_5_lut_LC_10_22_3.C_ON=1'b1;
    defparam add_741_5_lut_LC_10_22_3.SEQ_MODE=4'b0000;
    defparam add_741_5_lut_LC_10_22_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_741_5_lut_LC_10_22_3 (
            .in0(_gnd_net_),
            .in1(N__54701),
            .in2(N__41928),
            .in3(N__39894),
            .lcout(n2563),
            .ltout(),
            .carryin(n12498),
            .carryout(n12499),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_741_6_lut_LC_10_22_4.C_ON=1'b1;
    defparam add_741_6_lut_LC_10_22_4.SEQ_MODE=4'b0000;
    defparam add_741_6_lut_LC_10_22_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_741_6_lut_LC_10_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39873),
            .in3(N__39891),
            .lcout(n2562),
            .ltout(),
            .carryin(n12499),
            .carryout(n12500),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_741_7_lut_LC_10_22_5.C_ON=1'b0;
    defparam add_741_7_lut_LC_10_22_5.SEQ_MODE=4'b0000;
    defparam add_741_7_lut_LC_10_22_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 add_741_7_lut_LC_10_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40038),
            .in3(N__39888),
            .lcout(n2561),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10984_3_lut_LC_10_22_6.C_ON=1'b0;
    defparam i10984_3_lut_LC_10_22_6.SEQ_MODE=4'b0000;
    defparam i10984_3_lut_LC_10_22_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 i10984_3_lut_LC_10_22_6 (
            .in0(_gnd_net_),
            .in1(N__49496),
            .in2(N__41955),
            .in3(N__39879),
            .lcout(n830),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10983_3_lut_LC_10_22_7.C_ON=1'b0;
    defparam i10983_3_lut_LC_10_22_7.SEQ_MODE=4'b0000;
    defparam i10983_3_lut_LC_10_22_7.LUT_INIT=16'b1111110000110000;
    LogicCell40 i10983_3_lut_LC_10_22_7 (
            .in0(_gnd_net_),
            .in1(N__42193),
            .in2(N__42318),
            .in3(N__39885),
            .lcout(n13656),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i31_3_lut_LC_10_23_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i31_3_lut_LC_10_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i31_3_lut_LC_10_23_0.LUT_INIT=16'b1111101001010000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i31_3_lut_LC_10_23_0 (
            .in0(N__49547),
            .in1(_gnd_net_),
            .in2(N__42020),
            .in3(N__42220),
            .lcout(n403),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i27_3_lut_LC_10_23_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i27_3_lut_LC_10_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i27_3_lut_LC_10_23_1.LUT_INIT=16'b1111110000110000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i27_3_lut_LC_10_23_1 (
            .in0(_gnd_net_),
            .in1(N__49542),
            .in2(N__41829),
            .in3(N__41846),
            .lcout(n40),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut_LC_10_23_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut_LC_10_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut_LC_10_23_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut_LC_10_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47707),
            .lcout(n13_adj_631),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i29_3_lut_LC_10_23_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i29_3_lut_LC_10_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i29_3_lut_LC_10_23_3.LUT_INIT=16'b1111110000110000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i29_3_lut_LC_10_23_3 (
            .in0(_gnd_net_),
            .in1(N__49546),
            .in2(N__42075),
            .in3(N__42256),
            .lcout(n38),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_152_LC_10_23_4.C_ON=1'b0;
    defparam i1_3_lut_adj_152_LC_10_23_4.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_152_LC_10_23_4.LUT_INIT=16'b1100000000000000;
    LogicCell40 i1_3_lut_adj_152_LC_10_23_4 (
            .in0(_gnd_net_),
            .in1(N__42231),
            .in2(N__49598),
            .in3(N__42221),
            .lcout(n14568),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2181_2_lut_LC_10_23_5.C_ON=1'b0;
    defparam i2181_2_lut_LC_10_23_5.SEQ_MODE=4'b0000;
    defparam i2181_2_lut_LC_10_23_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 i2181_2_lut_LC_10_23_5 (
            .in0(_gnd_net_),
            .in1(N__49548),
            .in2(_gnd_net_),
            .in3(N__42428),
            .lcout(n402),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i28_3_lut_LC_10_23_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i28_3_lut_LC_10_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i28_3_lut_LC_10_23_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_mux_3_i28_3_lut_LC_10_23_6 (
            .in0(_gnd_net_),
            .in1(N__41787),
            .in2(N__49597),
            .in3(N__42340),
            .lcout(n39),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10981_3_lut_LC_10_23_7.C_ON=1'b0;
    defparam i10981_3_lut_LC_10_23_7.SEQ_MODE=4'b0000;
    defparam i10981_3_lut_LC_10_23_7.LUT_INIT=16'b1111110000110000;
    LogicCell40 i10981_3_lut_LC_10_23_7 (
            .in0(_gnd_net_),
            .in1(N__42194),
            .in2(N__42225),
            .in3(N__40020),
            .lcout(n13654),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dti_163_LC_10_24_1.C_ON=1'b0;
    defparam dti_163_LC_10_24_1.SEQ_MODE=4'b1000;
    defparam dti_163_LC_10_24_1.LUT_INIT=16'b1111111100110011;
    LogicCell40 dti_163_LC_10_24_1 (
            .in0(_gnd_net_),
            .in1(N__46601),
            .in2(_gnd_net_),
            .in3(N__46665),
            .lcout(dti),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56212),
            .ce(N__40014),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut_LC_10_24_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut_LC_10_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut_LC_10_24_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut_LC_10_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40002),
            .lcout(n22_adj_640),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut_LC_10_24_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut_LC_10_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut_LC_10_24_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut_LC_10_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39971),
            .lcout(n21_adj_639),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut_LC_10_24_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut_LC_10_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut_LC_10_24_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut_LC_10_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39930),
            .lcout(n20_adj_638),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut_LC_10_24_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut_LC_10_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut_LC_10_24_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut_LC_10_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43648),
            .lcout(n15_adj_633),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut_LC_10_24_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut_LC_10_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut_LC_10_24_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut_LC_10_24_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41786),
            .lcout(n6_adj_624),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.debounce_cnt_I_0_4_lut_LC_10_25_0 .C_ON=1'b0;
    defparam \quad_counter0.debounce_cnt_I_0_4_lut_LC_10_25_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.debounce_cnt_I_0_4_lut_LC_10_25_0 .LUT_INIT=16'b1000101010101000;
    LogicCell40 \quad_counter0.debounce_cnt_I_0_4_lut_LC_10_25_0  (
            .in0(N__46306),
            .in1(N__40362),
            .in2(N__46401),
            .in3(N__40542),
            .lcout(direction_N_537),
            .ltout(direction_N_537_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.direction_57_LC_10_25_1 .C_ON=1'b0;
    defparam \quad_counter0.direction_57_LC_10_25_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.direction_57_LC_10_25_1 .LUT_INIT=16'b0101110010101100;
    LogicCell40 \quad_counter0.direction_57_LC_10_25_1  (
            .in0(N__46400),
            .in1(N__40257),
            .in2(N__40260),
            .in3(N__46278),
            .lcout(n1302),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56215),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut_LC_10_25_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut_LC_10_25_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut_LC_10_25_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut_LC_10_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43916),
            .lcout(n8_adj_626),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut_LC_10_25_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut_LC_10_25_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut_LC_10_25_3.LUT_INIT=16'b0000111100001111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut_LC_10_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42074),
            .in3(_gnd_net_),
            .lcout(n5_adj_623),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut_LC_10_25_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut_LC_10_25_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut_LC_10_25_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut_LC_10_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49541),
            .lcout(n2_adj_620),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut_LC_10_25_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut_LC_10_25_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut_LC_10_25_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut_LC_10_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43801),
            .lcout(n9_adj_627),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i6_1_lut_LC_10_25_6.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i6_1_lut_LC_10_25_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i6_1_lut_LC_10_25_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i6_1_lut_LC_10_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40056),
            .lcout(n20_adj_556),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i2_1_lut_LC_10_25_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i2_1_lut_LC_10_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i2_1_lut_LC_10_25_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i2_1_lut_LC_10_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40371),
            .lcout(n24_adj_552),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i8_3_lut_3_lut_LC_10_26_0.C_ON=1'b0;
    defparam LessThan_299_i8_3_lut_3_lut_LC_10_26_0.SEQ_MODE=4'b0000;
    defparam LessThan_299_i8_3_lut_3_lut_LC_10_26_0.LUT_INIT=16'b1011101100100010;
    LogicCell40 LessThan_299_i8_3_lut_3_lut_LC_10_26_0 (
            .in0(N__42803),
            .in1(N__47979),
            .in2(_gnd_net_),
            .in3(N__40563),
            .lcout(n8_adj_657),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_prev_I_0_65_2_lut_LC_10_26_1 .C_ON=1'b0;
    defparam \quad_counter0.b_prev_I_0_65_2_lut_LC_10_26_1 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.b_prev_I_0_65_2_lut_LC_10_26_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \quad_counter0.b_prev_I_0_65_2_lut_LC_10_26_1  (
            .in0(_gnd_net_),
            .in1(N__46340),
            .in2(_gnd_net_),
            .in3(N__46277),
            .lcout(\quad_counter0.direction_N_540 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i10_1_lut_LC_10_26_2.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i10_1_lut_LC_10_26_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i10_1_lut_LC_10_26_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i10_1_lut_LC_10_26_2 (
            .in0(N__40356),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n16_adj_560),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i5_LC_10_26_3.C_ON=1'b0;
    defparam pwm_setpoint_i5_LC_10_26_3.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i5_LC_10_26_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 pwm_setpoint_i5_LC_10_26_3 (
            .in0(N__43968),
            .in1(N__42459),
            .in2(_gnd_net_),
            .in3(N__50907),
            .lcout(pwm_setpoint_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56216),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i21_1_lut_LC_10_26_4.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i21_1_lut_LC_10_26_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i21_1_lut_LC_10_26_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i21_1_lut_LC_10_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40347),
            .lcout(n5_adj_571),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i7_LC_10_26_5.C_ON=1'b0;
    defparam pwm_setpoint_i7_LC_10_26_5.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i7_LC_10_26_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 pwm_setpoint_i7_LC_10_26_5 (
            .in0(N__42441),
            .in1(N__50908),
            .in2(_gnd_net_),
            .in3(N__44340),
            .lcout(pwm_setpoint_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56216),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i4_LC_10_26_6.C_ON=1'b0;
    defparam pwm_setpoint_i4_LC_10_26_6.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i4_LC_10_26_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 pwm_setpoint_i4_LC_10_26_6 (
            .in0(N__50906),
            .in1(N__42474),
            .in2(_gnd_net_),
            .in3(N__43998),
            .lcout(pwm_setpoint_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56216),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i12_1_lut_LC_10_26_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i12_1_lut_LC_10_26_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i12_1_lut_LC_10_26_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i12_1_lut_LC_10_26_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40335),
            .lcout(n14_adj_562),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i13_LC_10_27_0.C_ON=1'b0;
    defparam pwm_setpoint_i13_LC_10_27_0.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i13_LC_10_27_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 pwm_setpoint_i13_LC_10_27_0 (
            .in0(N__50868),
            .in1(N__44151),
            .in2(_gnd_net_),
            .in3(N__42558),
            .lcout(pwm_setpoint_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56217),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i22_1_lut_LC_10_27_1.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i22_1_lut_LC_10_27_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i22_1_lut_LC_10_27_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i22_1_lut_LC_10_27_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40581),
            .lcout(n4_adj_572),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i20_1_lut_LC_10_27_2.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i20_1_lut_LC_10_27_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i20_1_lut_LC_10_27_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i20_1_lut_LC_10_27_2 (
            .in0(N__40572),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n6_adj_570),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i9_2_lut_LC_10_27_3.C_ON=1'b0;
    defparam LessThan_299_i9_2_lut_LC_10_27_3.SEQ_MODE=4'b0000;
    defparam LessThan_299_i9_2_lut_LC_10_27_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i9_2_lut_LC_10_27_3 (
            .in0(_gnd_net_),
            .in1(N__40562),
            .in2(_gnd_net_),
            .in3(N__48102),
            .lcout(n9_adj_658),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i23_1_lut_LC_10_27_4.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i23_1_lut_LC_10_27_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i23_1_lut_LC_10_27_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i23_1_lut_LC_10_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40551),
            .lcout(n3_adj_573),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i14_1_lut_LC_10_27_5.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i14_1_lut_LC_10_27_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i14_1_lut_LC_10_27_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i14_1_lut_LC_10_27_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44150),
            .lcout(n12_adj_584),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i11_LC_10_27_6.C_ON=1'b0;
    defparam pwm_setpoint_i11_LC_10_27_6.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i11_LC_10_27_6.LUT_INIT=16'b1110111001000100;
    LogicCell40 pwm_setpoint_i11_LC_10_27_6 (
            .in0(N__50867),
            .in1(N__44201),
            .in2(_gnd_net_),
            .in3(N__42576),
            .lcout(pwm_setpoint_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56217),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i8_LC_10_27_7.C_ON=1'b0;
    defparam pwm_setpoint_i8_LC_10_27_7.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i8_LC_10_27_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 pwm_setpoint_i8_LC_10_27_7 (
            .in0(N__44309),
            .in1(N__42627),
            .in2(_gnd_net_),
            .in3(N__50869),
            .lcout(pwm_setpoint_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56217),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.a_prev_51_LC_10_28_0 .C_ON=1'b0;
    defparam \quad_counter0.a_prev_51_LC_10_28_0 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_prev_51_LC_10_28_0 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \quad_counter0.a_prev_51_LC_10_28_0  (
            .in0(N__46395),
            .in1(N__40541),
            .in2(N__46308),
            .in3(N__46356),
            .lcout(\quad_counter0.a_prev ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56220),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_prev_I_0_63_2_lut_LC_10_28_5 .C_ON=1'b0;
    defparam \quad_counter0.b_prev_I_0_63_2_lut_LC_10_28_5 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.b_prev_I_0_63_2_lut_LC_10_28_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \quad_counter0.b_prev_I_0_63_2_lut_LC_10_28_5  (
            .in0(_gnd_net_),
            .in1(N__46394),
            .in2(_gnd_net_),
            .in3(N__46270),
            .lcout(\quad_counter0.direction_N_536 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.debounce_cnt_50_LC_10_28_6 .C_ON=1'b0;
    defparam \quad_counter0.debounce_cnt_50_LC_10_28_6 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.debounce_cnt_50_LC_10_28_6 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \quad_counter0.debounce_cnt_50_LC_10_28_6  (
            .in0(N__46396),
            .in1(N__46457),
            .in2(N__46347),
            .in3(N__46428),
            .lcout(\quad_counter0.debounce_cnt ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56220),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i0_LC_10_29_0.C_ON=1'b1;
    defparam blink_counter_663__i0_LC_10_29_0.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i0_LC_10_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i0_LC_10_29_0 (
            .in0(_gnd_net_),
            .in1(N__40644),
            .in2(_gnd_net_),
            .in3(N__40638),
            .lcout(n26_adj_703),
            .ltout(),
            .carryin(bfn_10_29_0_),
            .carryout(n13070),
            .clk(N__56224),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i1_LC_10_29_1.C_ON=1'b1;
    defparam blink_counter_663__i1_LC_10_29_1.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i1_LC_10_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i1_LC_10_29_1 (
            .in0(_gnd_net_),
            .in1(N__40635),
            .in2(_gnd_net_),
            .in3(N__40629),
            .lcout(n25_adj_702),
            .ltout(),
            .carryin(n13070),
            .carryout(n13071),
            .clk(N__56224),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i2_LC_10_29_2.C_ON=1'b1;
    defparam blink_counter_663__i2_LC_10_29_2.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i2_LC_10_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i2_LC_10_29_2 (
            .in0(_gnd_net_),
            .in1(N__40626),
            .in2(_gnd_net_),
            .in3(N__40620),
            .lcout(n24_adj_701),
            .ltout(),
            .carryin(n13071),
            .carryout(n13072),
            .clk(N__56224),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i3_LC_10_29_3.C_ON=1'b1;
    defparam blink_counter_663__i3_LC_10_29_3.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i3_LC_10_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i3_LC_10_29_3 (
            .in0(_gnd_net_),
            .in1(N__40617),
            .in2(_gnd_net_),
            .in3(N__40611),
            .lcout(n23_adj_700),
            .ltout(),
            .carryin(n13072),
            .carryout(n13073),
            .clk(N__56224),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i4_LC_10_29_4.C_ON=1'b1;
    defparam blink_counter_663__i4_LC_10_29_4.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i4_LC_10_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i4_LC_10_29_4 (
            .in0(_gnd_net_),
            .in1(N__40608),
            .in2(_gnd_net_),
            .in3(N__40602),
            .lcout(n22_adj_699),
            .ltout(),
            .carryin(n13073),
            .carryout(n13074),
            .clk(N__56224),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i5_LC_10_29_5.C_ON=1'b1;
    defparam blink_counter_663__i5_LC_10_29_5.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i5_LC_10_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i5_LC_10_29_5 (
            .in0(_gnd_net_),
            .in1(N__40599),
            .in2(_gnd_net_),
            .in3(N__40593),
            .lcout(n21_adj_698),
            .ltout(),
            .carryin(n13074),
            .carryout(n13075),
            .clk(N__56224),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i6_LC_10_29_6.C_ON=1'b1;
    defparam blink_counter_663__i6_LC_10_29_6.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i6_LC_10_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i6_LC_10_29_6 (
            .in0(_gnd_net_),
            .in1(N__40590),
            .in2(_gnd_net_),
            .in3(N__40584),
            .lcout(n20_adj_697),
            .ltout(),
            .carryin(n13075),
            .carryout(n13076),
            .clk(N__56224),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i7_LC_10_29_7.C_ON=1'b1;
    defparam blink_counter_663__i7_LC_10_29_7.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i7_LC_10_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i7_LC_10_29_7 (
            .in0(_gnd_net_),
            .in1(N__40725),
            .in2(_gnd_net_),
            .in3(N__40719),
            .lcout(n19_adj_696),
            .ltout(),
            .carryin(n13076),
            .carryout(n13077),
            .clk(N__56224),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i8_LC_10_30_0.C_ON=1'b1;
    defparam blink_counter_663__i8_LC_10_30_0.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i8_LC_10_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i8_LC_10_30_0 (
            .in0(_gnd_net_),
            .in1(N__40716),
            .in2(_gnd_net_),
            .in3(N__40710),
            .lcout(n18_adj_695),
            .ltout(),
            .carryin(bfn_10_30_0_),
            .carryout(n13078),
            .clk(N__56229),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i9_LC_10_30_1.C_ON=1'b1;
    defparam blink_counter_663__i9_LC_10_30_1.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i9_LC_10_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i9_LC_10_30_1 (
            .in0(_gnd_net_),
            .in1(N__40707),
            .in2(_gnd_net_),
            .in3(N__40701),
            .lcout(n17_adj_694),
            .ltout(),
            .carryin(n13078),
            .carryout(n13079),
            .clk(N__56229),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i10_LC_10_30_2.C_ON=1'b1;
    defparam blink_counter_663__i10_LC_10_30_2.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i10_LC_10_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i10_LC_10_30_2 (
            .in0(_gnd_net_),
            .in1(N__40698),
            .in2(_gnd_net_),
            .in3(N__40692),
            .lcout(n16_adj_693),
            .ltout(),
            .carryin(n13079),
            .carryout(n13080),
            .clk(N__56229),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i11_LC_10_30_3.C_ON=1'b1;
    defparam blink_counter_663__i11_LC_10_30_3.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i11_LC_10_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i11_LC_10_30_3 (
            .in0(_gnd_net_),
            .in1(N__40689),
            .in2(_gnd_net_),
            .in3(N__40683),
            .lcout(n15_adj_692),
            .ltout(),
            .carryin(n13080),
            .carryout(n13081),
            .clk(N__56229),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i12_LC_10_30_4.C_ON=1'b1;
    defparam blink_counter_663__i12_LC_10_30_4.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i12_LC_10_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i12_LC_10_30_4 (
            .in0(_gnd_net_),
            .in1(N__40680),
            .in2(_gnd_net_),
            .in3(N__40674),
            .lcout(n14_adj_691),
            .ltout(),
            .carryin(n13081),
            .carryout(n13082),
            .clk(N__56229),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i13_LC_10_30_5.C_ON=1'b1;
    defparam blink_counter_663__i13_LC_10_30_5.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i13_LC_10_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i13_LC_10_30_5 (
            .in0(_gnd_net_),
            .in1(N__40671),
            .in2(_gnd_net_),
            .in3(N__40665),
            .lcout(n13_adj_690),
            .ltout(),
            .carryin(n13082),
            .carryout(n13083),
            .clk(N__56229),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i14_LC_10_30_6.C_ON=1'b1;
    defparam blink_counter_663__i14_LC_10_30_6.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i14_LC_10_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i14_LC_10_30_6 (
            .in0(_gnd_net_),
            .in1(N__40662),
            .in2(_gnd_net_),
            .in3(N__40656),
            .lcout(n12_adj_689),
            .ltout(),
            .carryin(n13083),
            .carryout(n13084),
            .clk(N__56229),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i15_LC_10_30_7.C_ON=1'b1;
    defparam blink_counter_663__i15_LC_10_30_7.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i15_LC_10_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i15_LC_10_30_7 (
            .in0(_gnd_net_),
            .in1(N__40653),
            .in2(_gnd_net_),
            .in3(N__40647),
            .lcout(n11_adj_688),
            .ltout(),
            .carryin(n13084),
            .carryout(n13085),
            .clk(N__56229),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i16_LC_10_31_0.C_ON=1'b1;
    defparam blink_counter_663__i16_LC_10_31_0.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i16_LC_10_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i16_LC_10_31_0 (
            .in0(_gnd_net_),
            .in1(N__40830),
            .in2(_gnd_net_),
            .in3(N__40824),
            .lcout(n10_adj_687),
            .ltout(),
            .carryin(bfn_10_31_0_),
            .carryout(n13086),
            .clk(N__56236),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i17_LC_10_31_1.C_ON=1'b1;
    defparam blink_counter_663__i17_LC_10_31_1.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i17_LC_10_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i17_LC_10_31_1 (
            .in0(_gnd_net_),
            .in1(N__40821),
            .in2(_gnd_net_),
            .in3(N__40815),
            .lcout(n9_adj_686),
            .ltout(),
            .carryin(n13086),
            .carryout(n13087),
            .clk(N__56236),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i18_LC_10_31_2.C_ON=1'b1;
    defparam blink_counter_663__i18_LC_10_31_2.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i18_LC_10_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i18_LC_10_31_2 (
            .in0(_gnd_net_),
            .in1(N__40812),
            .in2(_gnd_net_),
            .in3(N__40806),
            .lcout(n8_adj_685),
            .ltout(),
            .carryin(n13087),
            .carryout(n13088),
            .clk(N__56236),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i19_LC_10_31_3.C_ON=1'b1;
    defparam blink_counter_663__i19_LC_10_31_3.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i19_LC_10_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i19_LC_10_31_3 (
            .in0(_gnd_net_),
            .in1(N__40803),
            .in2(_gnd_net_),
            .in3(N__40797),
            .lcout(n7_adj_684),
            .ltout(),
            .carryin(n13088),
            .carryout(n13089),
            .clk(N__56236),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i20_LC_10_31_4.C_ON=1'b1;
    defparam blink_counter_663__i20_LC_10_31_4.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i20_LC_10_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i20_LC_10_31_4 (
            .in0(_gnd_net_),
            .in1(N__40794),
            .in2(_gnd_net_),
            .in3(N__40788),
            .lcout(n6_adj_683),
            .ltout(),
            .carryin(n13089),
            .carryout(n13090),
            .clk(N__56236),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i21_LC_10_31_5.C_ON=1'b1;
    defparam blink_counter_663__i21_LC_10_31_5.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i21_LC_10_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i21_LC_10_31_5 (
            .in0(_gnd_net_),
            .in1(N__40780),
            .in2(_gnd_net_),
            .in3(N__40767),
            .lcout(blink_counter_21),
            .ltout(),
            .carryin(n13090),
            .carryout(n13091),
            .clk(N__56236),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i22_LC_10_31_6.C_ON=1'b1;
    defparam blink_counter_663__i22_LC_10_31_6.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i22_LC_10_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i22_LC_10_31_6 (
            .in0(_gnd_net_),
            .in1(N__40762),
            .in2(_gnd_net_),
            .in3(N__40749),
            .lcout(blink_counter_22),
            .ltout(),
            .carryin(n13091),
            .carryout(n13092),
            .clk(N__56236),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i23_LC_10_31_7.C_ON=1'b1;
    defparam blink_counter_663__i23_LC_10_31_7.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i23_LC_10_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i23_LC_10_31_7 (
            .in0(_gnd_net_),
            .in1(N__40741),
            .in2(_gnd_net_),
            .in3(N__40728),
            .lcout(blink_counter_23),
            .ltout(),
            .carryin(n13092),
            .carryout(n13093),
            .clk(N__56236),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i24_LC_10_32_0.C_ON=1'b1;
    defparam blink_counter_663__i24_LC_10_32_0.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i24_LC_10_32_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i24_LC_10_32_0 (
            .in0(_gnd_net_),
            .in1(N__40990),
            .in2(_gnd_net_),
            .in3(N__40977),
            .lcout(blink_counter_24),
            .ltout(),
            .carryin(bfn_10_32_0_),
            .carryout(n13094),
            .clk(N__56242),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_663__i25_LC_10_32_1.C_ON=1'b0;
    defparam blink_counter_663__i25_LC_10_32_1.SEQ_MODE=4'b1000;
    defparam blink_counter_663__i25_LC_10_32_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_663__i25_LC_10_32_1 (
            .in0(_gnd_net_),
            .in1(N__40970),
            .in2(_gnd_net_),
            .in3(N__40974),
            .lcout(blink_counter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56242),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1185_3_lut_LC_11_16_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1185_3_lut_LC_11_16_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1185_3_lut_LC_11_16_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i1185_3_lut_LC_11_16_2 (
            .in0(N__43692),
            .in1(N__43347),
            .in2(_gnd_net_),
            .in3(N__45476),
            .lcout(n1833),
            .ltout(n1833_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10012_4_lut_LC_11_16_3.C_ON=1'b0;
    defparam i10012_4_lut_LC_11_16_3.SEQ_MODE=4'b0000;
    defparam i10012_4_lut_LC_11_16_3.LUT_INIT=16'b1111111011001100;
    LogicCell40 i10012_4_lut_LC_11_16_3 (
            .in0(N__40949),
            .in1(N__40847),
            .in2(N__40959),
            .in3(N__40879),
            .lcout(n11989),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1184_3_lut_LC_11_16_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1184_3_lut_LC_11_16_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1184_3_lut_LC_11_16_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1184_3_lut_LC_11_16_5 (
            .in0(_gnd_net_),
            .in1(N__43332),
            .in2(N__45499),
            .in3(N__45537),
            .lcout(n1832),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_2_lut_LC_11_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_2_lut_LC_11_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_2_lut_LC_11_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_2_lut_LC_11_17_0 (
            .in0(_gnd_net_),
            .in1(N__40948),
            .in2(_gnd_net_),
            .in3(N__40914),
            .lcout(n1901),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(n12606),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_3_lut_LC_11_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_3_lut_LC_11_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_3_lut_LC_11_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_3_lut_LC_11_17_1 (
            .in0(_gnd_net_),
            .in1(N__55285),
            .in2(N__40910),
            .in3(N__40887),
            .lcout(n1900),
            .ltout(),
            .carryin(n12606),
            .carryout(n12607),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_4_lut_LC_11_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_4_lut_LC_11_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_4_lut_LC_11_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_4_lut_LC_11_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40884),
            .in3(N__40854),
            .lcout(n1899),
            .ltout(),
            .carryin(n12607),
            .carryout(n12608),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_5_lut_LC_11_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_5_lut_LC_11_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_5_lut_LC_11_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_5_lut_LC_11_17_3 (
            .in0(_gnd_net_),
            .in1(N__55286),
            .in2(N__40851),
            .in3(N__41058),
            .lcout(n1898),
            .ltout(),
            .carryin(n12608),
            .carryout(n12609),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_6_lut_LC_11_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_6_lut_LC_11_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_6_lut_LC_11_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_6_lut_LC_11_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43111),
            .in3(N__41049),
            .lcout(n1897),
            .ltout(),
            .carryin(n12609),
            .carryout(n12610),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_7_lut_LC_11_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_7_lut_LC_11_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_7_lut_LC_11_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_7_lut_LC_11_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41667),
            .in3(N__41040),
            .lcout(n1896),
            .ltout(),
            .carryin(n12610),
            .carryout(n12611),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_8_lut_LC_11_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_8_lut_LC_11_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_8_lut_LC_11_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_8_lut_LC_11_17_6 (
            .in0(_gnd_net_),
            .in1(N__55087),
            .in2(N__42848),
            .in3(N__41037),
            .lcout(n1895),
            .ltout(),
            .carryin(n12611),
            .carryout(n12612),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_9_lut_LC_11_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_9_lut_LC_11_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_9_lut_LC_11_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_9_lut_LC_11_17_7 (
            .in0(_gnd_net_),
            .in1(N__55287),
            .in2(N__43169),
            .in3(N__41034),
            .lcout(n1894),
            .ltout(),
            .carryin(n12612),
            .carryout(n12613),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_10_lut_LC_11_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_10_lut_LC_11_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_10_lut_LC_11_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_10_lut_LC_11_18_0 (
            .in0(_gnd_net_),
            .in1(N__55281),
            .in2(N__43082),
            .in3(N__41025),
            .lcout(n1893),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(n12614),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_11_lut_LC_11_18_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_11_lut_LC_11_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_11_lut_LC_11_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_11_lut_LC_11_18_1 (
            .in0(_gnd_net_),
            .in1(N__54955),
            .in2(N__42878),
            .in3(N__41022),
            .lcout(n1892),
            .ltout(),
            .carryin(n12614),
            .carryout(n12615),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_12_lut_LC_11_18_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_12_lut_LC_11_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_12_lut_LC_11_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_12_lut_LC_11_18_2 (
            .in0(_gnd_net_),
            .in1(N__55282),
            .in2(N__43058),
            .in3(N__41010),
            .lcout(n1891),
            .ltout(),
            .carryin(n12615),
            .carryout(n12616),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_13_lut_LC_11_18_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_13_lut_LC_11_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_13_lut_LC_11_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_13_lut_LC_11_18_3 (
            .in0(_gnd_net_),
            .in1(N__54956),
            .in2(N__43031),
            .in3(N__40995),
            .lcout(n1890),
            .ltout(),
            .carryin(n12616),
            .carryout(n12617),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_14_lut_LC_11_18_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_14_lut_LC_11_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_14_lut_LC_11_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_14_lut_LC_11_18_4 (
            .in0(_gnd_net_),
            .in1(N__55283),
            .in2(N__41087),
            .in3(N__41181),
            .lcout(n1889),
            .ltout(),
            .carryin(n12617),
            .carryout(n12618),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_15_lut_LC_11_18_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_15_lut_LC_11_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_15_lut_LC_11_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_15_lut_LC_11_18_5 (
            .in0(_gnd_net_),
            .in1(N__54957),
            .in2(N__43142),
            .in3(N__41178),
            .lcout(n1888),
            .ltout(),
            .carryin(n12618),
            .carryout(n12619),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_16_lut_LC_11_18_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_16_lut_LC_11_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_16_lut_LC_11_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_16_lut_LC_11_18_6 (
            .in0(_gnd_net_),
            .in1(N__55284),
            .in2(N__43193),
            .in3(N__41163),
            .lcout(n1887),
            .ltout(),
            .carryin(n12619),
            .carryout(n12620),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_17_lut_LC_11_18_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1235_17_lut_LC_11_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_17_lut_LC_11_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1235_17_lut_LC_11_18_7 (
            .in0(_gnd_net_),
            .in1(N__54958),
            .in2(N__41228),
            .in3(N__41148),
            .lcout(n1886),
            .ltout(),
            .carryin(n12620),
            .carryout(n12621),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1235_18_lut_LC_11_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1235_18_lut_LC_11_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1235_18_lut_LC_11_19_0.LUT_INIT=16'b1010010101011010;
    LogicCell40 encoder0_position_31__I_0_add_1235_18_lut_LC_11_19_0 (
            .in0(N__55280),
            .in1(_gnd_net_),
            .in2(N__43749),
            .in3(N__41145),
            .lcout(n1885),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1244_3_lut_LC_11_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1244_3_lut_LC_11_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1244_3_lut_LC_11_19_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1244_3_lut_LC_11_19_1 (
            .in0(_gnd_net_),
            .in1(N__42879),
            .in2(N__41142),
            .in3(N__41503),
            .lcout(n1924),
            .ltout(n1924_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_140_LC_11_19_2.C_ON=1'b0;
    defparam i1_3_lut_adj_140_LC_11_19_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_140_LC_11_19_2.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_140_LC_11_19_2 (
            .in0(_gnd_net_),
            .in1(N__41725),
            .in2(N__41106),
            .in3(N__41683),
            .lcout(n14438),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1174_3_lut_LC_11_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1174_3_lut_LC_11_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1174_3_lut_LC_11_19_3.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1174_3_lut_LC_11_19_3 (
            .in0(N__43467),
            .in1(_gnd_net_),
            .in2(N__45506),
            .in3(N__43487),
            .lcout(n1822),
            .ltout(n1822_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_139_LC_11_19_4.C_ON=1'b0;
    defparam i1_3_lut_adj_139_LC_11_19_4.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_139_LC_11_19_4.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_139_LC_11_19_4 (
            .in0(_gnd_net_),
            .in1(N__43186),
            .in2(N__41070),
            .in3(N__43135),
            .lcout(n14534),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1247_3_lut_LC_11_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1247_3_lut_LC_11_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1247_3_lut_LC_11_19_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1247_3_lut_LC_11_19_5 (
            .in0(_gnd_net_),
            .in1(N__42849),
            .in2(N__41757),
            .in3(N__41502),
            .lcout(n1927),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1246_3_lut_LC_11_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1246_3_lut_LC_11_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1246_3_lut_LC_11_19_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1246_3_lut_LC_11_19_7 (
            .in0(_gnd_net_),
            .in1(N__41712),
            .in2(N__43170),
            .in3(N__41501),
            .lcout(n1926),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1181_3_lut_LC_11_20_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1181_3_lut_LC_11_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1181_3_lut_LC_11_20_0.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1181_3_lut_LC_11_20_0 (
            .in0(_gnd_net_),
            .in1(N__43242),
            .in2(N__45501),
            .in3(N__45702),
            .lcout(n1829),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1237_3_lut_LC_11_20_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1237_3_lut_LC_11_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1237_3_lut_LC_11_20_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1237_3_lut_LC_11_20_2 (
            .in0(_gnd_net_),
            .in1(N__43735),
            .in2(N__41646),
            .in3(N__41505),
            .lcout(n1917),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i4_3_lut_LC_11_20_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i4_3_lut_LC_11_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i4_3_lut_LC_11_20_3.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i4_3_lut_LC_11_20_3 (
            .in0(N__41613),
            .in1(_gnd_net_),
            .in2(N__41601),
            .in3(N__49539),
            .lcout(n316),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1240_3_lut_LC_11_20_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1240_3_lut_LC_11_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1240_3_lut_LC_11_20_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1240_3_lut_LC_11_20_6 (
            .in0(_gnd_net_),
            .in1(N__41532),
            .in2(N__43143),
            .in3(N__41504),
            .lcout(n1920),
            .ltout(n1920_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1307_3_lut_LC_11_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1307_3_lut_LC_11_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1307_3_lut_LC_11_20_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1307_3_lut_LC_11_20_7 (
            .in0(_gnd_net_),
            .in1(N__41397),
            .in2(N__41385),
            .in3(N__41378),
            .lcout(n2019),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1171_3_lut_LC_11_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1171_3_lut_LC_11_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1171_3_lut_LC_11_21_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1171_3_lut_LC_11_21_0 (
            .in0(_gnd_net_),
            .in1(N__43368),
            .in2(N__43395),
            .in3(N__45502),
            .lcout(n1819),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i18_3_lut_LC_11_21_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i18_3_lut_LC_11_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i18_3_lut_LC_11_21_2.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_mux_3_i18_3_lut_LC_11_21_2 (
            .in0(N__41918),
            .in1(_gnd_net_),
            .in2(N__49553),
            .in3(N__41967),
            .lcout(n302),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i30_3_lut_LC_11_21_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i30_3_lut_LC_11_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i30_3_lut_LC_11_21_4.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_mux_3_i30_3_lut_LC_11_21_4 (
            .in0(_gnd_net_),
            .in1(N__41950),
            .in2(N__49552),
            .in3(N__42316),
            .lcout(n404),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut_LC_11_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut_LC_11_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut_LC_11_21_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut_LC_11_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41917),
            .lcout(n16_adj_634),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut_LC_11_21_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut_LC_11_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut_LC_11_21_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut_LC_11_21_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41817),
            .lcout(n7_adj_625),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut_LC_11_21_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut_LC_11_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut_LC_11_21_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut_LC_11_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42003),
            .lcout(n3_adj_621),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10989_3_lut_LC_11_22_0.C_ON=1'b0;
    defparam i10989_3_lut_LC_11_22_0.SEQ_MODE=4'b0000;
    defparam i10989_3_lut_LC_11_22_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 i10989_3_lut_LC_11_22_0 (
            .in0(_gnd_net_),
            .in1(N__41859),
            .in2(N__41853),
            .in3(N__42188),
            .lcout(),
            .ltout(n13662_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12421_3_lut_LC_11_22_1.C_ON=1'b0;
    defparam i12421_3_lut_LC_11_22_1.SEQ_MODE=4'b0000;
    defparam i12421_3_lut_LC_11_22_1.LUT_INIT=16'b1111001111000000;
    LogicCell40 i12421_3_lut_LC_11_22_1 (
            .in0(_gnd_net_),
            .in1(N__49493),
            .in2(N__41832),
            .in3(N__41821),
            .lcout(n833),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10987_3_lut_LC_11_22_2.C_ON=1'b0;
    defparam i10987_3_lut_LC_11_22_2.SEQ_MODE=4'b0000;
    defparam i10987_3_lut_LC_11_22_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 i10987_3_lut_LC_11_22_2 (
            .in0(_gnd_net_),
            .in1(N__42348),
            .in2(N__41796),
            .in3(N__42189),
            .lcout(),
            .ltout(n13660_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10988_3_lut_LC_11_22_3.C_ON=1'b0;
    defparam i10988_3_lut_LC_11_22_3.SEQ_MODE=4'b0000;
    defparam i10988_3_lut_LC_11_22_3.LUT_INIT=16'b1111000010101010;
    LogicCell40 i10988_3_lut_LC_11_22_3 (
            .in0(N__41784),
            .in1(_gnd_net_),
            .in2(N__41760),
            .in3(N__49494),
            .lcout(n832),
            .ltout(n832_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10050_4_lut_LC_11_22_4.C_ON=1'b0;
    defparam i10050_4_lut_LC_11_22_4.SEQ_MODE=4'b0000;
    defparam i10050_4_lut_LC_11_22_4.LUT_INIT=16'b1111111111100000;
    LogicCell40 i10050_4_lut_LC_11_22_4 (
            .in0(N__43585),
            .in1(N__43875),
            .in2(N__42087),
            .in3(N__42151),
            .lcout(n12027),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10985_3_lut_LC_11_22_5.C_ON=1'b0;
    defparam i10985_3_lut_LC_11_22_5.SEQ_MODE=4'b0000;
    defparam i10985_3_lut_LC_11_22_5.LUT_INIT=16'b1111110000001100;
    LogicCell40 i10985_3_lut_LC_11_22_5 (
            .in0(_gnd_net_),
            .in1(N__42264),
            .in2(N__42195),
            .in3(N__42084),
            .lcout(),
            .ltout(n13658_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10986_3_lut_LC_11_22_6.C_ON=1'b0;
    defparam i10986_3_lut_LC_11_22_6.SEQ_MODE=4'b0000;
    defparam i10986_3_lut_LC_11_22_6.LUT_INIT=16'b1111010110100000;
    LogicCell40 i10986_3_lut_LC_11_22_6 (
            .in0(N__49495),
            .in1(_gnd_net_),
            .in2(N__42078),
            .in3(N__42063),
            .lcout(n831),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i5_1_lut_LC_11_22_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i5_1_lut_LC_11_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i5_1_lut_LC_11_22_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i5_1_lut_LC_11_22_7 (
            .in0(N__42036),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n21_adj_555),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i569_3_lut_LC_11_23_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i569_3_lut_LC_11_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i569_3_lut_LC_11_23_0.LUT_INIT=16'b1111110000110000;
    LogicCell40 encoder0_position_31__I_0_i569_3_lut_LC_11_23_0 (
            .in0(_gnd_net_),
            .in1(N__44089),
            .in2(N__42125),
            .in3(N__42099),
            .lcout(n929),
            .ltout(n929_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_85_LC_11_23_1.C_ON=1'b0;
    defparam i1_2_lut_adj_85_LC_11_23_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_85_LC_11_23_1.LUT_INIT=16'b1111000000000000;
    LogicCell40 i1_2_lut_adj_85_LC_11_23_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42024),
            .in3(N__46096),
            .lcout(n14460),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10982_3_lut_LC_11_23_2.C_ON=1'b0;
    defparam i10982_3_lut_LC_11_23_2.SEQ_MODE=4'b0000;
    defparam i10982_3_lut_LC_11_23_2.LUT_INIT=16'b1111101001010000;
    LogicCell40 i10982_3_lut_LC_11_23_2 (
            .in0(N__49600),
            .in1(_gnd_net_),
            .in2(N__42021),
            .in3(N__41985),
            .lcout(n829),
            .ltout(n829_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10150_4_lut_LC_11_23_3.C_ON=1'b0;
    defparam i10150_4_lut_LC_11_23_3.SEQ_MODE=4'b0000;
    defparam i10150_4_lut_LC_11_23_3.LUT_INIT=16'b1110110011001100;
    LogicCell40 i10150_4_lut_LC_11_23_3 (
            .in0(N__42118),
            .in1(N__42377),
            .in2(N__41979),
            .in3(N__41976),
            .lcout(n861),
            .ltout(n861_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i570_3_lut_LC_11_23_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i570_3_lut_LC_11_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i570_3_lut_LC_11_23_4.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i570_3_lut_LC_11_23_4 (
            .in0(_gnd_net_),
            .in1(N__42155),
            .in2(N__41970),
            .in3(N__42135),
            .lcout(n930),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_83_LC_11_23_6.C_ON=1'b0;
    defparam i1_4_lut_adj_83_LC_11_23_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_83_LC_11_23_6.LUT_INIT=16'b1111111011001100;
    LogicCell40 i1_4_lut_adj_83_LC_11_23_6 (
            .in0(N__42347),
            .in1(N__42317),
            .in2(N__42281),
            .in3(N__42263),
            .lcout(n5_adj_682),
            .ltout(n5_adj_682_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_84_LC_11_23_7.C_ON=1'b0;
    defparam i1_3_lut_adj_84_LC_11_23_7.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_84_LC_11_23_7.LUT_INIT=16'b1100000000000000;
    LogicCell40 i1_3_lut_adj_84_LC_11_23_7 (
            .in0(_gnd_net_),
            .in1(N__42219),
            .in2(N__42198),
            .in3(N__42427),
            .lcout(n13653),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_2_lut_LC_11_24_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_565_2_lut_LC_11_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_2_lut_LC_11_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_565_2_lut_LC_11_24_0 (
            .in0(_gnd_net_),
            .in1(N__43874),
            .in2(_gnd_net_),
            .in3(N__42168),
            .lcout(n901),
            .ltout(),
            .carryin(bfn_11_24_0_),
            .carryout(n12501),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_3_lut_LC_11_24_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_565_3_lut_LC_11_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_3_lut_LC_11_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_565_3_lut_LC_11_24_1 (
            .in0(_gnd_net_),
            .in1(N__53813),
            .in2(N__43592),
            .in3(N__42165),
            .lcout(n900),
            .ltout(),
            .carryin(n12501),
            .carryout(n12502),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_4_lut_LC_11_24_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_565_4_lut_LC_11_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_4_lut_LC_11_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_565_4_lut_LC_11_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43620),
            .in3(N__42162),
            .lcout(n899),
            .ltout(),
            .carryin(n12502),
            .carryout(n12503),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_5_lut_LC_11_24_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_565_5_lut_LC_11_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_5_lut_LC_11_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_565_5_lut_LC_11_24_3 (
            .in0(_gnd_net_),
            .in1(N__53814),
            .in2(N__42159),
            .in3(N__42129),
            .lcout(n898),
            .ltout(),
            .carryin(n12503),
            .carryout(n12504),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_6_lut_LC_11_24_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_565_6_lut_LC_11_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_6_lut_LC_11_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_565_6_lut_LC_11_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42126),
            .in3(N__42093),
            .lcout(n897),
            .ltout(),
            .carryin(n12504),
            .carryout(n12505),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_7_lut_LC_11_24_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_565_7_lut_LC_11_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_7_lut_LC_11_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_565_7_lut_LC_11_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__44063),
            .in3(N__42090),
            .lcout(n896),
            .ltout(),
            .carryin(n12505),
            .carryout(n12506),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_565_8_lut_LC_11_24_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_565_8_lut_LC_11_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_565_8_lut_LC_11_24_6.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_565_8_lut_LC_11_24_6 (
            .in0(N__53815),
            .in1(N__44093),
            .in2(N__42381),
            .in3(N__42432),
            .lcout(n927),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i500_4_lut_LC_11_24_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i500_4_lut_LC_11_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i500_4_lut_LC_11_24_7.LUT_INIT=16'b1010100000001000;
    LogicCell40 encoder0_position_31__I_0_i500_4_lut_LC_11_24_7 (
            .in0(N__42429),
            .in1(N__49560),
            .in2(N__42399),
            .in3(N__42390),
            .lcout(n828),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i4_1_lut_LC_11_25_0.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i4_1_lut_LC_11_25_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i4_1_lut_LC_11_25_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i4_1_lut_LC_11_25_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42366),
            .lcout(n22_adj_554),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i7_1_lut_LC_11_25_1.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i7_1_lut_LC_11_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i7_1_lut_LC_11_25_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i7_1_lut_LC_11_25_1 (
            .in0(N__42357),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n19_adj_557),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i4_1_lut_LC_11_25_2.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i4_1_lut_LC_11_25_2.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i4_1_lut_LC_11_25_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i4_1_lut_LC_11_25_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46142),
            .lcout(n22_adj_594),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i8_1_lut_LC_11_25_3.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i8_1_lut_LC_11_25_3.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i8_1_lut_LC_11_25_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i8_1_lut_LC_11_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44333),
            .lcout(n18_adj_590),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i1_1_lut_LC_11_25_4.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i1_1_lut_LC_11_25_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i1_1_lut_LC_11_25_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i1_1_lut_LC_11_25_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44501),
            .lcout(n25_adj_597),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i6_1_lut_LC_11_25_5.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i6_1_lut_LC_11_25_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i6_1_lut_LC_11_25_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i6_1_lut_LC_11_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43958),
            .lcout(n20_adj_592),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i5_1_lut_LC_11_25_6.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i5_1_lut_LC_11_25_6.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i5_1_lut_LC_11_25_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i5_1_lut_LC_11_25_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43991),
            .lcout(n21_adj_593),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i3_1_lut_LC_11_25_7.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i3_1_lut_LC_11_25_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i3_1_lut_LC_11_25_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i3_1_lut_LC_11_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42513),
            .lcout(n23_adj_553),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_2_lut_LC_11_26_0.C_ON=1'b1;
    defparam unary_minus_13_add_3_2_lut_LC_11_26_0.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_2_lut_LC_11_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_2_lut_LC_11_26_0 (
            .in0(_gnd_net_),
            .in1(N__42504),
            .in2(_gnd_net_),
            .in3(N__42498),
            .lcout(pwm_setpoint_23_N_171_0),
            .ltout(),
            .carryin(bfn_11_26_0_),
            .carryout(n12426),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_3_lut_LC_11_26_1.C_ON=1'b1;
    defparam unary_minus_13_add_3_3_lut_LC_11_26_1.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_3_lut_LC_11_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_3_lut_LC_11_26_1 (
            .in0(_gnd_net_),
            .in1(N__47850),
            .in2(_gnd_net_),
            .in3(N__42495),
            .lcout(pwm_setpoint_23_N_171_1),
            .ltout(),
            .carryin(n12426),
            .carryout(n12427),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_4_lut_LC_11_26_2.C_ON=1'b1;
    defparam unary_minus_13_add_3_4_lut_LC_11_26_2.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_4_lut_LC_11_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_4_lut_LC_11_26_2 (
            .in0(_gnd_net_),
            .in1(N__46512),
            .in2(_gnd_net_),
            .in3(N__42492),
            .lcout(pwm_setpoint_23_N_171_2),
            .ltout(),
            .carryin(n12427),
            .carryout(n12428),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_5_lut_LC_11_26_3.C_ON=1'b1;
    defparam unary_minus_13_add_3_5_lut_LC_11_26_3.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_5_lut_LC_11_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_5_lut_LC_11_26_3 (
            .in0(_gnd_net_),
            .in1(N__42489),
            .in2(_gnd_net_),
            .in3(N__42483),
            .lcout(pwm_setpoint_23_N_171_3),
            .ltout(),
            .carryin(n12428),
            .carryout(n12429),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_6_lut_LC_11_26_4.C_ON=1'b1;
    defparam unary_minus_13_add_3_6_lut_LC_11_26_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_6_lut_LC_11_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_6_lut_LC_11_26_4 (
            .in0(_gnd_net_),
            .in1(N__42480),
            .in2(_gnd_net_),
            .in3(N__42468),
            .lcout(pwm_setpoint_23_N_171_4),
            .ltout(),
            .carryin(n12429),
            .carryout(n12430),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_7_lut_LC_11_26_5.C_ON=1'b1;
    defparam unary_minus_13_add_3_7_lut_LC_11_26_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_7_lut_LC_11_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_7_lut_LC_11_26_5 (
            .in0(_gnd_net_),
            .in1(N__42465),
            .in2(_gnd_net_),
            .in3(N__42453),
            .lcout(pwm_setpoint_23_N_171_5),
            .ltout(),
            .carryin(n12430),
            .carryout(n12431),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_8_lut_LC_11_26_6.C_ON=1'b1;
    defparam unary_minus_13_add_3_8_lut_LC_11_26_6.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_8_lut_LC_11_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_8_lut_LC_11_26_6 (
            .in0(_gnd_net_),
            .in1(N__47301),
            .in2(_gnd_net_),
            .in3(N__42450),
            .lcout(pwm_setpoint_23_N_171_6),
            .ltout(),
            .carryin(n12431),
            .carryout(n12432),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_9_lut_LC_11_26_7.C_ON=1'b1;
    defparam unary_minus_13_add_3_9_lut_LC_11_26_7.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_9_lut_LC_11_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_9_lut_LC_11_26_7 (
            .in0(_gnd_net_),
            .in1(N__42447),
            .in2(_gnd_net_),
            .in3(N__42435),
            .lcout(pwm_setpoint_23_N_171_7),
            .ltout(),
            .carryin(n12432),
            .carryout(n12433),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_10_lut_LC_11_27_0.C_ON=1'b1;
    defparam unary_minus_13_add_3_10_lut_LC_11_27_0.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_10_lut_LC_11_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_10_lut_LC_11_27_0 (
            .in0(_gnd_net_),
            .in1(N__42639),
            .in2(_gnd_net_),
            .in3(N__42621),
            .lcout(pwm_setpoint_23_N_171_8),
            .ltout(),
            .carryin(bfn_11_27_0_),
            .carryout(n12434),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_11_lut_LC_11_27_1.C_ON=1'b1;
    defparam unary_minus_13_add_3_11_lut_LC_11_27_1.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_11_lut_LC_11_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_11_lut_LC_11_27_1 (
            .in0(_gnd_net_),
            .in1(N__42618),
            .in2(_gnd_net_),
            .in3(N__42606),
            .lcout(pwm_setpoint_23_N_171_9),
            .ltout(),
            .carryin(n12434),
            .carryout(n12435),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_12_lut_LC_11_27_2.C_ON=1'b1;
    defparam unary_minus_13_add_3_12_lut_LC_11_27_2.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_12_lut_LC_11_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_12_lut_LC_11_27_2 (
            .in0(_gnd_net_),
            .in1(N__42603),
            .in2(_gnd_net_),
            .in3(N__42591),
            .lcout(pwm_setpoint_23_N_171_10),
            .ltout(),
            .carryin(n12435),
            .carryout(n12436),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_13_lut_LC_11_27_3.C_ON=1'b1;
    defparam unary_minus_13_add_3_13_lut_LC_11_27_3.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_13_lut_LC_11_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_13_lut_LC_11_27_3 (
            .in0(_gnd_net_),
            .in1(N__42588),
            .in2(_gnd_net_),
            .in3(N__42570),
            .lcout(pwm_setpoint_23_N_171_11),
            .ltout(),
            .carryin(n12436),
            .carryout(n12437),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_14_lut_LC_11_27_4.C_ON=1'b1;
    defparam unary_minus_13_add_3_14_lut_LC_11_27_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_14_lut_LC_11_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_14_lut_LC_11_27_4 (
            .in0(_gnd_net_),
            .in1(N__44937),
            .in2(_gnd_net_),
            .in3(N__42567),
            .lcout(pwm_setpoint_23_N_171_12),
            .ltout(),
            .carryin(n12437),
            .carryout(n12438),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_15_lut_LC_11_27_5.C_ON=1'b1;
    defparam unary_minus_13_add_3_15_lut_LC_11_27_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_15_lut_LC_11_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_15_lut_LC_11_27_5 (
            .in0(_gnd_net_),
            .in1(N__42564),
            .in2(_gnd_net_),
            .in3(N__42552),
            .lcout(pwm_setpoint_23_N_171_13),
            .ltout(),
            .carryin(n12438),
            .carryout(n12439),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_16_lut_LC_11_27_6.C_ON=1'b1;
    defparam unary_minus_13_add_3_16_lut_LC_11_27_6.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_16_lut_LC_11_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_16_lut_LC_11_27_6 (
            .in0(_gnd_net_),
            .in1(N__42549),
            .in2(_gnd_net_),
            .in3(N__42537),
            .lcout(pwm_setpoint_23_N_171_14),
            .ltout(),
            .carryin(n12439),
            .carryout(n12440),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_17_lut_LC_11_27_7.C_ON=1'b1;
    defparam unary_minus_13_add_3_17_lut_LC_11_27_7.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_17_lut_LC_11_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_17_lut_LC_11_27_7 (
            .in0(_gnd_net_),
            .in1(N__42534),
            .in2(_gnd_net_),
            .in3(N__42516),
            .lcout(pwm_setpoint_23_N_171_15),
            .ltout(),
            .carryin(n12440),
            .carryout(n12441),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_18_lut_LC_11_28_0.C_ON=1'b1;
    defparam unary_minus_13_add_3_18_lut_LC_11_28_0.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_18_lut_LC_11_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_18_lut_LC_11_28_0 (
            .in0(_gnd_net_),
            .in1(N__42684),
            .in2(_gnd_net_),
            .in3(N__42675),
            .lcout(pwm_setpoint_23_N_171_16),
            .ltout(),
            .carryin(bfn_11_28_0_),
            .carryout(n12442),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_19_lut_LC_11_28_1.C_ON=1'b1;
    defparam unary_minus_13_add_3_19_lut_LC_11_28_1.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_19_lut_LC_11_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_19_lut_LC_11_28_1 (
            .in0(_gnd_net_),
            .in1(N__44580),
            .in2(_gnd_net_),
            .in3(N__42672),
            .lcout(pwm_setpoint_23_N_171_17),
            .ltout(),
            .carryin(n12442),
            .carryout(n12443),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_20_lut_LC_11_28_2.C_ON=1'b1;
    defparam unary_minus_13_add_3_20_lut_LC_11_28_2.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_20_lut_LC_11_28_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_20_lut_LC_11_28_2 (
            .in0(_gnd_net_),
            .in1(N__44532),
            .in2(_gnd_net_),
            .in3(N__42657),
            .lcout(pwm_setpoint_23_N_171_18),
            .ltout(),
            .carryin(n12443),
            .carryout(n12444),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_21_lut_LC_11_28_3.C_ON=1'b1;
    defparam unary_minus_13_add_3_21_lut_LC_11_28_3.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_21_lut_LC_11_28_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_21_lut_LC_11_28_3 (
            .in0(_gnd_net_),
            .in1(N__46737),
            .in2(_gnd_net_),
            .in3(N__42654),
            .lcout(pwm_setpoint_23_N_171_19),
            .ltout(),
            .carryin(n12444),
            .carryout(n12445),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_22_lut_LC_11_28_4.C_ON=1'b1;
    defparam unary_minus_13_add_3_22_lut_LC_11_28_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_22_lut_LC_11_28_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_22_lut_LC_11_28_4 (
            .in0(_gnd_net_),
            .in1(N__44475),
            .in2(_gnd_net_),
            .in3(N__42651),
            .lcout(pwm_setpoint_23_N_171_20),
            .ltout(),
            .carryin(n12445),
            .carryout(n12446),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_23_lut_LC_11_28_5.C_ON=1'b1;
    defparam unary_minus_13_add_3_23_lut_LC_11_28_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_23_lut_LC_11_28_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_23_lut_LC_11_28_5 (
            .in0(_gnd_net_),
            .in1(N__44559),
            .in2(_gnd_net_),
            .in3(N__42648),
            .lcout(pwm_setpoint_23_N_171_21),
            .ltout(),
            .carryin(n12446),
            .carryout(n12447),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_add_3_24_lut_LC_11_28_6.C_ON=1'b1;
    defparam unary_minus_13_add_3_24_lut_LC_11_28_6.SEQ_MODE=4'b0000;
    defparam unary_minus_13_add_3_24_lut_LC_11_28_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 unary_minus_13_add_3_24_lut_LC_11_28_6 (
            .in0(_gnd_net_),
            .in1(N__44625),
            .in2(_gnd_net_),
            .in3(N__42645),
            .lcout(pwm_setpoint_23_N_171_22),
            .ltout(),
            .carryin(n12447),
            .carryout(n12448),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i23_LC_11_28_7.C_ON=1'b0;
    defparam pwm_setpoint_i23_LC_11_28_7.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i23_LC_11_28_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 pwm_setpoint_i23_LC_11_28_7 (
            .in0(_gnd_net_),
            .in1(N__47837),
            .in2(_gnd_net_),
            .in3(N__42642),
            .lcout(pwm_setpoint_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56225),
            .ce(),
            .sr(N__47838));
    defparam LessThan_299_i19_2_lut_LC_11_29_0.C_ON=1'b0;
    defparam LessThan_299_i19_2_lut_LC_11_29_0.SEQ_MODE=4'b0000;
    defparam LessThan_299_i19_2_lut_LC_11_29_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i19_2_lut_LC_11_29_0 (
            .in0(_gnd_net_),
            .in1(N__42703),
            .in2(_gnd_net_),
            .in3(N__48395),
            .lcout(n19_adj_666),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i16_3_lut_3_lut_LC_11_29_1.C_ON=1'b0;
    defparam LessThan_299_i16_3_lut_3_lut_LC_11_29_1.SEQ_MODE=4'b0000;
    defparam LessThan_299_i16_3_lut_3_lut_LC_11_29_1.LUT_INIT=16'b1011101100100010;
    LogicCell40 LessThan_299_i16_3_lut_3_lut_LC_11_29_1 (
            .in0(N__42704),
            .in1(N__48475),
            .in2(_gnd_net_),
            .in3(N__44878),
            .lcout(),
            .ltout(n16_adj_664_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i24_3_lut_LC_11_29_2.C_ON=1'b0;
    defparam LessThan_299_i24_3_lut_LC_11_29_2.SEQ_MODE=4'b0000;
    defparam LessThan_299_i24_3_lut_LC_11_29_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 LessThan_299_i24_3_lut_LC_11_29_2 (
            .in0(_gnd_net_),
            .in1(N__44715),
            .in2(N__42747),
            .in3(N__44677),
            .lcout(),
            .ltout(n24_adj_669_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12493_4_lut_LC_11_29_3.C_ON=1'b0;
    defparam i12493_4_lut_LC_11_29_3.SEQ_MODE=4'b0000;
    defparam i12493_4_lut_LC_11_29_3.LUT_INIT=16'b1111000111100000;
    LogicCell40 i12493_4_lut_LC_11_29_3 (
            .in0(N__44678),
            .in1(N__42729),
            .in2(N__42744),
            .in3(N__42741),
            .lcout(n15223),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12414_2_lut_4_lut_LC_11_29_4.C_ON=1'b0;
    defparam i12414_2_lut_4_lut_LC_11_29_4.SEQ_MODE=4'b0000;
    defparam i12414_2_lut_4_lut_LC_11_29_4.LUT_INIT=16'b0111101111011110;
    LogicCell40 i12414_2_lut_4_lut_LC_11_29_4 (
            .in0(N__44879),
            .in1(N__42705),
            .in2(N__48477),
            .in3(N__48396),
            .lcout(n15144),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i23_2_lut_LC_11_29_5.C_ON=1'b0;
    defparam LessThan_299_i23_2_lut_LC_11_29_5.SEQ_MODE=4'b0000;
    defparam LessThan_299_i23_2_lut_LC_11_29_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i23_2_lut_LC_11_29_5 (
            .in0(_gnd_net_),
            .in1(N__42929),
            .in2(_gnd_net_),
            .in3(N__48344),
            .lcout(n23_adj_668),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i21_LC_11_29_6.C_ON=1'b0;
    defparam pwm_setpoint_i21_LC_11_29_6.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i21_LC_11_29_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 pwm_setpoint_i21_LC_11_29_6 (
            .in0(N__42723),
            .in1(N__50892),
            .in2(_gnd_net_),
            .in3(N__44574),
            .lcout(pwm_setpoint_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56230),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i9_LC_11_29_7.C_ON=1'b0;
    defparam pwm_setpoint_i9_LC_11_29_7.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i9_LC_11_29_7.LUT_INIT=16'b1111010110100000;
    LogicCell40 pwm_setpoint_i9_LC_11_29_7 (
            .in0(N__50893),
            .in1(_gnd_net_),
            .in2(N__42717),
            .in3(N__44271),
            .lcout(pwm_setpoint_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56230),
            .ce(),
            .sr(_gnd_net_));
    defparam i12448_4_lut_LC_11_30_0.C_ON=1'b0;
    defparam i12448_4_lut_LC_11_30_0.SEQ_MODE=4'b0000;
    defparam i12448_4_lut_LC_11_30_0.LUT_INIT=16'b1111111111001101;
    LogicCell40 i12448_4_lut_LC_11_30_0 (
            .in0(N__42815),
            .in1(N__46809),
            .in2(N__46239),
            .in3(N__44747),
            .lcout(n15178),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i14_LC_11_30_1.C_ON=1'b0;
    defparam pwm_setpoint_i14_LC_11_30_1.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i14_LC_11_30_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 pwm_setpoint_i14_LC_11_30_1 (
            .in0(N__50894),
            .in1(N__44120),
            .in2(_gnd_net_),
            .in3(N__42693),
            .lcout(pwm_setpoint_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56237),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i22_LC_11_30_2.C_ON=1'b0;
    defparam pwm_setpoint_i22_LC_11_30_2.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i22_LC_11_30_2.LUT_INIT=16'b1110111000100010;
    LogicCell40 pwm_setpoint_i22_LC_11_30_2 (
            .in0(N__44643),
            .in1(N__50895),
            .in2(_gnd_net_),
            .in3(N__42825),
            .lcout(pwm_setpoint_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56237),
            .ce(),
            .sr(_gnd_net_));
    defparam i12380_4_lut_LC_11_30_3.C_ON=1'b0;
    defparam i12380_4_lut_LC_11_30_3.SEQ_MODE=4'b0000;
    defparam i12380_4_lut_LC_11_30_3.LUT_INIT=16'b1010101010101011;
    LogicCell40 i12380_4_lut_LC_11_30_3 (
            .in0(N__47144),
            .in1(N__42780),
            .in2(N__42789),
            .in3(N__42816),
            .lcout(n15110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i15_2_lut_LC_11_30_4.C_ON=1'b0;
    defparam LessThan_299_i15_2_lut_LC_11_30_4.SEQ_MODE=4'b0000;
    defparam LessThan_299_i15_2_lut_LC_11_30_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i15_2_lut_LC_11_30_4 (
            .in0(_gnd_net_),
            .in1(N__48017),
            .in2(_gnd_net_),
            .in3(N__42965),
            .lcout(n15_adj_663),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i17_2_lut_LC_11_30_5.C_ON=1'b0;
    defparam LessThan_299_i17_2_lut_LC_11_30_5.SEQ_MODE=4'b0000;
    defparam LessThan_299_i17_2_lut_LC_11_30_5.LUT_INIT=16'b0101010110101010;
    LogicCell40 LessThan_299_i17_2_lut_LC_11_30_5 (
            .in0(N__42804),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47978),
            .lcout(n17_adj_665),
            .ltout(n17_adj_665_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12444_4_lut_LC_11_30_6.C_ON=1'b0;
    defparam i12444_4_lut_LC_11_30_6.SEQ_MODE=4'b0000;
    defparam i12444_4_lut_LC_11_30_6.LUT_INIT=16'b1111101011111011;
    LogicCell40 i12444_4_lut_LC_11_30_6 (
            .in0(N__42779),
            .in1(N__42771),
            .in2(N__42765),
            .in3(N__44733),
            .lcout(n15174),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i33_2_lut_LC_11_31_0.C_ON=1'b0;
    defparam LessThan_299_i33_2_lut_LC_11_31_0.SEQ_MODE=4'b0000;
    defparam LessThan_299_i33_2_lut_LC_11_31_0.LUT_INIT=16'b0101010110101010;
    LogicCell40 LessThan_299_i33_2_lut_LC_11_31_0 (
            .in0(N__42981),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48213),
            .lcout(n33_adj_675),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12367_2_lut_4_lut_LC_11_31_1.C_ON=1'b0;
    defparam i12367_2_lut_4_lut_LC_11_31_1.SEQ_MODE=4'b0000;
    defparam i12367_2_lut_4_lut_LC_11_31_1.LUT_INIT=16'b0110111111110110;
    LogicCell40 i12367_2_lut_4_lut_LC_11_31_1 (
            .in0(N__48212),
            .in1(N__42980),
            .in2(N__42969),
            .in3(N__48018),
            .lcout(n15097),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12435_3_lut_LC_11_31_2.C_ON=1'b0;
    defparam i12435_3_lut_LC_11_31_2.SEQ_MODE=4'b0000;
    defparam i12435_3_lut_LC_11_31_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 i12435_3_lut_LC_11_31_2 (
            .in0(N__44808),
            .in1(N__44820),
            .in2(_gnd_net_),
            .in3(N__42906),
            .lcout(n15165),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i16_LC_11_31_3.C_ON=1'b0;
    defparam pwm_setpoint_i16_LC_11_31_3.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i16_LC_11_31_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 pwm_setpoint_i16_LC_11_31_3 (
            .in0(N__42762),
            .in1(N__50900),
            .in2(_gnd_net_),
            .in3(N__44454),
            .lcout(pwm_setpoint_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56243),
            .ce(),
            .sr(_gnd_net_));
    defparam i12507_4_lut_LC_11_31_5.C_ON=1'b0;
    defparam i12507_4_lut_LC_11_31_5.SEQ_MODE=4'b0000;
    defparam i12507_4_lut_LC_11_31_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12507_4_lut_LC_11_31_5 (
            .in0(N__42753),
            .in1(N__44789),
            .in2(N__47145),
            .in3(N__44807),
            .lcout(n15237),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i17_LC_11_31_6.C_ON=1'b0;
    defparam pwm_setpoint_i17_LC_11_31_6.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i17_LC_11_31_6.LUT_INIT=16'b1110111001000100;
    LogicCell40 pwm_setpoint_i17_LC_11_31_6 (
            .in0(N__50901),
            .in1(N__44598),
            .in2(_gnd_net_),
            .in3(N__42990),
            .lcout(pwm_setpoint_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56243),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i12_3_lut_3_lut_LC_11_31_7.C_ON=1'b0;
    defparam LessThan_299_i12_3_lut_3_lut_LC_11_31_7.SEQ_MODE=4'b0000;
    defparam LessThan_299_i12_3_lut_3_lut_LC_11_31_7.LUT_INIT=16'b1101110101000100;
    LogicCell40 LessThan_299_i12_3_lut_3_lut_LC_11_31_7 (
            .in0(N__48211),
            .in1(N__42979),
            .in2(_gnd_net_),
            .in3(N__42964),
            .lcout(n12_adj_661),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i10_LC_11_32_1.C_ON=1'b0;
    defparam pwm_setpoint_i10_LC_11_32_1.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i10_LC_11_32_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 pwm_setpoint_i10_LC_11_32_1 (
            .in0(N__50910),
            .in1(N__42939),
            .in2(_gnd_net_),
            .in3(N__44235),
            .lcout(pwm_setpoint_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56249),
            .ce(),
            .sr(_gnd_net_));
    defparam i12474_3_lut_LC_11_32_3.C_ON=1'b0;
    defparam i12474_3_lut_LC_11_32_3.SEQ_MODE=4'b0000;
    defparam i12474_3_lut_LC_11_32_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 i12474_3_lut_LC_11_32_3 (
            .in0(N__47094),
            .in1(N__42930),
            .in2(_gnd_net_),
            .in3(N__44790),
            .lcout(n15204),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i35_2_lut_LC_11_32_5.C_ON=1'b0;
    defparam LessThan_299_i35_2_lut_LC_11_32_5.SEQ_MODE=4'b0000;
    defparam LessThan_299_i35_2_lut_LC_11_32_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i35_2_lut_LC_11_32_5 (
            .in0(_gnd_net_),
            .in1(N__42896),
            .in2(_gnd_net_),
            .in3(N__48582),
            .lcout(n35),
            .ltout(n35_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i30_3_lut_LC_11_32_6.C_ON=1'b0;
    defparam LessThan_299_i30_3_lut_LC_11_32_6.SEQ_MODE=4'b0000;
    defparam LessThan_299_i30_3_lut_LC_11_32_6.LUT_INIT=16'b1010111110100000;
    LogicCell40 LessThan_299_i30_3_lut_LC_11_32_6 (
            .in0(N__42897),
            .in1(_gnd_net_),
            .in2(N__42888),
            .in3(N__42885),
            .lcout(n30_adj_673),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1177_3_lut_LC_12_17_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1177_3_lut_LC_12_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1177_3_lut_LC_12_17_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1177_3_lut_LC_12_17_0 (
            .in0(_gnd_net_),
            .in1(N__43553),
            .in2(N__43539),
            .in3(N__45457),
            .lcout(n1825),
            .ltout(n1825_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_136_LC_12_17_1.C_ON=1'b0;
    defparam i1_4_lut_adj_136_LC_12_17_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_136_LC_12_17_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_136_LC_12_17_1 (
            .in0(N__43075),
            .in1(N__42841),
            .in2(N__42861),
            .in3(N__43162),
            .lcout(n14520),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1180_3_lut_LC_12_17_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1180_3_lut_LC_12_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1180_3_lut_LC_12_17_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1180_3_lut_LC_12_17_2 (
            .in0(_gnd_net_),
            .in1(N__43233),
            .in2(N__45681),
            .in3(N__45456),
            .lcout(n1828),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1182_3_lut_LC_12_17_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1182_3_lut_LC_12_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1182_3_lut_LC_12_17_3.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i1182_3_lut_LC_12_17_3 (
            .in0(N__43272),
            .in1(_gnd_net_),
            .in2(N__45486),
            .in3(N__43254),
            .lcout(n1830),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12904_4_lut_LC_12_17_4.C_ON=1'b0;
    defparam i12904_4_lut_LC_12_17_4.SEQ_MODE=4'b0000;
    defparam i12904_4_lut_LC_12_17_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12904_4_lut_LC_12_17_4 (
            .in0(N__43418),
            .in1(N__43390),
            .in2(N__45341),
            .in3(N__42996),
            .lcout(n1752),
            .ltout(n1752_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12480_3_lut_LC_12_17_5.C_ON=1'b0;
    defparam i12480_3_lut_LC_12_17_5.SEQ_MODE=4'b0000;
    defparam i12480_3_lut_LC_12_17_5.LUT_INIT=16'b1100111111000000;
    LogicCell40 i12480_3_lut_LC_12_17_5 (
            .in0(_gnd_net_),
            .in1(N__45314),
            .in2(N__43086),
            .in3(N__43206),
            .lcout(n1826),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1176_3_lut_LC_12_17_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1176_3_lut_LC_12_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1176_3_lut_LC_12_17_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1176_3_lut_LC_12_17_6 (
            .in0(_gnd_net_),
            .in1(N__43521),
            .in2(N__45210),
            .in3(N__45461),
            .lcout(n1824),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1175_3_lut_LC_12_17_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1175_3_lut_LC_12_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1175_3_lut_LC_12_17_7.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1175_3_lut_LC_12_17_7 (
            .in0(_gnd_net_),
            .in1(N__45245),
            .in2(N__45485),
            .in3(N__43506),
            .lcout(n1823),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12478_3_lut_LC_12_18_1.C_ON=1'b0;
    defparam i12478_3_lut_LC_12_18_1.SEQ_MODE=4'b0000;
    defparam i12478_3_lut_LC_12_18_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 i12478_3_lut_LC_12_18_1 (
            .in0(_gnd_net_),
            .in1(N__45135),
            .in2(N__47211),
            .in3(N__45608),
            .lcout(n1726),
            .ltout(n1726_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_132_LC_12_18_2.C_ON=1'b0;
    defparam i1_3_lut_adj_132_LC_12_18_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_132_LC_12_18_2.LUT_INIT=16'b1111111111111010;
    LogicCell40 i1_3_lut_adj_132_LC_12_18_2 (
            .in0(N__45277),
            .in1(_gnd_net_),
            .in2(N__43005),
            .in3(N__45310),
            .lcout(),
            .ltout(n14244_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_133_LC_12_18_3.C_ON=1'b0;
    defparam i1_4_lut_adj_133_LC_12_18_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_133_LC_12_18_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_133_LC_12_18_3 (
            .in0(N__45235),
            .in1(N__45196),
            .in2(N__43002),
            .in3(N__43483),
            .lcout(),
            .ltout(n14250_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_135_LC_12_18_4.C_ON=1'b0;
    defparam i1_4_lut_adj_135_LC_12_18_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_135_LC_12_18_4.LUT_INIT=16'b1111111011111010;
    LogicCell40 i1_4_lut_adj_135_LC_12_18_4 (
            .in0(N__43448),
            .in1(N__43353),
            .in2(N__42999),
            .in3(N__45654),
            .lcout(n14254),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1105_3_lut_LC_12_18_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1105_3_lut_LC_12_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1105_3_lut_LC_12_18_5.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1105_3_lut_LC_12_18_5 (
            .in0(_gnd_net_),
            .in1(N__47181),
            .in2(N__45099),
            .in3(N__45609),
            .lcout(n1721),
            .ltout(n1721_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1172_3_lut_LC_12_18_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1172_3_lut_LC_12_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1172_3_lut_LC_12_18_6.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1172_3_lut_LC_12_18_6 (
            .in0(N__45455),
            .in1(_gnd_net_),
            .in2(N__43197),
            .in3(N__43407),
            .lcout(n1820),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1179_3_lut_LC_12_18_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1179_3_lut_LC_12_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1179_3_lut_LC_12_18_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1179_3_lut_LC_12_18_7 (
            .in0(_gnd_net_),
            .in1(N__45278),
            .in2(N__43221),
            .in3(N__45454),
            .lcout(n1827),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1104_3_lut_LC_12_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1104_3_lut_LC_12_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1104_3_lut_LC_12_19_1.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1104_3_lut_LC_12_19_1 (
            .in0(N__45087),
            .in1(_gnd_net_),
            .in2(N__45372),
            .in3(N__45604),
            .lcout(n1720),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1107_3_lut_LC_12_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1107_3_lut_LC_12_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1107_3_lut_LC_12_19_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1107_3_lut_LC_12_19_2 (
            .in0(N__45602),
            .in1(_gnd_net_),
            .in2(N__47283),
            .in3(N__45120),
            .lcout(n1723),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1106_3_lut_LC_12_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1106_3_lut_LC_12_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1106_3_lut_LC_12_19_3.LUT_INIT=16'b1111110000110000;
    LogicCell40 encoder0_position_31__I_0_i1106_3_lut_LC_12_19_3 (
            .in0(_gnd_net_),
            .in1(N__45603),
            .in2(N__45111),
            .in3(N__47253),
            .lcout(n1722),
            .ltout(n1722_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1173_3_lut_LC_12_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1173_3_lut_LC_12_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1173_3_lut_LC_12_19_4.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i1173_3_lut_LC_12_19_4 (
            .in0(N__45484),
            .in1(_gnd_net_),
            .in2(N__43146),
            .in3(N__43437),
            .lcout(n1821),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1116_3_lut_LC_12_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1116_3_lut_LC_12_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1116_3_lut_LC_12_19_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1116_3_lut_LC_12_19_5 (
            .in0(_gnd_net_),
            .in1(N__44985),
            .in2(N__48756),
            .in3(N__45598),
            .lcout(n1732),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1115_3_lut_LC_12_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1115_3_lut_LC_12_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1115_3_lut_LC_12_19_6.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i1115_3_lut_LC_12_19_6 (
            .in0(N__44973),
            .in1(_gnd_net_),
            .in2(N__45616),
            .in3(N__48810),
            .lcout(n1731),
            .ltout(n1731_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10014_4_lut_LC_12_19_7.C_ON=1'b0;
    defparam i10014_4_lut_LC_12_19_7.SEQ_MODE=4'b0000;
    defparam i10014_4_lut_LC_12_19_7.LUT_INIT=16'b1111110011111000;
    LogicCell40 i10014_4_lut_LC_12_19_7 (
            .in0(N__43687),
            .in1(N__43303),
            .in2(N__43356),
            .in3(N__45526),
            .lcout(n11991),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_2_lut_LC_12_20_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_2_lut_LC_12_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_2_lut_LC_12_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_2_lut_LC_12_20_0 (
            .in0(_gnd_net_),
            .in1(N__43688),
            .in2(_gnd_net_),
            .in3(N__43335),
            .lcout(n1801),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(n12591),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_3_lut_LC_12_20_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_3_lut_LC_12_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_3_lut_LC_12_20_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_3_lut_LC_12_20_1 (
            .in0(_gnd_net_),
            .in1(N__54881),
            .in2(N__45533),
            .in3(N__43320),
            .lcout(n1800),
            .ltout(),
            .carryin(n12591),
            .carryout(n12592),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_4_lut_LC_12_20_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_4_lut_LC_12_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_4_lut_LC_12_20_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_4_lut_LC_12_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43310),
            .in3(N__43275),
            .lcout(n1799),
            .ltout(),
            .carryin(n12592),
            .carryout(n12593),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_5_lut_LC_12_20_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_5_lut_LC_12_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_5_lut_LC_12_20_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_5_lut_LC_12_20_3 (
            .in0(_gnd_net_),
            .in1(N__54882),
            .in2(N__43271),
            .in3(N__43245),
            .lcout(n1798),
            .ltout(),
            .carryin(n12593),
            .carryout(n12594),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_6_lut_LC_12_20_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_6_lut_LC_12_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_6_lut_LC_12_20_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_6_lut_LC_12_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45701),
            .in3(N__43236),
            .lcout(n1797),
            .ltout(),
            .carryin(n12594),
            .carryout(n12595),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_7_lut_LC_12_20_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_7_lut_LC_12_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_7_lut_LC_12_20_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_7_lut_LC_12_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45677),
            .in3(N__43224),
            .lcout(n1796),
            .ltout(),
            .carryin(n12595),
            .carryout(n12596),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_8_lut_LC_12_20_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_8_lut_LC_12_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_8_lut_LC_12_20_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_8_lut_LC_12_20_6 (
            .in0(_gnd_net_),
            .in1(N__55086),
            .in2(N__45282),
            .in3(N__43209),
            .lcout(n1795),
            .ltout(),
            .carryin(n12596),
            .carryout(n12597),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_9_lut_LC_12_20_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_9_lut_LC_12_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_9_lut_LC_12_20_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_9_lut_LC_12_20_7 (
            .in0(_gnd_net_),
            .in1(N__54883),
            .in2(N__45318),
            .in3(N__43563),
            .lcout(n1794),
            .ltout(),
            .carryin(n12597),
            .carryout(n12598),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_10_lut_LC_12_21_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_10_lut_LC_12_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_10_lut_LC_12_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_10_lut_LC_12_21_0 (
            .in0(_gnd_net_),
            .in1(N__54586),
            .in2(N__43560),
            .in3(N__43524),
            .lcout(n1793),
            .ltout(),
            .carryin(bfn_12_21_0_),
            .carryout(n12599),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_11_lut_LC_12_21_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_11_lut_LC_12_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_11_lut_LC_12_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_11_lut_LC_12_21_1 (
            .in0(_gnd_net_),
            .in1(N__54590),
            .in2(N__45209),
            .in3(N__43509),
            .lcout(n1792),
            .ltout(),
            .carryin(n12599),
            .carryout(n12600),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_12_lut_LC_12_21_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_12_lut_LC_12_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_12_lut_LC_12_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_12_lut_LC_12_21_2 (
            .in0(_gnd_net_),
            .in1(N__54587),
            .in2(N__45246),
            .in3(N__43494),
            .lcout(n1791),
            .ltout(),
            .carryin(n12600),
            .carryout(n12601),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_13_lut_LC_12_21_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_13_lut_LC_12_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_13_lut_LC_12_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_13_lut_LC_12_21_3 (
            .in0(_gnd_net_),
            .in1(N__54591),
            .in2(N__43491),
            .in3(N__43458),
            .lcout(n1790),
            .ltout(),
            .carryin(n12601),
            .carryout(n12602),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_14_lut_LC_12_21_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_14_lut_LC_12_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_14_lut_LC_12_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_14_lut_LC_12_21_4 (
            .in0(_gnd_net_),
            .in1(N__54588),
            .in2(N__43455),
            .in3(N__43428),
            .lcout(n1789),
            .ltout(),
            .carryin(n12602),
            .carryout(n12603),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_15_lut_LC_12_21_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_15_lut_LC_12_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_15_lut_LC_12_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_15_lut_LC_12_21_5 (
            .in0(_gnd_net_),
            .in1(N__54592),
            .in2(N__43425),
            .in3(N__43398),
            .lcout(n1788),
            .ltout(),
            .carryin(n12603),
            .carryout(n12604),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_16_lut_LC_12_21_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1168_16_lut_LC_12_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_16_lut_LC_12_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1168_16_lut_LC_12_21_6 (
            .in0(_gnd_net_),
            .in1(N__43391),
            .in2(N__54880),
            .in3(N__43362),
            .lcout(n1787),
            .ltout(),
            .carryin(n12604),
            .carryout(n12605),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1168_17_lut_LC_12_21_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1168_17_lut_LC_12_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1168_17_lut_LC_12_21_7.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1168_17_lut_LC_12_21_7 (
            .in0(N__54589),
            .in1(N__45345),
            .in2(N__45389),
            .in3(N__43359),
            .lcout(n1818),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut_LC_12_22_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut_LC_12_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut_LC_12_22_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut_LC_12_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43838),
            .lcout(n10_adj_628),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i17_3_lut_LC_12_22_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i17_3_lut_LC_12_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i17_3_lut_LC_12_22_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i17_3_lut_LC_12_22_5 (
            .in0(N__49611),
            .in1(N__43704),
            .in2(_gnd_net_),
            .in3(N__45759),
            .lcout(n303),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i19_3_lut_LC_12_22_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i19_3_lut_LC_12_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i19_3_lut_LC_12_22_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i19_3_lut_LC_12_22_6 (
            .in0(N__43668),
            .in1(N__49610),
            .in2(_gnd_net_),
            .in3(N__43655),
            .lcout(n301),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i571_3_lut_LC_12_23_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i571_3_lut_LC_12_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i571_3_lut_LC_12_23_0.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i571_3_lut_LC_12_23_0 (
            .in0(_gnd_net_),
            .in1(N__43626),
            .in2(N__43619),
            .in3(N__44090),
            .lcout(n931),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i636_3_lut_LC_12_23_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i636_3_lut_LC_12_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i636_3_lut_LC_12_23_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i636_3_lut_LC_12_23_1 (
            .in0(_gnd_net_),
            .in1(N__46064),
            .in2(N__46013),
            .in3(N__46050),
            .lcout(n1028),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i572_3_lut_LC_12_23_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i572_3_lut_LC_12_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i572_3_lut_LC_12_23_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i572_3_lut_LC_12_23_2 (
            .in0(_gnd_net_),
            .in1(N__43599),
            .in2(N__43593),
            .in3(N__44092),
            .lcout(n932),
            .ltout(n932_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i639_3_lut_LC_12_23_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i639_3_lut_LC_12_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i639_3_lut_LC_12_23_3.LUT_INIT=16'b1111101001010000;
    LogicCell40 encoder0_position_31__I_0_i639_3_lut_LC_12_23_3 (
            .in0(N__46004),
            .in1(_gnd_net_),
            .in2(N__43566),
            .in3(N__45864),
            .lcout(n1031),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i641_3_lut_LC_12_23_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i641_3_lut_LC_12_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i641_3_lut_LC_12_23_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i641_3_lut_LC_12_23_4 (
            .in0(N__45924),
            .in1(N__45912),
            .in2(_gnd_net_),
            .in3(N__46002),
            .lcout(n1033),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i26_3_lut_LC_12_23_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i26_3_lut_LC_12_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i26_3_lut_LC_12_23_5.LUT_INIT=16'b1111110000110000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i26_3_lut_LC_12_23_5 (
            .in0(_gnd_net_),
            .in1(N__49599),
            .in2(N__43920),
            .in3(N__43887),
            .lcout(n41),
            .ltout(n41_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i573_3_lut_LC_12_23_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i573_3_lut_LC_12_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i573_3_lut_LC_12_23_6.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i573_3_lut_LC_12_23_6 (
            .in0(N__43863),
            .in1(_gnd_net_),
            .in2(N__43857),
            .in3(N__44091),
            .lcout(n933),
            .ltout(n933_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i640_3_lut_LC_12_23_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i640_3_lut_LC_12_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i640_3_lut_LC_12_23_7.LUT_INIT=16'b1111101001010000;
    LogicCell40 encoder0_position_31__I_0_i640_3_lut_LC_12_23_7 (
            .in0(N__46003),
            .in1(_gnd_net_),
            .in2(N__43854),
            .in3(N__45888),
            .lcout(n1032),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i635_rep_47_3_lut_LC_12_24_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i635_rep_47_3_lut_LC_12_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i635_rep_47_3_lut_LC_12_24_0.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i635_rep_47_3_lut_LC_12_24_0 (
            .in0(_gnd_net_),
            .in1(N__46037),
            .in2(N__46014),
            .in3(N__46023),
            .lcout(n1027),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i24_3_lut_LC_12_24_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i24_3_lut_LC_12_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i24_3_lut_LC_12_24_1.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i24_3_lut_LC_12_24_1 (
            .in0(_gnd_net_),
            .in1(N__49602),
            .in2(N__43851),
            .in3(N__43839),
            .lcout(n296),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i25_3_lut_LC_12_24_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i25_3_lut_LC_12_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i25_3_lut_LC_12_24_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 encoder0_position_31__I_0_mux_3_i25_3_lut_LC_12_24_3 (
            .in0(N__43808),
            .in1(N__49601),
            .in2(_gnd_net_),
            .in3(N__43779),
            .lcout(n295),
            .ltout(n295_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9978_4_lut_LC_12_24_4.C_ON=1'b0;
    defparam i9978_4_lut_LC_12_24_4.SEQ_MODE=4'b0000;
    defparam i9978_4_lut_LC_12_24_4.LUT_INIT=16'b1111111010101010;
    LogicCell40 i9978_4_lut_LC_12_24_4 (
            .in0(N__45850),
            .in1(N__45899),
            .in2(N__43764),
            .in3(N__45875),
            .lcout(),
            .ltout(n11955_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_86_LC_12_24_5.C_ON=1'b0;
    defparam i1_4_lut_adj_86_LC_12_24_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_86_LC_12_24_5.LUT_INIT=16'b1111111011101110;
    LogicCell40 i1_4_lut_adj_86_LC_12_24_5 (
            .in0(N__46036),
            .in1(N__45968),
            .in2(N__43761),
            .in3(N__43758),
            .lcout(n960),
            .ltout(n960_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i637_3_lut_LC_12_24_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i637_3_lut_LC_12_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i637_3_lut_LC_12_24_6.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i637_3_lut_LC_12_24_6 (
            .in0(N__46100),
            .in1(_gnd_net_),
            .in2(N__43752),
            .in3(N__46080),
            .lcout(n1029),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i568_3_lut_LC_12_24_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i568_3_lut_LC_12_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i568_3_lut_LC_12_24_7.LUT_INIT=16'b1111110000110000;
    LogicCell40 encoder0_position_31__I_0_i568_3_lut_LC_12_24_7 (
            .in0(_gnd_net_),
            .in1(N__44094),
            .in2(N__44064),
            .in3(N__44046),
            .lcout(n928),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i0_LC_12_25_0.C_ON=1'b1;
    defparam duty_i0_LC_12_25_0.SEQ_MODE=4'b1000;
    defparam duty_i0_LC_12_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i0_LC_12_25_0 (
            .in0(_gnd_net_),
            .in1(N__45945),
            .in2(N__49770),
            .in3(N__44040),
            .lcout(duty_0),
            .ltout(),
            .carryin(bfn_12_25_0_),
            .carryout(n12473),
            .clk(N__56218),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i1_LC_12_25_1.C_ON=1'b1;
    defparam duty_i1_LC_12_25_1.SEQ_MODE=4'b1000;
    defparam duty_i1_LC_12_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i1_LC_12_25_1 (
            .in0(_gnd_net_),
            .in1(N__44037),
            .in2(N__49740),
            .in3(N__44028),
            .lcout(duty_1),
            .ltout(),
            .carryin(n12473),
            .carryout(n12474),
            .clk(N__56218),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i2_LC_12_25_2.C_ON=1'b1;
    defparam duty_i2_LC_12_25_2.SEQ_MODE=4'b1000;
    defparam duty_i2_LC_12_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i2_LC_12_25_2 (
            .in0(_gnd_net_),
            .in1(N__44025),
            .in2(N__49704),
            .in3(N__44019),
            .lcout(duty_2),
            .ltout(),
            .carryin(n12474),
            .carryout(n12475),
            .clk(N__56218),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i3_LC_12_25_3.C_ON=1'b1;
    defparam duty_i3_LC_12_25_3.SEQ_MODE=4'b1000;
    defparam duty_i3_LC_12_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i3_LC_12_25_3 (
            .in0(_gnd_net_),
            .in1(N__44016),
            .in2(N__50352),
            .in3(N__44010),
            .lcout(duty_3),
            .ltout(),
            .carryin(n12475),
            .carryout(n12476),
            .clk(N__56218),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i4_LC_12_25_4.C_ON=1'b1;
    defparam duty_i4_LC_12_25_4.SEQ_MODE=4'b1000;
    defparam duty_i4_LC_12_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i4_LC_12_25_4 (
            .in0(_gnd_net_),
            .in1(N__44007),
            .in2(N__50319),
            .in3(N__43980),
            .lcout(duty_4),
            .ltout(),
            .carryin(n12476),
            .carryout(n12477),
            .clk(N__56218),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i5_LC_12_25_5.C_ON=1'b1;
    defparam duty_i5_LC_12_25_5.SEQ_MODE=4'b1000;
    defparam duty_i5_LC_12_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i5_LC_12_25_5 (
            .in0(_gnd_net_),
            .in1(N__43977),
            .in2(N__50274),
            .in3(N__43947),
            .lcout(duty_5),
            .ltout(),
            .carryin(n12477),
            .carryout(n12478),
            .clk(N__56218),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i6_LC_12_25_6.C_ON=1'b1;
    defparam duty_i6_LC_12_25_6.SEQ_MODE=4'b1000;
    defparam duty_i6_LC_12_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i6_LC_12_25_6 (
            .in0(_gnd_net_),
            .in1(N__43944),
            .in2(N__50238),
            .in3(N__43938),
            .lcout(duty_6),
            .ltout(),
            .carryin(n12478),
            .carryout(n12479),
            .clk(N__56218),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i7_LC_12_25_7.C_ON=1'b1;
    defparam duty_i7_LC_12_25_7.SEQ_MODE=4'b1000;
    defparam duty_i7_LC_12_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i7_LC_12_25_7 (
            .in0(_gnd_net_),
            .in1(N__43935),
            .in2(N__50202),
            .in3(N__44322),
            .lcout(duty_7),
            .ltout(),
            .carryin(n12479),
            .carryout(n12480),
            .clk(N__56218),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i8_LC_12_26_0.C_ON=1'b1;
    defparam duty_i8_LC_12_26_0.SEQ_MODE=4'b1000;
    defparam duty_i8_LC_12_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i8_LC_12_26_0 (
            .in0(_gnd_net_),
            .in1(N__44319),
            .in2(N__50157),
            .in3(N__44283),
            .lcout(duty_8),
            .ltout(),
            .carryin(bfn_12_26_0_),
            .carryout(n12481),
            .clk(N__56221),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i9_LC_12_26_1.C_ON=1'b1;
    defparam duty_i9_LC_12_26_1.SEQ_MODE=4'b1000;
    defparam duty_i9_LC_12_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i9_LC_12_26_1 (
            .in0(_gnd_net_),
            .in1(N__44280),
            .in2(N__50118),
            .in3(N__44247),
            .lcout(duty_9),
            .ltout(),
            .carryin(n12481),
            .carryout(n12482),
            .clk(N__56221),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i10_LC_12_26_2.C_ON=1'b1;
    defparam duty_i10_LC_12_26_2.SEQ_MODE=4'b1000;
    defparam duty_i10_LC_12_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i10_LC_12_26_2 (
            .in0(_gnd_net_),
            .in1(N__44244),
            .in2(N__50076),
            .in3(N__44214),
            .lcout(duty_10),
            .ltout(),
            .carryin(n12482),
            .carryout(n12483),
            .clk(N__56221),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i11_LC_12_26_3.C_ON=1'b1;
    defparam duty_i11_LC_12_26_3.SEQ_MODE=4'b1000;
    defparam duty_i11_LC_12_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i11_LC_12_26_3 (
            .in0(_gnd_net_),
            .in1(N__44211),
            .in2(N__50709),
            .in3(N__44178),
            .lcout(duty_11),
            .ltout(),
            .carryin(n12483),
            .carryout(n12484),
            .clk(N__56221),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i12_LC_12_26_4.C_ON=1'b1;
    defparam duty_i12_LC_12_26_4.SEQ_MODE=4'b1000;
    defparam duty_i12_LC_12_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i12_LC_12_26_4 (
            .in0(_gnd_net_),
            .in1(N__50674),
            .in2(N__44175),
            .in3(N__44163),
            .lcout(duty_12),
            .ltout(),
            .carryin(n12484),
            .carryout(n12485),
            .clk(N__56221),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i13_LC_12_26_5.C_ON=1'b1;
    defparam duty_i13_LC_12_26_5.SEQ_MODE=4'b1000;
    defparam duty_i13_LC_12_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i13_LC_12_26_5 (
            .in0(_gnd_net_),
            .in1(N__44160),
            .in2(N__50637),
            .in3(N__44133),
            .lcout(duty_13),
            .ltout(),
            .carryin(n12485),
            .carryout(n12486),
            .clk(N__56221),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i14_LC_12_26_6.C_ON=1'b1;
    defparam duty_i14_LC_12_26_6.SEQ_MODE=4'b1000;
    defparam duty_i14_LC_12_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i14_LC_12_26_6 (
            .in0(_gnd_net_),
            .in1(N__44130),
            .in2(N__50598),
            .in3(N__44097),
            .lcout(duty_14),
            .ltout(),
            .carryin(n12486),
            .carryout(n12487),
            .clk(N__56221),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i15_LC_12_26_7.C_ON=1'b1;
    defparam duty_i15_LC_12_26_7.SEQ_MODE=4'b1000;
    defparam duty_i15_LC_12_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i15_LC_12_26_7 (
            .in0(_gnd_net_),
            .in1(N__44469),
            .in2(N__50565),
            .in3(N__44457),
            .lcout(duty_15),
            .ltout(),
            .carryin(n12487),
            .carryout(n12488),
            .clk(N__56221),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i16_LC_12_27_0.C_ON=1'b1;
    defparam duty_i16_LC_12_27_0.SEQ_MODE=4'b1000;
    defparam duty_i16_LC_12_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i16_LC_12_27_0 (
            .in0(_gnd_net_),
            .in1(N__47883),
            .in2(N__50517),
            .in3(N__44433),
            .lcout(duty_16),
            .ltout(),
            .carryin(bfn_12_27_0_),
            .carryout(n12489),
            .clk(N__56226),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i17_LC_12_27_1.C_ON=1'b1;
    defparam duty_i17_LC_12_27_1.SEQ_MODE=4'b1000;
    defparam duty_i17_LC_12_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i17_LC_12_27_1 (
            .in0(_gnd_net_),
            .in1(N__44430),
            .in2(N__50481),
            .in3(N__44418),
            .lcout(duty_17),
            .ltout(),
            .carryin(n12489),
            .carryout(n12490),
            .clk(N__56226),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i18_LC_12_27_2.C_ON=1'b1;
    defparam duty_i18_LC_12_27_2.SEQ_MODE=4'b1000;
    defparam duty_i18_LC_12_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i18_LC_12_27_2 (
            .in0(_gnd_net_),
            .in1(N__44415),
            .in2(N__50436),
            .in3(N__44406),
            .lcout(duty_18),
            .ltout(),
            .carryin(n12490),
            .carryout(n12491),
            .clk(N__56226),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i19_LC_12_27_3.C_ON=1'b1;
    defparam duty_i19_LC_12_27_3.SEQ_MODE=4'b1000;
    defparam duty_i19_LC_12_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i19_LC_12_27_3 (
            .in0(_gnd_net_),
            .in1(N__44403),
            .in2(N__50396),
            .in3(N__44394),
            .lcout(duty_19),
            .ltout(),
            .carryin(n12491),
            .carryout(n12492),
            .clk(N__56226),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i20_LC_12_27_4.C_ON=1'b1;
    defparam duty_i20_LC_12_27_4.SEQ_MODE=4'b1000;
    defparam duty_i20_LC_12_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i20_LC_12_27_4 (
            .in0(_gnd_net_),
            .in1(N__44391),
            .in2(N__51300),
            .in3(N__44379),
            .lcout(duty_20),
            .ltout(),
            .carryin(n12492),
            .carryout(n12493),
            .clk(N__56226),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i21_LC_12_27_5.C_ON=1'b1;
    defparam duty_i21_LC_12_27_5.SEQ_MODE=4'b1000;
    defparam duty_i21_LC_12_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i21_LC_12_27_5 (
            .in0(_gnd_net_),
            .in1(N__44376),
            .in2(N__51270),
            .in3(N__44367),
            .lcout(duty_21),
            .ltout(),
            .carryin(n12493),
            .carryout(n12494),
            .clk(N__56226),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i22_LC_12_27_6.C_ON=1'b1;
    defparam duty_i22_LC_12_27_6.SEQ_MODE=4'b1000;
    defparam duty_i22_LC_12_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 duty_i22_LC_12_27_6 (
            .in0(_gnd_net_),
            .in1(N__44364),
            .in2(N__51228),
            .in3(N__44355),
            .lcout(duty_22),
            .ltout(),
            .carryin(n12494),
            .carryout(n12495),
            .clk(N__56226),
            .ce(),
            .sr(_gnd_net_));
    defparam duty_i23_LC_12_27_7.C_ON=1'b0;
    defparam duty_i23_LC_12_27_7.SEQ_MODE=4'b1000;
    defparam duty_i23_LC_12_27_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 duty_i23_LC_12_27_7 (
            .in0(N__51054),
            .in1(N__44352),
            .in2(_gnd_net_),
            .in3(N__44343),
            .lcout(duty_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56226),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i18_1_lut_LC_12_28_0.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i18_1_lut_LC_12_28_0.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i18_1_lut_LC_12_28_0.LUT_INIT=16'b0011001100110011;
    LogicCell40 unary_minus_13_inv_0_i18_1_lut_LC_12_28_0 (
            .in0(_gnd_net_),
            .in1(N__44591),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n8_adj_580),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i22_1_lut_LC_12_28_1.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i22_1_lut_LC_12_28_1.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i22_1_lut_LC_12_28_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i22_1_lut_LC_12_28_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44570),
            .lcout(n4_adj_576),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i19_1_lut_LC_12_28_2.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i19_1_lut_LC_12_28_2.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i19_1_lut_LC_12_28_2.LUT_INIT=16'b0101010101010101;
    LogicCell40 unary_minus_13_inv_0_i19_1_lut_LC_12_28_2 (
            .in0(N__44543),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n7_adj_579),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i19_LC_12_28_3.C_ON=1'b0;
    defparam pwm_setpoint_i19_LC_12_28_3.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i19_LC_12_28_3.LUT_INIT=16'b1111101001010000;
    LogicCell40 pwm_setpoint_i19_LC_12_28_3 (
            .in0(N__50833),
            .in1(_gnd_net_),
            .in2(N__46752),
            .in3(N__44526),
            .lcout(pwm_setpoint_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56231),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i20_LC_12_28_4.C_ON=1'b0;
    defparam pwm_setpoint_i20_LC_12_28_4.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i20_LC_12_28_4.LUT_INIT=16'b1110111000100010;
    LogicCell40 pwm_setpoint_i20_LC_12_28_4 (
            .in0(N__44484),
            .in1(N__50834),
            .in2(_gnd_net_),
            .in3(N__44520),
            .lcout(pwm_setpoint_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56231),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i4_4_lut_LC_12_28_5.C_ON=1'b0;
    defparam LessThan_299_i4_4_lut_LC_12_28_5.SEQ_MODE=4'b0000;
    defparam LessThan_299_i4_4_lut_LC_12_28_5.LUT_INIT=16'b0100110101000100;
    LogicCell40 LessThan_299_i4_4_lut_LC_12_28_5 (
            .in0(N__48156),
            .in1(N__47940),
            .in2(N__48177),
            .in3(N__44490),
            .lcout(n4_adj_655),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i0_LC_12_28_6.C_ON=1'b0;
    defparam pwm_setpoint_i0_LC_12_28_6.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i0_LC_12_28_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 pwm_setpoint_i0_LC_12_28_6 (
            .in0(N__44514),
            .in1(N__50832),
            .in2(_gnd_net_),
            .in3(N__44505),
            .lcout(pwm_setpoint_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56231),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i21_1_lut_LC_12_28_7.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i21_1_lut_LC_12_28_7.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i21_1_lut_LC_12_28_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i21_1_lut_LC_12_28_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44483),
            .lcout(n5_adj_577),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i45_2_lut_LC_12_29_0.C_ON=1'b0;
    defparam LessThan_299_i45_2_lut_LC_12_29_0.SEQ_MODE=4'b0000;
    defparam LessThan_299_i45_2_lut_LC_12_29_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i45_2_lut_LC_12_29_0 (
            .in0(_gnd_net_),
            .in1(N__44711),
            .in2(_gnd_net_),
            .in3(N__48432),
            .lcout(n45),
            .ltout(n45_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12515_4_lut_LC_12_29_1.C_ON=1'b0;
    defparam i12515_4_lut_LC_12_29_1.SEQ_MODE=4'b0000;
    defparam i12515_4_lut_LC_12_29_1.LUT_INIT=16'b1010101110101000;
    LogicCell40 i12515_4_lut_LC_12_29_1 (
            .in0(N__44649),
            .in1(N__44838),
            .in2(N__44700),
            .in3(N__44685),
            .lcout(n15245),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i41_2_lut_LC_12_29_2.C_ON=1'b0;
    defparam LessThan_299_i41_2_lut_LC_12_29_2.SEQ_MODE=4'b0000;
    defparam LessThan_299_i41_2_lut_LC_12_29_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i41_2_lut_LC_12_29_2 (
            .in0(_gnd_net_),
            .in1(N__44696),
            .in2(_gnd_net_),
            .in3(N__48504),
            .lcout(n41_adj_678),
            .ltout(n41_adj_678_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12522_3_lut_LC_12_29_3.C_ON=1'b0;
    defparam i12522_3_lut_LC_12_29_3.SEQ_MODE=4'b0000;
    defparam i12522_3_lut_LC_12_29_3.LUT_INIT=16'b1010111110100000;
    LogicCell40 i12522_3_lut_LC_12_29_3 (
            .in0(N__44697),
            .in1(_gnd_net_),
            .in2(N__44688),
            .in3(N__44604),
            .lcout(n40_adj_677),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12513_4_lut_LC_12_29_4.C_ON=1'b0;
    defparam i12513_4_lut_LC_12_29_4.SEQ_MODE=4'b0000;
    defparam i12513_4_lut_LC_12_29_4.LUT_INIT=16'b1100110111001000;
    LogicCell40 i12513_4_lut_LC_12_29_4 (
            .in0(N__44679),
            .in1(N__44664),
            .in2(N__44757),
            .in3(N__44658),
            .lcout(n15243),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i23_1_lut_LC_12_29_5.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i23_1_lut_LC_12_29_5.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i23_1_lut_LC_12_29_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i23_1_lut_LC_12_29_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44639),
            .lcout(n3_adj_575),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i13_2_lut_LC_12_29_6.C_ON=1'b0;
    defparam LessThan_299_i13_2_lut_LC_12_29_6.SEQ_MODE=4'b0000;
    defparam LessThan_299_i13_2_lut_LC_12_29_6.LUT_INIT=16'b0101010110101010;
    LogicCell40 LessThan_299_i13_2_lut_LC_12_29_6 (
            .in0(N__46208),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48056),
            .lcout(n13_adj_662),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i39_2_lut_LC_12_30_0.C_ON=1'b0;
    defparam LessThan_299_i39_2_lut_LC_12_30_0.SEQ_MODE=4'b0000;
    defparam LessThan_299_i39_2_lut_LC_12_30_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i39_2_lut_LC_12_30_0 (
            .in0(_gnd_net_),
            .in1(N__44618),
            .in2(_gnd_net_),
            .in3(N__48528),
            .lcout(n39_adj_676),
            .ltout(n39_adj_676_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12524_3_lut_LC_12_30_1.C_ON=1'b0;
    defparam i12524_3_lut_LC_12_30_1.SEQ_MODE=4'b0000;
    defparam i12524_3_lut_LC_12_30_1.LUT_INIT=16'b1010111110100000;
    LogicCell40 i12524_3_lut_LC_12_30_1 (
            .in0(N__44619),
            .in1(_gnd_net_),
            .in2(N__44607),
            .in3(N__44997),
            .lcout(n15254),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i43_2_lut_LC_12_30_2.C_ON=1'b0;
    defparam LessThan_299_i43_2_lut_LC_12_30_2.SEQ_MODE=4'b0000;
    defparam LessThan_299_i43_2_lut_LC_12_30_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i43_2_lut_LC_12_30_2 (
            .in0(_gnd_net_),
            .in1(N__48476),
            .in2(_gnd_net_),
            .in3(N__44880),
            .lcout(n43),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i12_LC_12_30_3.C_ON=1'b0;
    defparam pwm_setpoint_i12_LC_12_30_3.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i12_LC_12_30_3.LUT_INIT=16'b1110111001000100;
    LogicCell40 pwm_setpoint_i12_LC_12_30_3 (
            .in0(N__50873),
            .in1(N__44955),
            .in2(_gnd_net_),
            .in3(N__44865),
            .lcout(pwm_setpoint_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56244),
            .ce(),
            .sr(_gnd_net_));
    defparam i12361_4_lut_LC_12_30_4.C_ON=1'b0;
    defparam i12361_4_lut_LC_12_30_4.SEQ_MODE=4'b0000;
    defparam i12361_4_lut_LC_12_30_4.LUT_INIT=16'b1010101010101011;
    LogicCell40 i12361_4_lut_LC_12_30_4 (
            .in0(N__44766),
            .in1(N__44856),
            .in2(N__44850),
            .in3(N__44907),
            .lcout(n15091),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12499_3_lut_LC_12_30_5.C_ON=1'b0;
    defparam i12499_3_lut_LC_12_30_5.SEQ_MODE=4'b0000;
    defparam i12499_3_lut_LC_12_30_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 i12499_3_lut_LC_12_30_5 (
            .in0(N__46575),
            .in1(N__46540),
            .in2(_gnd_net_),
            .in3(N__44829),
            .lcout(n15229),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i25_2_lut_LC_12_30_6.C_ON=1'b0;
    defparam LessThan_299_i25_2_lut_LC_12_30_6.SEQ_MODE=4'b0000;
    defparam LessThan_299_i25_2_lut_LC_12_30_6.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i25_2_lut_LC_12_30_6 (
            .in0(_gnd_net_),
            .in1(N__44819),
            .in2(_gnd_net_),
            .in3(N__48318),
            .lcout(n25_adj_670),
            .ltout(n25_adj_670_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12416_4_lut_LC_12_30_7.C_ON=1'b0;
    defparam i12416_4_lut_LC_12_30_7.SEQ_MODE=4'b0000;
    defparam i12416_4_lut_LC_12_30_7.LUT_INIT=16'b1111111100000001;
    LogicCell40 i12416_4_lut_LC_12_30_7 (
            .in0(N__44799),
            .in1(N__44788),
            .in2(N__44769),
            .in3(N__44765),
            .lcout(n15146),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam commutation_state_i1_LC_12_31_0.C_ON=1'b0;
    defparam commutation_state_i1_LC_12_31_0.SEQ_MODE=4'b1000;
    defparam commutation_state_i1_LC_12_31_0.LUT_INIT=16'b1010001100100010;
    LogicCell40 commutation_state_i1_LC_12_31_0 (
            .in0(N__47005),
            .in1(N__46957),
            .in2(N__46905),
            .in3(N__56319),
            .lcout(commutation_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56250),
            .ce(),
            .sr(_gnd_net_));
    defparam i12374_4_lut_LC_12_31_1.C_ON=1'b0;
    defparam i12374_4_lut_LC_12_31_1.SEQ_MODE=4'b0000;
    defparam i12374_4_lut_LC_12_31_1.LUT_INIT=16'b1010101010101011;
    LogicCell40 i12374_4_lut_LC_12_31_1 (
            .in0(N__46547),
            .in1(N__44748),
            .in2(N__46805),
            .in3(N__44732),
            .lcout(n15104),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12500_3_lut_LC_12_31_2.C_ON=1'b0;
    defparam i12500_3_lut_LC_12_31_2.SEQ_MODE=4'b0000;
    defparam i12500_3_lut_LC_12_31_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 i12500_3_lut_LC_12_31_2 (
            .in0(N__46784),
            .in1(N__46765),
            .in2(_gnd_net_),
            .in3(N__44721),
            .lcout(n15230),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i10_3_lut_3_lut_LC_12_31_3.C_ON=1'b0;
    defparam LessThan_299_i10_3_lut_3_lut_LC_12_31_3.SEQ_MODE=4'b0000;
    defparam LessThan_299_i10_3_lut_3_lut_LC_12_31_3.LUT_INIT=16'b1000100011101110;
    LogicCell40 LessThan_299_i10_3_lut_3_lut_LC_12_31_3 (
            .in0(N__46830),
            .in1(N__46212),
            .in2(_gnd_net_),
            .in3(N__48057),
            .lcout(n10_adj_659),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i13_1_lut_LC_12_31_4.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i13_1_lut_LC_12_31_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i13_1_lut_LC_12_31_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i13_1_lut_LC_12_31_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44954),
            .lcout(n13_adj_585),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_3_lut_LC_12_31_5.C_ON=1'b0;
    defparam i2_2_lut_3_lut_LC_12_31_5.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_LC_12_31_5.LUT_INIT=16'b0000000000100010;
    LogicCell40 i2_2_lut_3_lut_LC_12_31_5 (
            .in0(N__46956),
            .in1(N__47004),
            .in2(_gnd_net_),
            .in3(N__46899),
            .lcout(commutation_state_7__N_261),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i31_2_lut_LC_12_31_6.C_ON=1'b0;
    defparam LessThan_299_i31_2_lut_LC_12_31_6.SEQ_MODE=4'b0000;
    defparam LessThan_299_i31_2_lut_LC_12_31_6.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i31_2_lut_LC_12_31_6 (
            .in0(_gnd_net_),
            .in1(N__46475),
            .in2(_gnd_net_),
            .in3(N__48242),
            .lcout(n31_adj_674),
            .ltout(n31_adj_674_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12490_3_lut_LC_12_31_7.C_ON=1'b0;
    defparam i12490_3_lut_LC_12_31_7.SEQ_MODE=4'b0000;
    defparam i12490_3_lut_LC_12_31_7.LUT_INIT=16'b1010111110100000;
    LogicCell40 i12490_3_lut_LC_12_31_7 (
            .in0(N__46476),
            .in1(_gnd_net_),
            .in2(N__44925),
            .in3(N__44922),
            .lcout(n15220),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12465_4_lut_LC_12_32_0.C_ON=1'b0;
    defparam i12465_4_lut_LC_12_32_0.SEQ_MODE=4'b0000;
    defparam i12465_4_lut_LC_12_32_0.LUT_INIT=16'b1111111111111011;
    LogicCell40 i12465_4_lut_LC_12_32_0 (
            .in0(N__45060),
            .in1(N__44916),
            .in2(N__46770),
            .in3(N__46548),
            .lcout(),
            .ltout(n15195_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12511_4_lut_LC_12_32_1.C_ON=1'b0;
    defparam i12511_4_lut_LC_12_32_1.SEQ_MODE=4'b0000;
    defparam i12511_4_lut_LC_12_32_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12511_4_lut_LC_12_32_1 (
            .in0(N__45078),
            .in1(N__45006),
            .in2(N__44910),
            .in3(N__45050),
            .lcout(n15241),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i37_2_lut_LC_12_32_3.C_ON=1'b0;
    defparam LessThan_299_i37_2_lut_LC_12_32_3.SEQ_MODE=4'b0000;
    defparam LessThan_299_i37_2_lut_LC_12_32_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i37_2_lut_LC_12_32_3 (
            .in0(_gnd_net_),
            .in1(N__45020),
            .in2(_gnd_net_),
            .in3(N__48555),
            .lcout(n37),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12517_4_lut_LC_12_32_4.C_ON=1'b0;
    defparam i12517_4_lut_LC_12_32_4.SEQ_MODE=4'b0000;
    defparam i12517_4_lut_LC_12_32_4.LUT_INIT=16'b1111111000000100;
    LogicCell40 i12517_4_lut_LC_12_32_4 (
            .in0(N__44898),
            .in1(N__44892),
            .in2(N__45051),
            .in3(N__44886),
            .lcout(n15247),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12369_4_lut_LC_12_32_5.C_ON=1'b0;
    defparam i12369_4_lut_LC_12_32_5.SEQ_MODE=4'b0000;
    defparam i12369_4_lut_LC_12_32_5.LUT_INIT=16'b1010101010101011;
    LogicCell40 i12369_4_lut_LC_12_32_5 (
            .in0(N__45077),
            .in1(N__46766),
            .in2(N__45069),
            .in3(N__45059),
            .lcout(),
            .ltout(n15099_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12527_4_lut_LC_12_32_6.C_ON=1'b0;
    defparam i12527_4_lut_LC_12_32_6.SEQ_MODE=4'b0000;
    defparam i12527_4_lut_LC_12_32_6.LUT_INIT=16'b1100110111001000;
    LogicCell40 i12527_4_lut_LC_12_32_6 (
            .in0(N__45049),
            .in1(N__45036),
            .in2(N__45030),
            .in3(N__45027),
            .lcout(),
            .ltout(n15257_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12528_3_lut_LC_12_32_7.C_ON=1'b0;
    defparam i12528_3_lut_LC_12_32_7.SEQ_MODE=4'b0000;
    defparam i12528_3_lut_LC_12_32_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 i12528_3_lut_LC_12_32_7 (
            .in0(_gnd_net_),
            .in1(N__45021),
            .in2(N__45009),
            .in3(N__45005),
            .lcout(n15258),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_2_lut_LC_13_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_2_lut_LC_13_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_2_lut_LC_13_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_2_lut_LC_13_17_0 (
            .in0(_gnd_net_),
            .in1(N__48788),
            .in2(_gnd_net_),
            .in3(N__44988),
            .lcout(n1701),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(n12577),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_3_lut_LC_13_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_3_lut_LC_13_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_3_lut_LC_13_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_3_lut_LC_13_17_1 (
            .in0(_gnd_net_),
            .in1(N__53850),
            .in2(N__48749),
            .in3(N__44976),
            .lcout(n1700),
            .ltout(),
            .carryin(n12577),
            .carryout(n12578),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_4_lut_LC_13_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_4_lut_LC_13_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_4_lut_LC_13_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_4_lut_LC_13_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__48809),
            .in3(N__44964),
            .lcout(n1699),
            .ltout(),
            .carryin(n12578),
            .carryout(n12579),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_5_lut_LC_13_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_5_lut_LC_13_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_5_lut_LC_13_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_5_lut_LC_13_17_3 (
            .in0(_gnd_net_),
            .in1(N__53851),
            .in2(N__48926),
            .in3(N__44961),
            .lcout(n1698),
            .ltout(),
            .carryin(n12579),
            .carryout(n12580),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_6_lut_LC_13_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_6_lut_LC_13_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_6_lut_LC_13_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_6_lut_LC_13_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47081),
            .in3(N__44958),
            .lcout(n1697),
            .ltout(),
            .carryin(n12580),
            .carryout(n12581),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_7_lut_LC_13_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_7_lut_LC_13_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_7_lut_LC_13_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_7_lut_LC_13_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47063),
            .in3(N__45141),
            .lcout(n1696),
            .ltout(),
            .carryin(n12581),
            .carryout(n12582),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_8_lut_LC_13_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_8_lut_LC_13_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_8_lut_LC_13_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_8_lut_LC_13_17_6 (
            .in0(_gnd_net_),
            .in1(N__47406),
            .in2(N__54246),
            .in3(N__45138),
            .lcout(n1695),
            .ltout(),
            .carryin(n12582),
            .carryout(n12583),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_9_lut_LC_13_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_9_lut_LC_13_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_9_lut_LC_13_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_9_lut_LC_13_17_7 (
            .in0(_gnd_net_),
            .in1(N__53855),
            .in2(N__47207),
            .in3(N__45129),
            .lcout(n1694),
            .ltout(),
            .carryin(n12583),
            .carryout(n12584),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_10_lut_LC_13_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_10_lut_LC_13_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_10_lut_LC_13_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_10_lut_LC_13_18_0 (
            .in0(_gnd_net_),
            .in1(N__53841),
            .in2(N__47340),
            .in3(N__45126),
            .lcout(n1693_adj_614),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(n12585),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_11_lut_LC_13_18_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_11_lut_LC_13_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_11_lut_LC_13_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_11_lut_LC_13_18_1 (
            .in0(_gnd_net_),
            .in1(N__54953),
            .in2(N__45156),
            .in3(N__45123),
            .lcout(n1692),
            .ltout(),
            .carryin(n12585),
            .carryout(n12586),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_12_lut_LC_13_18_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_12_lut_LC_13_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_12_lut_LC_13_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_12_lut_LC_13_18_2 (
            .in0(_gnd_net_),
            .in1(N__53842),
            .in2(N__47276),
            .in3(N__45114),
            .lcout(n1691),
            .ltout(),
            .carryin(n12586),
            .carryout(n12587),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_13_lut_LC_13_18_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_13_lut_LC_13_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_13_lut_LC_13_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_13_lut_LC_13_18_3 (
            .in0(_gnd_net_),
            .in1(N__47246),
            .in2(N__54244),
            .in3(N__45102),
            .lcout(n1690),
            .ltout(),
            .carryin(n12587),
            .carryout(n12588),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_14_lut_LC_13_18_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_14_lut_LC_13_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_14_lut_LC_13_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_14_lut_LC_13_18_4 (
            .in0(_gnd_net_),
            .in1(N__53846),
            .in2(N__47180),
            .in3(N__45090),
            .lcout(n1689),
            .ltout(),
            .carryin(n12588),
            .carryout(n12589),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_15_lut_LC_13_18_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1101_15_lut_LC_13_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_15_lut_LC_13_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1101_15_lut_LC_13_18_5 (
            .in0(_gnd_net_),
            .in1(N__45371),
            .in2(N__54245),
            .in3(N__45081),
            .lcout(n1688),
            .ltout(),
            .carryin(n12589),
            .carryout(n12590),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1101_16_lut_LC_13_18_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1101_16_lut_LC_13_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1101_16_lut_LC_13_18_6.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_1101_16_lut_LC_13_18_6 (
            .in0(N__54954),
            .in1(N__45167),
            .in2(N__52443),
            .in3(N__45348),
            .lcout(n1719),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1111_3_lut_LC_13_18_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1111_3_lut_LC_13_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1111_3_lut_LC_13_18_7.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1111_3_lut_LC_13_18_7 (
            .in0(_gnd_net_),
            .in1(N__45324),
            .in2(N__45617),
            .in3(N__47405),
            .lcout(n1727),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12884_4_lut_LC_13_19_0.C_ON=1'b0;
    defparam i12884_4_lut_LC_13_19_0.SEQ_MODE=4'b0000;
    defparam i12884_4_lut_LC_13_19_0.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12884_4_lut_LC_13_19_0 (
            .in0(N__47173),
            .in1(N__45364),
            .in2(N__47220),
            .in3(N__52439),
            .lcout(n1653),
            .ltout(n1653_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1112_3_lut_LC_13_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1112_3_lut_LC_13_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1112_3_lut_LC_13_19_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1112_3_lut_LC_13_19_1 (
            .in0(_gnd_net_),
            .in1(N__45294),
            .in2(N__45285),
            .in3(N__47064),
            .lcout(n1728),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1113_3_lut_LC_13_19_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1113_3_lut_LC_13_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1113_3_lut_LC_13_19_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1113_3_lut_LC_13_19_2 (
            .in0(_gnd_net_),
            .in1(N__47082),
            .in2(N__45264),
            .in3(N__45586),
            .lcout(n1729),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1108_3_lut_LC_13_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1108_3_lut_LC_13_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1108_3_lut_LC_13_19_3.LUT_INIT=16'b1100101011001010;
    LogicCell40 encoder0_position_31__I_0_i1108_3_lut_LC_13_19_3 (
            .in0(N__45252),
            .in1(N__45155),
            .in2(N__45613),
            .in3(_gnd_net_),
            .lcout(n1724),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1109_3_lut_LC_13_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1109_3_lut_LC_13_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1109_3_lut_LC_13_19_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1109_3_lut_LC_13_19_4 (
            .in0(_gnd_net_),
            .in1(N__47336),
            .in2(N__45219),
            .in3(N__45587),
            .lcout(n1725),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12881_1_lut_LC_13_19_5.C_ON=1'b0;
    defparam i12881_1_lut_LC_13_19_5.SEQ_MODE=4'b0000;
    defparam i12881_1_lut_LC_13_19_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12881_1_lut_LC_13_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45614),
            .in3(_gnd_net_),
            .lcout(n15611),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1041_3_lut_LC_13_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1041_3_lut_LC_13_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1041_3_lut_LC_13_19_6.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i1041_3_lut_LC_13_19_6 (
            .in0(N__51969),
            .in1(_gnd_net_),
            .in2(N__51999),
            .in3(N__48877),
            .lcout(n1625_adj_605),
            .ltout(n1625_adj_605_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_122_LC_13_19_7.C_ON=1'b0;
    defparam i1_4_lut_adj_122_LC_13_19_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_122_LC_13_19_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_122_LC_13_19_7 (
            .in0(N__47335),
            .in1(N__47200),
            .in2(N__45714),
            .in3(N__47401),
            .lcout(n14502),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1114_3_lut_LC_13_20_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1114_3_lut_LC_13_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1114_3_lut_LC_13_20_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1114_3_lut_LC_13_20_0 (
            .in0(_gnd_net_),
            .in1(N__45711),
            .in2(N__48930),
            .in3(N__45597),
            .lcout(n1730),
            .ltout(n1730_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_134_LC_13_20_1.C_ON=1'b0;
    defparam i1_2_lut_adj_134_LC_13_20_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_134_LC_13_20_1.LUT_INIT=16'b1111000000000000;
    LogicCell40 i1_2_lut_adj_134_LC_13_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45684),
            .in3(N__45670),
            .lcout(n14514),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut_LC_13_20_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut_LC_13_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut_LC_13_20_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut_LC_13_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47365),
            .lcout(n11_adj_629),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1117_3_lut_LC_13_20_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1117_3_lut_LC_13_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1117_3_lut_LC_13_20_3.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1117_3_lut_LC_13_20_3 (
            .in0(_gnd_net_),
            .in1(N__45630),
            .in2(N__45615),
            .in3(N__48789),
            .lcout(n1733),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12900_1_lut_LC_13_20_4.C_ON=1'b0;
    defparam i12900_1_lut_LC_13_20_4.SEQ_MODE=4'b0000;
    defparam i12900_1_lut_LC_13_20_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12900_1_lut_LC_13_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45480),
            .lcout(n15630),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1037_3_lut_LC_13_20_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1037_3_lut_LC_13_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1037_3_lut_LC_13_20_5.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i1037_3_lut_LC_13_20_5 (
            .in0(N__52536),
            .in1(N__52509),
            .in2(N__48893),
            .in3(_gnd_net_),
            .lcout(n1621_adj_601),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_new_i1_LC_13_21_1 .C_ON=1'b0;
    defparam \quad_counter0.b_new_i1_LC_13_21_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_new_i1_LC_13_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter0.b_new_i1_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46417),
            .lcout(\quad_counter0.b_new_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56213),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_new_i0_LC_13_21_4 .C_ON=1'b0;
    defparam \quad_counter0.b_new_i0_LC_13_21_4 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_new_i0_LC_13_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter0.b_new_i0_LC_13_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45822),
            .lcout(\quad_counter0.b_new_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56213),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i707_3_lut_LC_13_22_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i707_3_lut_LC_13_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i707_3_lut_LC_13_22_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i707_3_lut_LC_13_22_0 (
            .in0(_gnd_net_),
            .in1(N__53017),
            .in2(N__49860),
            .in3(N__52995),
            .lcout(n1131),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut_LC_13_22_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut_LC_13_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut_LC_13_22_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut_LC_13_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45800),
            .lcout(n32_adj_650),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut_LC_13_22_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut_LC_13_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut_LC_13_22_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut_LC_13_22_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45758),
            .lcout(n17_adj_635),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i705_3_lut_LC_13_22_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i705_3_lut_LC_13_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i705_3_lut_LC_13_22_4.LUT_INIT=16'b1111010110100000;
    LogicCell40 encoder0_position_31__I_0_i705_3_lut_LC_13_22_4 (
            .in0(N__49842),
            .in1(_gnd_net_),
            .in2(N__52937),
            .in3(N__52911),
            .lcout(n1129),
            .ltout(n1129_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_99_LC_13_22_5.C_ON=1'b0;
    defparam i1_2_lut_adj_99_LC_13_22_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_99_LC_13_22_5.LUT_INIT=16'b1111000000000000;
    LogicCell40 i1_2_lut_adj_99_LC_13_22_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45717),
            .in3(N__47536),
            .lcout(n14464),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i706_3_lut_LC_13_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i706_3_lut_LC_13_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i706_3_lut_LC_13_22_7.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i706_3_lut_LC_13_22_7 (
            .in0(_gnd_net_),
            .in1(N__49841),
            .in2(N__52979),
            .in3(N__52953),
            .lcout(n1130),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i702_3_lut_LC_13_23_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i702_3_lut_LC_13_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i702_3_lut_LC_13_23_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i702_3_lut_LC_13_23_0 (
            .in0(_gnd_net_),
            .in1(N__55592),
            .in2(N__49868),
            .in3(N__55575),
            .lcout(n1126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i638_3_lut_LC_13_23_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i638_3_lut_LC_13_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i638_3_lut_LC_13_23_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i638_3_lut_LC_13_23_1 (
            .in0(_gnd_net_),
            .in1(N__45854),
            .in2(N__45834),
            .in3(N__46008),
            .lcout(n1030),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9957_3_lut_LC_13_23_2.C_ON=1'b0;
    defparam i9957_3_lut_LC_13_23_2.SEQ_MODE=4'b0000;
    defparam i9957_3_lut_LC_13_23_2.LUT_INIT=16'b1111000011000000;
    LogicCell40 i9957_3_lut_LC_13_23_2 (
            .in0(_gnd_net_),
            .in1(N__53083),
            .in2(N__53021),
            .in3(N__53050),
            .lcout(),
            .ltout(n11933_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_92_LC_13_23_3.C_ON=1'b0;
    defparam i1_4_lut_adj_92_LC_13_23_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_92_LC_13_23_3.LUT_INIT=16'b1010100000000000;
    LogicCell40 i1_4_lut_adj_92_LC_13_23_3 (
            .in0(N__52885),
            .in1(N__52972),
            .in2(N__45936),
            .in3(N__52930),
            .lcout(),
            .ltout(n13728_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12781_4_lut_LC_13_23_4.C_ON=1'b0;
    defparam i12781_4_lut_LC_13_23_4.SEQ_MODE=4'b0000;
    defparam i12781_4_lut_LC_13_23_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12781_4_lut_LC_13_23_4 (
            .in0(N__52852),
            .in1(N__53377),
            .in2(N__45933),
            .in3(N__55591),
            .lcout(n1059),
            .ltout(n1059_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i709_3_lut_LC_13_23_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i709_3_lut_LC_13_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i709_3_lut_LC_13_23_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i709_3_lut_LC_13_23_5 (
            .in0(N__53084),
            .in1(_gnd_net_),
            .in2(N__45930),
            .in3(N__53070),
            .lcout(n1133),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i708_3_lut_LC_13_23_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i708_3_lut_LC_13_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i708_3_lut_LC_13_23_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i708_3_lut_LC_13_23_6 (
            .in0(_gnd_net_),
            .in1(N__53034),
            .in2(N__49867),
            .in3(N__53051),
            .lcout(n1132),
            .ltout(n1132_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10042_4_lut_LC_13_23_7.C_ON=1'b0;
    defparam i10042_4_lut_LC_13_23_7.SEQ_MODE=4'b0000;
    defparam i10042_4_lut_LC_13_23_7.LUT_INIT=16'b1111101011101010;
    LogicCell40 i10042_4_lut_LC_13_23_7 (
            .in0(N__47572),
            .in1(N__47647),
            .in2(N__45927),
            .in3(N__47611),
            .lcout(n12019),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_2_lut_LC_13_24_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_2_lut_LC_13_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_2_lut_LC_13_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_2_lut_LC_13_24_0 (
            .in0(_gnd_net_),
            .in1(N__45923),
            .in2(_gnd_net_),
            .in3(N__45906),
            .lcout(n1001),
            .ltout(),
            .carryin(bfn_13_24_0_),
            .carryout(n12507),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_3_lut_LC_13_24_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_3_lut_LC_13_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_3_lut_LC_13_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_3_lut_LC_13_24_1 (
            .in0(_gnd_net_),
            .in1(N__53785),
            .in2(N__45903),
            .in3(N__45882),
            .lcout(n1000),
            .ltout(),
            .carryin(n12507),
            .carryout(n12508),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_4_lut_LC_13_24_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_4_lut_LC_13_24_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_4_lut_LC_13_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_4_lut_LC_13_24_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45879),
            .in3(N__45858),
            .lcout(n999),
            .ltout(),
            .carryin(n12508),
            .carryout(n12509),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_5_lut_LC_13_24_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_5_lut_LC_13_24_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_5_lut_LC_13_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_5_lut_LC_13_24_3 (
            .in0(_gnd_net_),
            .in1(N__53786),
            .in2(N__45855),
            .in3(N__46110),
            .lcout(n998),
            .ltout(),
            .carryin(n12509),
            .carryout(n12510),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_6_lut_LC_13_24_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_6_lut_LC_13_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_6_lut_LC_13_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_6_lut_LC_13_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46107),
            .in3(N__46074),
            .lcout(n997),
            .ltout(),
            .carryin(n12510),
            .carryout(n12511),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_7_lut_LC_13_24_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_7_lut_LC_13_24_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_7_lut_LC_13_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_7_lut_LC_13_24_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46071),
            .in3(N__46044),
            .lcout(n996),
            .ltout(),
            .carryin(n12511),
            .carryout(n12512),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_8_lut_LC_13_24_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_632_8_lut_LC_13_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_8_lut_LC_13_24_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_632_8_lut_LC_13_24_6 (
            .in0(_gnd_net_),
            .in1(N__53787),
            .in2(N__46041),
            .in3(N__46017),
            .lcout(n995),
            .ltout(),
            .carryin(n12512),
            .carryout(n12513),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_632_9_lut_LC_13_24_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_632_9_lut_LC_13_24_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_632_9_lut_LC_13_24_7.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_632_9_lut_LC_13_24_7 (
            .in0(N__53788),
            .in1(N__46012),
            .in2(N__45975),
            .in3(N__45957),
            .lcout(n1026),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i1_1_lut_LC_13_25_1.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i1_1_lut_LC_13_25_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i1_1_lut_LC_13_25_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i1_1_lut_LC_13_25_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45954),
            .lcout(n25_adj_551),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9898_2_lut_LC_13_25_2.C_ON=1'b0;
    defparam i9898_2_lut_LC_13_25_2.SEQ_MODE=4'b0000;
    defparam i9898_2_lut_LC_13_25_2.LUT_INIT=16'b1111111111001100;
    LogicCell40 i9898_2_lut_LC_13_25_2 (
            .in0(_gnd_net_),
            .in1(N__50265),
            .in2(_gnd_net_),
            .in3(N__50310),
            .lcout(),
            .ltout(n11872_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_adj_52_LC_13_25_3.C_ON=1'b0;
    defparam i4_4_lut_adj_52_LC_13_25_3.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_52_LC_13_25_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 i4_4_lut_adj_52_LC_13_25_3 (
            .in0(N__50071),
            .in1(N__50191),
            .in2(N__45939),
            .in3(N__50232),
            .lcout(n10_adj_681),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_LC_13_25_4.C_ON=1'b0;
    defparam i3_4_lut_LC_13_25_4.SEQ_MODE=4'b0000;
    defparam i3_4_lut_LC_13_25_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i3_4_lut_LC_13_25_4 (
            .in0(N__49763),
            .in1(N__50347),
            .in2(N__49736),
            .in3(N__49699),
            .lcout(),
            .ltout(n14034_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_LC_13_25_5.C_ON=1'b0;
    defparam i2_3_lut_LC_13_25_5.SEQ_MODE=4'b0000;
    defparam i2_3_lut_LC_13_25_5.LUT_INIT=16'b1010000000000000;
    LogicCell40 i2_3_lut_LC_13_25_5 (
            .in0(N__50266),
            .in1(_gnd_net_),
            .in2(N__46173),
            .in3(N__50318),
            .lcout(),
            .ltout(n14116_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_51_LC_13_25_6.C_ON=1'b0;
    defparam i1_4_lut_adj_51_LC_13_25_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_51_LC_13_25_6.LUT_INIT=16'b1100110011001000;
    LogicCell40 i1_4_lut_adj_51_LC_13_25_6 (
            .in0(N__50117),
            .in1(N__50476),
            .in2(N__46170),
            .in3(N__46167),
            .lcout(n15_adj_680),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_LC_13_25_7.C_ON=1'b0;
    defparam i4_4_lut_LC_13_25_7.SEQ_MODE=4'b0000;
    defparam i4_4_lut_LC_13_25_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i4_4_lut_LC_13_25_7 (
            .in0(N__50072),
            .in1(N__50233),
            .in2(N__50198),
            .in3(N__50153),
            .lcout(n10_adj_598),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_LC_13_26_0.C_ON=1'b0;
    defparam i10_4_lut_LC_13_26_0.SEQ_MODE=4'b0000;
    defparam i10_4_lut_LC_13_26_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 i10_4_lut_LC_13_26_0 (
            .in0(N__51266),
            .in1(N__50557),
            .in2(N__50397),
            .in3(N__51050),
            .lcout(n24_adj_653),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i2_LC_13_26_1.C_ON=1'b0;
    defparam pwm_setpoint_i2_LC_13_26_1.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i2_LC_13_26_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 pwm_setpoint_i2_LC_13_26_1 (
            .in0(N__50836),
            .in1(N__46161),
            .in2(_gnd_net_),
            .in3(N__46526),
            .lcout(pwm_setpoint_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56227),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i3_LC_13_26_2.C_ON=1'b0;
    defparam pwm_setpoint_i3_LC_13_26_2.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i3_LC_13_26_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 pwm_setpoint_i3_LC_13_26_2 (
            .in0(N__50837),
            .in1(N__46152),
            .in2(_gnd_net_),
            .in3(N__46143),
            .lcout(pwm_setpoint_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56227),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_70_LC_13_26_3.C_ON=1'b0;
    defparam i1_4_lut_adj_70_LC_13_26_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_70_LC_13_26_3.LUT_INIT=16'b1110101010101010;
    LogicCell40 i1_4_lut_adj_70_LC_13_26_3 (
            .in0(N__50392),
            .in1(N__50107),
            .in2(N__46131),
            .in3(N__50151),
            .lcout(n15_adj_711),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_adj_53_LC_13_26_5.C_ON=1'b0;
    defparam i2_2_lut_adj_53_LC_13_26_5.SEQ_MODE=4'b0000;
    defparam i2_2_lut_adj_53_LC_13_26_5.LUT_INIT=16'b1111111110101010;
    LogicCell40 i2_2_lut_adj_53_LC_13_26_5 (
            .in0(N__50670),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51265),
            .lcout(),
            .ltout(n16_adj_710_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11_4_lut_adj_73_LC_13_26_6.C_ON=1'b0;
    defparam i11_4_lut_adj_73_LC_13_26_6.SEQ_MODE=4'b0000;
    defparam i11_4_lut_adj_73_LC_13_26_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i11_4_lut_adj_73_LC_13_26_6 (
            .in0(N__50630),
            .in1(N__51227),
            .in2(N__46122),
            .in3(N__46119),
            .lcout(n25_adj_707),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i3_1_lut_LC_13_27_0.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i3_1_lut_LC_13_27_0.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i3_1_lut_LC_13_27_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i3_1_lut_LC_13_27_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46527),
            .lcout(n23_adj_595),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i15_LC_13_27_4.C_ON=1'b0;
    defparam pwm_setpoint_i15_LC_13_27_4.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i15_LC_13_27_4.LUT_INIT=16'b1110111001000100;
    LogicCell40 pwm_setpoint_i15_LC_13_27_4 (
            .in0(N__50835),
            .in1(N__46499),
            .in2(_gnd_net_),
            .in3(N__46485),
            .lcout(pwm_setpoint_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56232),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.a_new_i1_LC_13_27_5 .C_ON=1'b0;
    defparam \quad_counter0.a_new_i1_LC_13_27_5 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.a_new_i1_LC_13_27_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \quad_counter0.a_new_i1_LC_13_27_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46461),
            .lcout(a_new_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56232),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.i12534_4_lut_LC_13_28_0 .C_ON=1'b0;
    defparam \quad_counter0.i12534_4_lut_LC_13_28_0 .SEQ_MODE=4'b0000;
    defparam \quad_counter0.i12534_4_lut_LC_13_28_0 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \quad_counter0.i12534_4_lut_LC_13_28_0  (
            .in0(N__46456),
            .in1(N__46424),
            .in2(N__46393),
            .in3(N__46332),
            .lcout(\quad_counter0.a_prev_N_543 ),
            .ltout(\quad_counter0.a_prev_N_543_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \quad_counter0.b_prev_52_LC_13_28_1 .C_ON=1'b0;
    defparam \quad_counter0.b_prev_52_LC_13_28_1 .SEQ_MODE=4'b1000;
    defparam \quad_counter0.b_prev_52_LC_13_28_1 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \quad_counter0.b_prev_52_LC_13_28_1  (
            .in0(N__46333),
            .in1(N__46307),
            .in2(N__46281),
            .in3(N__46269),
            .lcout(b_prev),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56238),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i2_3_lut_LC_13_28_2 .C_ON=1'b0;
    defparam \PWM.i2_3_lut_LC_13_28_2 .SEQ_MODE=4'b0000;
    defparam \PWM.i2_3_lut_LC_13_28_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \PWM.i2_3_lut_LC_13_28_2  (
            .in0(N__48080),
            .in1(N__48048),
            .in2(_gnd_net_),
            .in3(N__48009),
            .lcout(\PWM.n13991 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12391_3_lut_4_lut_LC_13_28_3.C_ON=1'b0;
    defparam i12391_3_lut_4_lut_LC_13_28_3.SEQ_MODE=4'b0000;
    defparam i12391_3_lut_4_lut_LC_13_28_3.LUT_INIT=16'b0111101111011110;
    LogicCell40 i12391_3_lut_4_lut_LC_13_28_3 (
            .in0(N__46196),
            .in1(N__46184),
            .in2(N__48138),
            .in3(N__48118),
            .lcout(n15121),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i6_LC_13_28_4.C_ON=1'b0;
    defparam pwm_setpoint_i6_LC_13_28_4.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i6_LC_13_28_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 pwm_setpoint_i6_LC_13_28_4 (
            .in0(N__50838),
            .in1(N__46224),
            .in2(_gnd_net_),
            .in3(N__47321),
            .lcout(pwm_setpoint_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56238),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i6_3_lut_3_lut_LC_13_28_5.C_ON=1'b0;
    defparam LessThan_299_i6_3_lut_3_lut_LC_13_28_5.SEQ_MODE=4'b0000;
    defparam LessThan_299_i6_3_lut_3_lut_LC_13_28_5.LUT_INIT=16'b1000100011101110;
    LogicCell40 LessThan_299_i6_3_lut_3_lut_LC_13_28_5 (
            .in0(N__46197),
            .in1(N__46185),
            .in2(_gnd_net_),
            .in3(N__48119),
            .lcout(n6_adj_656),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i20_1_lut_LC_13_28_7.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i20_1_lut_LC_13_28_7.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i20_1_lut_LC_13_28_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 unary_minus_13_inv_0_i20_1_lut_LC_13_28_7 (
            .in0(N__46748),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n6_adj_578),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i1_4_lut_LC_13_29_1 .C_ON=1'b0;
    defparam \PWM.i1_4_lut_LC_13_29_1 .SEQ_MODE=4'b0000;
    defparam \PWM.i1_4_lut_LC_13_29_1 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \PWM.i1_4_lut_LC_13_29_1  (
            .in0(N__48526),
            .in1(N__48394),
            .in2(N__47977),
            .in3(N__46728),
            .lcout(\PWM.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_80_LC_13_29_2.C_ON=1'b0;
    defparam i1_4_lut_adj_80_LC_13_29_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_80_LC_13_29_2.LUT_INIT=16'b0111101111011110;
    LogicCell40 i1_4_lut_adj_80_LC_13_29_2 (
            .in0(N__47013),
            .in1(N__56320),
            .in2(N__56405),
            .in3(N__46671),
            .lcout(n4_adj_599),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam commutation_state_prev_i1_LC_13_29_3.C_ON=1'b0;
    defparam commutation_state_prev_i1_LC_13_29_3.SEQ_MODE=4'b1000;
    defparam commutation_state_prev_i1_LC_13_29_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 commutation_state_prev_i1_LC_13_29_3 (
            .in0(N__56322),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(commutation_state_prev_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56245),
            .ce(),
            .sr(_gnd_net_));
    defparam i12529_4_lut_LC_13_29_4.C_ON=1'b0;
    defparam i12529_4_lut_LC_13_29_4.SEQ_MODE=4'b0000;
    defparam i12529_4_lut_LC_13_29_4.LUT_INIT=16'b1000101110111011;
    LogicCell40 i12529_4_lut_LC_13_29_4 (
            .in0(N__46664),
            .in1(N__46622),
            .in2(N__56406),
            .in3(N__56321),
            .lcout(n5201),
            .ltout(n5201_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3271_2_lut_LC_13_29_5.C_ON=1'b0;
    defparam i3271_2_lut_LC_13_29_5.SEQ_MODE=4'b0000;
    defparam i3271_2_lut_LC_13_29_5.LUT_INIT=16'b1010000010100000;
    LogicCell40 i3271_2_lut_LC_13_29_5 (
            .in0(N__46623),
            .in1(_gnd_net_),
            .in2(N__46578),
            .in3(_gnd_net_),
            .lcout(n5253),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i27_2_lut_LC_13_29_6.C_ON=1'b0;
    defparam LessThan_299_i27_2_lut_LC_13_29_6.SEQ_MODE=4'b0000;
    defparam LessThan_299_i27_2_lut_LC_13_29_6.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i27_2_lut_LC_13_29_6 (
            .in0(_gnd_net_),
            .in1(N__46571),
            .in2(_gnd_net_),
            .in3(N__48289),
            .lcout(n27_adj_671),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i11_4_lut_LC_13_29_7 .C_ON=1'b0;
    defparam \PWM.i11_4_lut_LC_13_29_7 .SEQ_MODE=4'b0000;
    defparam \PWM.i11_4_lut_LC_13_29_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \PWM.i11_4_lut_LC_13_29_7  (
            .in0(N__48345),
            .in1(N__48367),
            .in2(N__48270),
            .in3(N__48499),
            .lcout(\PWM.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i12_4_lut_LC_13_30_0 .C_ON=1'b0;
    defparam \PWM.i12_4_lut_LC_13_30_0 .SEQ_MODE=4'b0000;
    defparam \PWM.i12_4_lut_LC_13_30_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \PWM.i12_4_lut_LC_13_30_0  (
            .in0(N__50980),
            .in1(N__48291),
            .in2(N__48210),
            .in3(N__48577),
            .lcout(\PWM.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i10_4_lut_LC_13_30_2 .C_ON=1'b0;
    defparam \PWM.i10_4_lut_LC_13_30_2 .SEQ_MODE=4'b0000;
    defparam \PWM.i10_4_lut_LC_13_30_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \PWM.i10_4_lut_LC_13_30_2  (
            .in0(N__48427),
            .in1(N__48550),
            .in2(N__48243),
            .in3(N__48462),
            .lcout(),
            .ltout(\PWM.n26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i13_4_lut_LC_13_30_3 .C_ON=1'b0;
    defparam \PWM.i13_4_lut_LC_13_30_3 .SEQ_MODE=4'b0000;
    defparam \PWM.i13_4_lut_LC_13_30_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \PWM.i13_4_lut_LC_13_30_3  (
            .in0(N__48314),
            .in1(N__47037),
            .in2(N__47031),
            .in3(N__50934),
            .lcout(),
            .ltout(\PWM.n29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.i9630_4_lut_LC_13_30_4 .C_ON=1'b0;
    defparam \PWM.i9630_4_lut_LC_13_30_4 .SEQ_MODE=4'b0000;
    defparam \PWM.i9630_4_lut_LC_13_30_4 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \PWM.i9630_4_lut_LC_13_30_4  (
            .in0(N__47028),
            .in1(N__50951),
            .in2(N__47022),
            .in3(N__47019),
            .lcout(\PWM.pwm_counter_31__N_407 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam commutation_state_i2_LC_13_30_5.C_ON=1'b0;
    defparam commutation_state_i2_LC_13_30_5.SEQ_MODE=4'b1000;
    defparam commutation_state_i2_LC_13_30_5.LUT_INIT=16'b1000111100000100;
    LogicCell40 commutation_state_i2_LC_13_30_5 (
            .in0(N__47007),
            .in1(N__56404),
            .in2(N__46904),
            .in3(N__46959),
            .lcout(commutation_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56251),
            .ce(),
            .sr(_gnd_net_));
    defparam commutation_state_prev_i2_LC_13_30_6.C_ON=1'b0;
    defparam commutation_state_prev_i2_LC_13_30_6.SEQ_MODE=4'b1000;
    defparam commutation_state_prev_i2_LC_13_30_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 commutation_state_prev_i2_LC_13_30_6 (
            .in0(N__56403),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(commutation_state_prev_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56251),
            .ce(),
            .sr(_gnd_net_));
    defparam commutation_state_i0_LC_13_31_0.C_ON=1'b0;
    defparam commutation_state_i0_LC_13_31_0.SEQ_MODE=4'b1001;
    defparam commutation_state_i0_LC_13_31_0.LUT_INIT=16'b0001000100100010;
    LogicCell40 commutation_state_i0_LC_13_31_0 (
            .in0(N__47006),
            .in1(N__46958),
            .in2(_gnd_net_),
            .in3(N__46903),
            .lcout(commutation_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56255),
            .ce(N__46845),
            .sr(N__46836));
    defparam LessThan_299_i11_2_lut_LC_13_31_1.C_ON=1'b0;
    defparam LessThan_299_i11_2_lut_LC_13_31_1.SEQ_MODE=4'b0000;
    defparam LessThan_299_i11_2_lut_LC_13_31_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 LessThan_299_i11_2_lut_LC_13_31_1 (
            .in0(_gnd_net_),
            .in1(N__46829),
            .in2(_gnd_net_),
            .in3(N__48081),
            .lcout(n11_adj_660),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i29_2_lut_LC_13_31_3.C_ON=1'b0;
    defparam LessThan_299_i29_2_lut_LC_13_31_3.SEQ_MODE=4'b0000;
    defparam LessThan_299_i29_2_lut_LC_13_31_3.LUT_INIT=16'b0101010110101010;
    LogicCell40 LessThan_299_i29_2_lut_LC_13_31_3 (
            .in0(N__48266),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46788),
            .lcout(n29_adj_672),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_13_32_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_13_32_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_13_32_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_13_32_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LessThan_299_i21_2_lut_LC_13_32_6.C_ON=1'b0;
    defparam LessThan_299_i21_2_lut_LC_13_32_6.SEQ_MODE=4'b0000;
    defparam LessThan_299_i21_2_lut_LC_13_32_6.LUT_INIT=16'b0101010110101010;
    LogicCell40 LessThan_299_i21_2_lut_LC_13_32_6 (
            .in0(N__48369),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47117),
            .lcout(n21_adj_667),
            .ltout(n21_adj_667_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12473_3_lut_LC_13_32_7.C_ON=1'b0;
    defparam i12473_3_lut_LC_13_32_7.SEQ_MODE=4'b0000;
    defparam i12473_3_lut_LC_13_32_7.LUT_INIT=16'b1010111110100000;
    LogicCell40 i12473_3_lut_LC_13_32_7 (
            .in0(N__47118),
            .in1(_gnd_net_),
            .in2(N__47106),
            .in3(N__47103),
            .lcout(n15203),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1039_3_lut_LC_14_17_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1039_3_lut_LC_14_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1039_3_lut_LC_14_17_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i1039_3_lut_LC_14_17_0 (
            .in0(_gnd_net_),
            .in1(N__51905),
            .in2(N__48884),
            .in3(N__51891),
            .lcout(n1623_adj_603),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1045_3_lut_LC_14_17_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1045_3_lut_LC_14_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1045_3_lut_LC_14_17_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1045_3_lut_LC_14_17_1 (
            .in0(_gnd_net_),
            .in1(N__52125),
            .in2(N__52149),
            .in3(N__48861),
            .lcout(n1629_adj_609),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_112_LC_14_17_3.C_ON=1'b0;
    defparam i1_2_lut_adj_112_LC_14_17_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_112_LC_14_17_3.LUT_INIT=16'b1111111111110000;
    LogicCell40 i1_2_lut_adj_112_LC_14_17_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__52075),
            .in3(N__52027),
            .lcout(),
            .ltout(n14420_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_118_LC_14_17_4.C_ON=1'b0;
    defparam i1_4_lut_adj_118_LC_14_17_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_118_LC_14_17_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_118_LC_14_17_4 (
            .in0(N__51985),
            .in1(N__51943),
            .in2(N__47085),
            .in3(N__51904),
            .lcout(n14426),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1046_3_lut_LC_14_17_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1046_3_lut_LC_14_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1046_3_lut_LC_14_17_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1046_3_lut_LC_14_17_5 (
            .in0(_gnd_net_),
            .in1(N__51573),
            .in2(N__51594),
            .in3(N__48862),
            .lcout(n1630_adj_610),
            .ltout(n1630_adj_610_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_123_LC_14_17_6.C_ON=1'b0;
    defparam i1_4_lut_adj_123_LC_14_17_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_123_LC_14_17_6.LUT_INIT=16'b1100000010000000;
    LogicCell40 i1_4_lut_adj_123_LC_14_17_6 (
            .in0(N__48913),
            .in1(N__47056),
            .in2(N__47040),
            .in3(N__48726),
            .lcout(n13748),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1049_3_lut_LC_14_17_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1049_3_lut_LC_14_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1049_3_lut_LC_14_17_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i1049_3_lut_LC_14_17_7 (
            .in0(N__51678),
            .in1(N__51710),
            .in2(_gnd_net_),
            .in3(N__48860),
            .lcout(n1633_adj_613),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1040_3_lut_LC_14_18_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1040_3_lut_LC_14_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1040_3_lut_LC_14_18_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1040_3_lut_LC_14_18_0 (
            .in0(_gnd_net_),
            .in1(N__51927),
            .in2(N__51953),
            .in3(N__48875),
            .lcout(n1624_adj_604),
            .ltout(n1624_adj_604_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_124_LC_14_18_1.C_ON=1'b0;
    defparam i1_4_lut_adj_124_LC_14_18_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_124_LC_14_18_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_124_LC_14_18_1 (
            .in0(N__47259),
            .in1(N__47245),
            .in2(N__47229),
            .in3(N__47226),
            .lcout(n14508),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12477_3_lut_LC_14_18_2.C_ON=1'b0;
    defparam i12477_3_lut_LC_14_18_2.SEQ_MODE=4'b0000;
    defparam i12477_3_lut_LC_14_18_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 i12477_3_lut_LC_14_18_2 (
            .in0(_gnd_net_),
            .in1(N__52050),
            .in2(N__52077),
            .in3(N__48874),
            .lcout(n1627_adj_607),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i971_3_lut_LC_14_18_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i971_3_lut_LC_14_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i971_3_lut_LC_14_18_3.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i971_3_lut_LC_14_18_3 (
            .in0(N__51804),
            .in1(_gnd_net_),
            .in2(N__51834),
            .in3(N__48993),
            .lcout(n1523),
            .ltout(n1523_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1038_3_lut_LC_14_18_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1038_3_lut_LC_14_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1038_3_lut_LC_14_18_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1038_3_lut_LC_14_18_4 (
            .in0(_gnd_net_),
            .in1(N__52554),
            .in2(N__47184),
            .in3(N__48876),
            .lcout(n1622_adj_602),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_119_LC_14_18_5.C_ON=1'b0;
    defparam i1_4_lut_adj_119_LC_14_18_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_119_LC_14_18_5.LUT_INIT=16'b1111111110000000;
    LogicCell40 i1_4_lut_adj_119_LC_14_18_5 (
            .in0(N__52141),
            .in1(N__52105),
            .in2(N__49023),
            .in3(N__47157),
            .lcout(),
            .ltout(n14428_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12864_4_lut_LC_14_18_6.C_ON=1'b0;
    defparam i12864_4_lut_LC_14_18_6.SEQ_MODE=4'b0000;
    defparam i12864_4_lut_LC_14_18_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12864_4_lut_LC_14_18_6 (
            .in0(N__52525),
            .in1(N__51866),
            .in2(N__47151),
            .in3(N__52496),
            .lcout(n1554),
            .ltout(n1554_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12861_1_lut_LC_14_18_7.C_ON=1'b0;
    defparam i12861_1_lut_LC_14_18_7.SEQ_MODE=4'b0000;
    defparam i12861_1_lut_LC_14_18_7.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12861_1_lut_LC_14_18_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47148),
            .in3(_gnd_net_),
            .lcout(n15591),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i908_3_lut_LC_14_19_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i908_3_lut_LC_14_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i908_3_lut_LC_14_19_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i908_3_lut_LC_14_19_0 (
            .in0(_gnd_net_),
            .in1(N__47445),
            .in2(N__49188),
            .in3(N__52332),
            .lcout(n1428),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i907_3_lut_LC_14_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i907_3_lut_LC_14_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i907_3_lut_LC_14_19_1.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i907_3_lut_LC_14_19_1 (
            .in0(_gnd_net_),
            .in1(N__49287),
            .in2(N__52348),
            .in3(N__47436),
            .lcout(n1427),
            .ltout(n1427_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_107_LC_14_19_2.C_ON=1'b0;
    defparam i1_2_lut_adj_107_LC_14_19_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_107_LC_14_19_2.LUT_INIT=16'b1111111111110000;
    LogicCell40 i1_2_lut_adj_107_LC_14_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47409),
            .in3(N__51388),
            .lcout(n14484),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1044_rep_29_3_lut_LC_14_19_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1044_rep_29_3_lut_LC_14_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1044_rep_29_3_lut_LC_14_19_3.LUT_INIT=16'b1010110010101100;
    LogicCell40 encoder0_position_31__I_0_i1044_rep_29_3_lut_LC_14_19_3 (
            .in0(N__52109),
            .in1(N__52089),
            .in2(N__48886),
            .in3(_gnd_net_),
            .lcout(n1628_adj_608),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i904_3_lut_LC_14_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i904_3_lut_LC_14_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i904_3_lut_LC_14_19_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i904_3_lut_LC_14_19_4 (
            .in0(_gnd_net_),
            .in1(N__47421),
            .in2(N__49668),
            .in3(N__52336),
            .lcout(n1424),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i23_3_lut_LC_14_19_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i23_3_lut_LC_14_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i23_3_lut_LC_14_19_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i23_3_lut_LC_14_19_5 (
            .in0(N__47385),
            .in1(N__49606),
            .in2(_gnd_net_),
            .in3(N__47370),
            .lcout(n297),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1042_3_lut_LC_14_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1042_3_lut_LC_14_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1042_3_lut_LC_14_19_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i1042_3_lut_LC_14_19_6 (
            .in0(_gnd_net_),
            .in1(N__52011),
            .in2(N__52035),
            .in3(N__48870),
            .lcout(n1626_adj_606),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i7_1_lut_LC_14_19_7.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i7_1_lut_LC_14_19_7.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i7_1_lut_LC_14_19_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i7_1_lut_LC_14_19_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47322),
            .lcout(n19_adj_591),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_2_lut_LC_14_20_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_2_lut_LC_14_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_2_lut_LC_14_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_2_lut_LC_14_20_0 (
            .in0(_gnd_net_),
            .in1(N__49138),
            .in2(_gnd_net_),
            .in3(N__47289),
            .lcout(n1401),
            .ltout(),
            .carryin(bfn_14_20_0_),
            .carryout(n12541),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_3_lut_LC_14_20_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_3_lut_LC_14_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_3_lut_LC_14_20_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_3_lut_LC_14_20_1 (
            .in0(_gnd_net_),
            .in1(N__54890),
            .in2(N__49080),
            .in3(N__47286),
            .lcout(n1400),
            .ltout(),
            .carryin(n12541),
            .carryout(n12542),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_4_lut_LC_14_20_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_4_lut_LC_14_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_4_lut_LC_14_20_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_4_lut_LC_14_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__49212),
            .in3(N__47454),
            .lcout(n1399),
            .ltout(),
            .carryin(n12542),
            .carryout(n12543),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_5_lut_LC_14_20_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_5_lut_LC_14_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_5_lut_LC_14_20_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_5_lut_LC_14_20_3 (
            .in0(_gnd_net_),
            .in1(N__54891),
            .in2(N__49233),
            .in3(N__47451),
            .lcout(n1398),
            .ltout(),
            .carryin(n12543),
            .carryout(n12544),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_6_lut_LC_14_20_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_6_lut_LC_14_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_6_lut_LC_14_20_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_6_lut_LC_14_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__53121),
            .in3(N__47448),
            .lcout(n1397),
            .ltout(),
            .carryin(n12544),
            .carryout(n12545),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_7_lut_LC_14_20_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_7_lut_LC_14_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_7_lut_LC_14_20_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_7_lut_LC_14_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__49184),
            .in3(N__47439),
            .lcout(n1396),
            .ltout(),
            .carryin(n12545),
            .carryout(n12546),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_8_lut_LC_14_20_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_8_lut_LC_14_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_8_lut_LC_14_20_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_8_lut_LC_14_20_6 (
            .in0(_gnd_net_),
            .in1(N__54893),
            .in2(N__49286),
            .in3(N__47430),
            .lcout(n1395),
            .ltout(),
            .carryin(n12546),
            .carryout(n12547),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_9_lut_LC_14_20_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_9_lut_LC_14_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_9_lut_LC_14_20_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_9_lut_LC_14_20_7 (
            .in0(_gnd_net_),
            .in1(N__54892),
            .in2(N__49256),
            .in3(N__47427),
            .lcout(n1394),
            .ltout(),
            .carryin(n12547),
            .carryout(n12548),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_10_lut_LC_14_21_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_10_lut_LC_14_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_10_lut_LC_14_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_10_lut_LC_14_21_0 (
            .in0(_gnd_net_),
            .in1(N__54661),
            .in2(N__49376),
            .in3(N__47424),
            .lcout(n1393),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(n12549),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_11_lut_LC_14_21_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_11_lut_LC_14_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_11_lut_LC_14_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_11_lut_LC_14_21_1 (
            .in0(_gnd_net_),
            .in1(N__54657),
            .in2(N__49664),
            .in3(N__47412),
            .lcout(n1392),
            .ltout(),
            .carryin(n12549),
            .carryout(n12550),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_12_lut_LC_14_21_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_900_12_lut_LC_14_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_12_lut_LC_14_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_900_12_lut_LC_14_21_2 (
            .in0(_gnd_net_),
            .in1(N__50001),
            .in2(N__54952),
            .in3(N__47508),
            .lcout(n1391),
            .ltout(),
            .carryin(n12550),
            .carryout(n12551),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_900_13_lut_LC_14_21_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_900_13_lut_LC_14_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_900_13_lut_LC_14_21_3.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_900_13_lut_LC_14_21_3 (
            .in0(N__54662),
            .in1(N__47489),
            .in2(N__52581),
            .in3(N__47505),
            .lcout(n1422),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12823_1_lut_LC_14_21_4.C_ON=1'b0;
    defparam i12823_1_lut_LC_14_21_4.SEQ_MODE=4'b0000;
    defparam i12823_1_lut_LC_14_21_4.LUT_INIT=16'b0000111100001111;
    LogicCell40 i12823_1_lut_LC_14_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__52347),
            .in3(_gnd_net_),
            .lcout(n15553),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i774_3_lut_LC_14_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i774_3_lut_LC_14_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i774_3_lut_LC_14_21_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i774_3_lut_LC_14_21_5 (
            .in0(_gnd_net_),
            .in1(N__47556),
            .in2(N__47580),
            .in3(N__49934),
            .lcout(n1230),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i845_3_lut_LC_14_21_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i845_3_lut_LC_14_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i845_3_lut_LC_14_21_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i845_3_lut_LC_14_21_6 (
            .in0(N__52230),
            .in1(N__52248),
            .in2(_gnd_net_),
            .in3(N__53174),
            .lcout(n1333),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i913_3_lut_LC_14_21_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i913_3_lut_LC_14_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i913_3_lut_LC_14_21_7.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_i913_3_lut_LC_14_21_7 (
            .in0(N__49139),
            .in1(_gnd_net_),
            .in2(N__47478),
            .in3(N__52327),
            .lcout(n1433),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_96_LC_14_22_0.C_ON=1'b0;
    defparam i1_3_lut_adj_96_LC_14_22_0.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_96_LC_14_22_0.LUT_INIT=16'b1111111111111010;
    LogicCell40 i1_3_lut_adj_96_LC_14_22_0 (
            .in0(N__49307),
            .in1(_gnd_net_),
            .in2(N__49805),
            .in3(N__50026),
            .lcout(),
            .ltout(n14406_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12795_4_lut_LC_14_22_1.C_ON=1'b0;
    defparam i12795_4_lut_LC_14_22_1.SEQ_MODE=4'b0000;
    defparam i12795_4_lut_LC_14_22_1.LUT_INIT=16'b0000000100000011;
    LogicCell40 i12795_4_lut_LC_14_22_1 (
            .in0(N__47469),
            .in1(N__47681),
            .in2(N__47463),
            .in3(N__47460),
            .lcout(n1158),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i773_3_lut_LC_14_22_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i773_3_lut_LC_14_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i773_3_lut_LC_14_22_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i773_3_lut_LC_14_22_2 (
            .in0(_gnd_net_),
            .in1(N__47520),
            .in2(N__47544),
            .in3(N__49924),
            .lcout(n1229),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12765_2_lut_LC_14_22_3.C_ON=1'b0;
    defparam i12765_2_lut_LC_14_22_3.SEQ_MODE=4'b0000;
    defparam i12765_2_lut_LC_14_22_3.LUT_INIT=16'b0000000011001100;
    LogicCell40 i12765_2_lut_LC_14_22_3 (
            .in0(_gnd_net_),
            .in1(N__55761),
            .in2(_gnd_net_),
            .in3(N__47661),
            .lcout(n5215),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i776_3_lut_LC_14_22_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i776_3_lut_LC_14_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i776_3_lut_LC_14_22_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i776_3_lut_LC_14_22_4 (
            .in0(_gnd_net_),
            .in1(N__47615),
            .in2(N__47595),
            .in3(N__49923),
            .lcout(n1232),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i777_3_lut_LC_14_22_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i777_3_lut_LC_14_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i777_3_lut_LC_14_22_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 encoder0_position_31__I_0_i777_3_lut_LC_14_22_6 (
            .in0(N__47625),
            .in1(N__47649),
            .in2(_gnd_net_),
            .in3(N__49922),
            .lcout(n1233),
            .ltout(n1233_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9951_3_lut_LC_14_22_7.C_ON=1'b0;
    defparam i9951_3_lut_LC_14_22_7.SEQ_MODE=4'b0000;
    defparam i9951_3_lut_LC_14_22_7.LUT_INIT=16'b1111101000000000;
    LogicCell40 i9951_3_lut_LC_14_22_7 (
            .in0(N__52246),
            .in1(_gnd_net_),
            .in2(N__47652),
            .in3(N__52177),
            .lcout(n11927),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_2_lut_LC_14_23_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_2_lut_LC_14_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_2_lut_LC_14_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_2_lut_LC_14_23_0 (
            .in0(_gnd_net_),
            .in1(N__47648),
            .in2(_gnd_net_),
            .in3(N__47619),
            .lcout(n1201),
            .ltout(),
            .carryin(bfn_14_23_0_),
            .carryout(n12522),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_3_lut_LC_14_23_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_3_lut_LC_14_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_3_lut_LC_14_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_3_lut_LC_14_23_1 (
            .in0(_gnd_net_),
            .in1(N__54247),
            .in2(N__47616),
            .in3(N__47586),
            .lcout(n1200),
            .ltout(),
            .carryin(n12522),
            .carryout(n12523),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_4_lut_LC_14_23_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_4_lut_LC_14_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_4_lut_LC_14_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_4_lut_LC_14_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__49328),
            .in3(N__47583),
            .lcout(n1199),
            .ltout(),
            .carryin(n12523),
            .carryout(n12524),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_5_lut_LC_14_23_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_5_lut_LC_14_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_5_lut_LC_14_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_5_lut_LC_14_23_3 (
            .in0(_gnd_net_),
            .in1(N__54248),
            .in2(N__47579),
            .in3(N__47547),
            .lcout(n1198),
            .ltout(),
            .carryin(n12524),
            .carryout(n12525),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_6_lut_LC_14_23_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_6_lut_LC_14_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_6_lut_LC_14_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_6_lut_LC_14_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__47543),
            .in3(N__47514),
            .lcout(n1197),
            .ltout(),
            .carryin(n12525),
            .carryout(n12526),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_7_lut_LC_14_23_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_7_lut_LC_14_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_7_lut_LC_14_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_7_lut_LC_14_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__49979),
            .in3(N__47511),
            .lcout(n1196),
            .ltout(),
            .carryin(n12526),
            .carryout(n12527),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_8_lut_LC_14_23_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_8_lut_LC_14_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_8_lut_LC_14_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_8_lut_LC_14_23_6 (
            .in0(_gnd_net_),
            .in1(N__49801),
            .in2(N__54656),
            .in3(N__47757),
            .lcout(n1195),
            .ltout(),
            .carryin(n12527),
            .carryout(n12528),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_9_lut_LC_14_23_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_9_lut_LC_14_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_9_lut_LC_14_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_9_lut_LC_14_23_7 (
            .in0(_gnd_net_),
            .in1(N__54252),
            .in2(N__49311),
            .in3(N__47754),
            .lcout(n1194),
            .ltout(),
            .carryin(n12528),
            .carryout(n12529),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_10_lut_LC_14_24_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_766_10_lut_LC_14_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_10_lut_LC_14_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_766_10_lut_LC_14_24_0 (
            .in0(_gnd_net_),
            .in1(N__53789),
            .in2(N__50033),
            .in3(N__47751),
            .lcout(n1193),
            .ltout(),
            .carryin(bfn_14_24_0_),
            .carryout(n12530),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_766_11_lut_LC_14_24_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_766_11_lut_LC_14_24_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_766_11_lut_LC_14_24_1.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_766_11_lut_LC_14_24_1 (
            .in0(N__53790),
            .in1(N__47738),
            .in2(N__47682),
            .in3(N__47748),
            .lcout(n1224),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12792_1_lut_LC_14_24_3.C_ON=1'b0;
    defparam i12792_1_lut_LC_14_24_3.SEQ_MODE=4'b0000;
    defparam i12792_1_lut_LC_14_24_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12792_1_lut_LC_14_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49941),
            .lcout(n15522),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i21_3_lut_LC_14_24_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i21_3_lut_LC_14_24_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i21_3_lut_LC_14_24_4.LUT_INIT=16'b1010101011110000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i21_3_lut_LC_14_24_4 (
            .in0(N__47727),
            .in1(_gnd_net_),
            .in2(N__47715),
            .in3(N__49603),
            .lcout(n299),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i701_3_lut_LC_14_24_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i701_3_lut_LC_14_24_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i701_3_lut_LC_14_24_6.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i701_3_lut_LC_14_24_6 (
            .in0(_gnd_net_),
            .in1(N__49854),
            .in2(N__53384),
            .in3(N__53355),
            .lcout(n1125),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_3_lut_LC_14_25_2.C_ON=1'b0;
    defparam i7_3_lut_LC_14_25_2.SEQ_MODE=4'b0000;
    defparam i7_3_lut_LC_14_25_2.LUT_INIT=16'b1111111111101110;
    LogicCell40 i7_3_lut_LC_14_25_2 (
            .in0(N__53346),
            .in1(N__55716),
            .in2(_gnd_net_),
            .in3(N__53328),
            .lcout(),
            .ltout(n20_adj_618_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12_4_lut_LC_14_25_3.C_ON=1'b0;
    defparam i12_4_lut_LC_14_25_3.SEQ_MODE=4'b0000;
    defparam i12_4_lut_LC_14_25_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12_4_lut_LC_14_25_3 (
            .in0(N__55629),
            .in1(N__53247),
            .in2(N__47664),
            .in3(N__47904),
            .lcout(n13197),
            .ltout(n13197_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam direction_167_LC_14_25_4.C_ON=1'b0;
    defparam direction_167_LC_14_25_4.SEQ_MODE=4'b1000;
    defparam direction_167_LC_14_25_4.LUT_INIT=16'b1100110011000110;
    LogicCell40 direction_167_LC_14_25_4 (
            .in0(N__55760),
            .in1(N__51117),
            .in2(N__47823),
            .in3(N__47805),
            .lcout(direction_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56228),
            .ce(),
            .sr(_gnd_net_));
    defparam i9624_4_lut_LC_14_25_5.C_ON=1'b0;
    defparam i9624_4_lut_LC_14_25_5.SEQ_MODE=4'b0000;
    defparam i9624_4_lut_LC_14_25_5.LUT_INIT=16'b1000111100001111;
    LogicCell40 i9624_4_lut_LC_14_25_5 (
            .in0(N__47820),
            .in1(N__47772),
            .in2(N__51049),
            .in3(N__47919),
            .lcout(direction_N_342),
            .ltout(direction_N_342_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_303_i1_3_lut_LC_14_25_6.C_ON=1'b0;
    defparam mux_303_i1_3_lut_LC_14_25_6.SEQ_MODE=4'b0000;
    defparam mux_303_i1_3_lut_LC_14_25_6.LUT_INIT=16'b0000111111001100;
    LogicCell40 mux_303_i1_3_lut_LC_14_25_6 (
            .in0(_gnd_net_),
            .in1(N__47789),
            .in2(N__47814),
            .in3(N__51115),
            .lcout(n1693),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i20_3_lut_LC_14_25_7.C_ON=1'b0;
    defparam i20_3_lut_LC_14_25_7.SEQ_MODE=4'b0000;
    defparam i20_3_lut_LC_14_25_7.LUT_INIT=16'b1110111001000100;
    LogicCell40 i20_3_lut_LC_14_25_7 (
            .in0(N__51116),
            .in1(N__47790),
            .in2(_gnd_net_),
            .in3(N__47811),
            .lcout(n13675),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9_4_lut_adj_72_LC_14_26_0.C_ON=1'b0;
    defparam i9_4_lut_adj_72_LC_14_26_0.SEQ_MODE=4'b0000;
    defparam i9_4_lut_adj_72_LC_14_26_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i9_4_lut_adj_72_LC_14_26_0 (
            .in0(N__50586),
            .in1(N__50418),
            .in2(N__50510),
            .in3(N__50544),
            .lcout(),
            .ltout(n23_adj_709_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i831_4_lut_LC_14_26_1.C_ON=1'b0;
    defparam i831_4_lut_LC_14_26_1.SEQ_MODE=4'b0000;
    defparam i831_4_lut_LC_14_26_1.LUT_INIT=16'b1010101010101011;
    LogicCell40 i831_4_lut_LC_14_26_1 (
            .in0(N__51039),
            .in1(N__47778),
            .in2(N__47799),
            .in3(N__47796),
            .lcout(direction_N_340),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_adj_71_LC_14_26_2.C_ON=1'b0;
    defparam i10_4_lut_adj_71_LC_14_26_2.SEQ_MODE=4'b0000;
    defparam i10_4_lut_adj_71_LC_14_26_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i10_4_lut_adj_71_LC_14_26_2 (
            .in0(N__51038),
            .in1(N__50463),
            .in2(N__50705),
            .in3(N__51291),
            .lcout(n24_adj_708),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9_4_lut_LC_14_26_3.C_ON=1'b0;
    defparam i9_4_lut_LC_14_26_3.SEQ_MODE=4'b0000;
    defparam i9_4_lut_LC_14_26_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 i9_4_lut_LC_14_26_3 (
            .in0(N__50625),
            .in1(N__50419),
            .in2(N__50676),
            .in3(N__50587),
            .lcout(n23_adj_654),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_setpoint_i1_LC_14_26_5.C_ON=1'b0;
    defparam pwm_setpoint_i1_LC_14_26_5.SEQ_MODE=4'b1000;
    defparam pwm_setpoint_i1_LC_14_26_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 pwm_setpoint_i1_LC_14_26_5 (
            .in0(N__50905),
            .in1(N__47766),
            .in2(_gnd_net_),
            .in3(N__47874),
            .lcout(pwm_setpoint_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56233),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_LC_14_26_6.C_ON=1'b0;
    defparam i2_2_lut_LC_14_26_6.SEQ_MODE=4'b0000;
    defparam i2_2_lut_LC_14_26_6.LUT_INIT=16'b1000100010001000;
    LogicCell40 i2_2_lut_LC_14_26_6 (
            .in0(N__50700),
            .in1(N__51216),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(n16_adj_679_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11_4_lut_LC_14_26_7.C_ON=1'b0;
    defparam i11_4_lut_LC_14_26_7.SEQ_MODE=4'b0000;
    defparam i11_4_lut_LC_14_26_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 i11_4_lut_LC_14_26_7 (
            .in0(N__51292),
            .in1(N__50505),
            .in2(N__47928),
            .in3(N__47925),
            .lcout(n25_adj_652),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9_4_lut_adj_76_LC_14_27_0.C_ON=1'b0;
    defparam i9_4_lut_adj_76_LC_14_27_0.SEQ_MODE=4'b0000;
    defparam i9_4_lut_adj_76_LC_14_27_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i9_4_lut_adj_76_LC_14_27_0 (
            .in0(N__53310),
            .in1(N__53289),
            .in2(N__55674),
            .in3(N__55938),
            .lcout(n22_adj_617),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_2_lut_LC_14_27_1.C_ON=1'b0;
    defparam i3_2_lut_LC_14_27_1.SEQ_MODE=4'b0000;
    defparam i3_2_lut_LC_14_27_1.LUT_INIT=16'b1111111111001100;
    LogicCell40 i3_2_lut_LC_14_27_1 (
            .in0(_gnd_net_),
            .in1(N__55650),
            .in2(_gnd_net_),
            .in3(N__55959),
            .lcout(),
            .ltout(n16_adj_619_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11_4_lut_adj_77_LC_14_27_2.C_ON=1'b0;
    defparam i11_4_lut_adj_77_LC_14_27_2.SEQ_MODE=4'b0000;
    defparam i11_4_lut_adj_77_LC_14_27_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i11_4_lut_adj_77_LC_14_27_2 (
            .in0(N__55698),
            .in1(N__53268),
            .in2(N__47913),
            .in3(N__47910),
            .lcout(n24_adj_616),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_23__I_0_204_inv_0_i17_1_lut_LC_14_27_3.C_ON=1'b0;
    defparam encoder0_position_target_23__I_0_204_inv_0_i17_1_lut_LC_14_27_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_target_23__I_0_204_inv_0_i17_1_lut_LC_14_27_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_target_23__I_0_204_inv_0_i17_1_lut_LC_14_27_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47895),
            .lcout(n9_adj_567),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam unary_minus_13_inv_0_i2_1_lut_LC_14_27_4.C_ON=1'b0;
    defparam unary_minus_13_inv_0_i2_1_lut_LC_14_27_4.SEQ_MODE=4'b0000;
    defparam unary_minus_13_inv_0_i2_1_lut_LC_14_27_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 unary_minus_13_inv_0_i2_1_lut_LC_14_27_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47873),
            .lcout(n24_adj_596),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2178_1_lut_LC_14_27_7.C_ON=1'b0;
    defparam i2178_1_lut_LC_14_27_7.SEQ_MODE=4'b0000;
    defparam i2178_1_lut_LC_14_27_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 i2178_1_lut_LC_14_27_7 (
            .in0(N__50863),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(pwm_setpoint_23__N_195),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWM.pwm_counter_664__i0_LC_14_28_0 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i0_LC_14_28_0 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i0_LC_14_28_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i0_LC_14_28_0  (
            .in0(_gnd_net_),
            .in1(N__48173),
            .in2(_gnd_net_),
            .in3(N__48159),
            .lcout(pwm_counter_0),
            .ltout(),
            .carryin(bfn_14_28_0_),
            .carryout(\PWM.n13022 ),
            .clk(N__56246),
            .ce(),
            .sr(N__48702));
    defparam \PWM.pwm_counter_664__i1_LC_14_28_1 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i1_LC_14_28_1 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i1_LC_14_28_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i1_LC_14_28_1  (
            .in0(_gnd_net_),
            .in1(N__48155),
            .in2(_gnd_net_),
            .in3(N__48141),
            .lcout(pwm_counter_1),
            .ltout(),
            .carryin(\PWM.n13022 ),
            .carryout(\PWM.n13023 ),
            .clk(N__56246),
            .ce(),
            .sr(N__48702));
    defparam \PWM.pwm_counter_664__i2_LC_14_28_2 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i2_LC_14_28_2 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i2_LC_14_28_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i2_LC_14_28_2  (
            .in0(_gnd_net_),
            .in1(N__48137),
            .in2(_gnd_net_),
            .in3(N__48123),
            .lcout(pwm_counter_2),
            .ltout(),
            .carryin(\PWM.n13023 ),
            .carryout(\PWM.n13024 ),
            .clk(N__56246),
            .ce(),
            .sr(N__48702));
    defparam \PWM.pwm_counter_664__i3_LC_14_28_3 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i3_LC_14_28_3 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i3_LC_14_28_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i3_LC_14_28_3  (
            .in0(_gnd_net_),
            .in1(N__48120),
            .in2(_gnd_net_),
            .in3(N__48105),
            .lcout(pwm_counter_3),
            .ltout(),
            .carryin(\PWM.n13024 ),
            .carryout(\PWM.n13025 ),
            .clk(N__56246),
            .ce(),
            .sr(N__48702));
    defparam \PWM.pwm_counter_664__i4_LC_14_28_4 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i4_LC_14_28_4 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i4_LC_14_28_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i4_LC_14_28_4  (
            .in0(_gnd_net_),
            .in1(N__48098),
            .in2(_gnd_net_),
            .in3(N__48084),
            .lcout(pwm_counter_4),
            .ltout(),
            .carryin(\PWM.n13025 ),
            .carryout(\PWM.n13026 ),
            .clk(N__56246),
            .ce(),
            .sr(N__48702));
    defparam \PWM.pwm_counter_664__i5_LC_14_28_5 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i5_LC_14_28_5 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i5_LC_14_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i5_LC_14_28_5  (
            .in0(_gnd_net_),
            .in1(N__48079),
            .in2(_gnd_net_),
            .in3(N__48060),
            .lcout(pwm_counter_5),
            .ltout(),
            .carryin(\PWM.n13026 ),
            .carryout(\PWM.n13027 ),
            .clk(N__56246),
            .ce(),
            .sr(N__48702));
    defparam \PWM.pwm_counter_664__i6_LC_14_28_6 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i6_LC_14_28_6 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i6_LC_14_28_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i6_LC_14_28_6  (
            .in0(_gnd_net_),
            .in1(N__48049),
            .in2(_gnd_net_),
            .in3(N__48021),
            .lcout(pwm_counter_6),
            .ltout(),
            .carryin(\PWM.n13027 ),
            .carryout(\PWM.n13028 ),
            .clk(N__56246),
            .ce(),
            .sr(N__48702));
    defparam \PWM.pwm_counter_664__i7_LC_14_28_7 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i7_LC_14_28_7 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i7_LC_14_28_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i7_LC_14_28_7  (
            .in0(_gnd_net_),
            .in1(N__48010),
            .in2(_gnd_net_),
            .in3(N__47982),
            .lcout(pwm_counter_7),
            .ltout(),
            .carryin(\PWM.n13028 ),
            .carryout(\PWM.n13029 ),
            .clk(N__56246),
            .ce(),
            .sr(N__48702));
    defparam \PWM.pwm_counter_664__i8_LC_14_29_0 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i8_LC_14_29_0 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i8_LC_14_29_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i8_LC_14_29_0  (
            .in0(_gnd_net_),
            .in1(N__47967),
            .in2(_gnd_net_),
            .in3(N__47943),
            .lcout(pwm_counter_8),
            .ltout(),
            .carryin(bfn_14_29_0_),
            .carryout(\PWM.n13030 ),
            .clk(N__56252),
            .ce(),
            .sr(N__48694));
    defparam \PWM.pwm_counter_664__i9_LC_14_29_1 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i9_LC_14_29_1 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i9_LC_14_29_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i9_LC_14_29_1  (
            .in0(_gnd_net_),
            .in1(N__48393),
            .in2(_gnd_net_),
            .in3(N__48372),
            .lcout(pwm_counter_9),
            .ltout(),
            .carryin(\PWM.n13030 ),
            .carryout(\PWM.n13031 ),
            .clk(N__56252),
            .ce(),
            .sr(N__48694));
    defparam \PWM.pwm_counter_664__i10_LC_14_29_2 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i10_LC_14_29_2 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i10_LC_14_29_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i10_LC_14_29_2  (
            .in0(_gnd_net_),
            .in1(N__48368),
            .in2(_gnd_net_),
            .in3(N__48348),
            .lcout(pwm_counter_10),
            .ltout(),
            .carryin(\PWM.n13031 ),
            .carryout(\PWM.n13032 ),
            .clk(N__56252),
            .ce(),
            .sr(N__48694));
    defparam \PWM.pwm_counter_664__i11_LC_14_29_3 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i11_LC_14_29_3 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i11_LC_14_29_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i11_LC_14_29_3  (
            .in0(_gnd_net_),
            .in1(N__48340),
            .in2(_gnd_net_),
            .in3(N__48321),
            .lcout(pwm_counter_11),
            .ltout(),
            .carryin(\PWM.n13032 ),
            .carryout(\PWM.n13033 ),
            .clk(N__56252),
            .ce(),
            .sr(N__48694));
    defparam \PWM.pwm_counter_664__i12_LC_14_29_4 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i12_LC_14_29_4 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i12_LC_14_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i12_LC_14_29_4  (
            .in0(_gnd_net_),
            .in1(N__48313),
            .in2(_gnd_net_),
            .in3(N__48294),
            .lcout(pwm_counter_12),
            .ltout(),
            .carryin(\PWM.n13033 ),
            .carryout(\PWM.n13034 ),
            .clk(N__56252),
            .ce(),
            .sr(N__48694));
    defparam \PWM.pwm_counter_664__i13_LC_14_29_5 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i13_LC_14_29_5 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i13_LC_14_29_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i13_LC_14_29_5  (
            .in0(_gnd_net_),
            .in1(N__48290),
            .in2(_gnd_net_),
            .in3(N__48273),
            .lcout(pwm_counter_13),
            .ltout(),
            .carryin(\PWM.n13034 ),
            .carryout(\PWM.n13035 ),
            .clk(N__56252),
            .ce(),
            .sr(N__48694));
    defparam \PWM.pwm_counter_664__i14_LC_14_29_6 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i14_LC_14_29_6 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i14_LC_14_29_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i14_LC_14_29_6  (
            .in0(_gnd_net_),
            .in1(N__48265),
            .in2(_gnd_net_),
            .in3(N__48246),
            .lcout(pwm_counter_14),
            .ltout(),
            .carryin(\PWM.n13035 ),
            .carryout(\PWM.n13036 ),
            .clk(N__56252),
            .ce(),
            .sr(N__48694));
    defparam \PWM.pwm_counter_664__i15_LC_14_29_7 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i15_LC_14_29_7 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i15_LC_14_29_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i15_LC_14_29_7  (
            .in0(_gnd_net_),
            .in1(N__48235),
            .in2(_gnd_net_),
            .in3(N__48216),
            .lcout(pwm_counter_15),
            .ltout(),
            .carryin(\PWM.n13036 ),
            .carryout(\PWM.n13037 ),
            .clk(N__56252),
            .ce(),
            .sr(N__48694));
    defparam \PWM.pwm_counter_664__i16_LC_14_30_0 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i16_LC_14_30_0 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i16_LC_14_30_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i16_LC_14_30_0  (
            .in0(_gnd_net_),
            .in1(N__48202),
            .in2(_gnd_net_),
            .in3(N__48180),
            .lcout(pwm_counter_16),
            .ltout(),
            .carryin(bfn_14_30_0_),
            .carryout(\PWM.n13038 ),
            .clk(N__56256),
            .ce(),
            .sr(N__48693));
    defparam \PWM.pwm_counter_664__i17_LC_14_30_1 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i17_LC_14_30_1 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i17_LC_14_30_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i17_LC_14_30_1  (
            .in0(_gnd_net_),
            .in1(N__48578),
            .in2(_gnd_net_),
            .in3(N__48558),
            .lcout(pwm_counter_17),
            .ltout(),
            .carryin(\PWM.n13038 ),
            .carryout(\PWM.n13039 ),
            .clk(N__56256),
            .ce(),
            .sr(N__48693));
    defparam \PWM.pwm_counter_664__i18_LC_14_30_2 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i18_LC_14_30_2 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i18_LC_14_30_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i18_LC_14_30_2  (
            .in0(_gnd_net_),
            .in1(N__48554),
            .in2(_gnd_net_),
            .in3(N__48531),
            .lcout(pwm_counter_18),
            .ltout(),
            .carryin(\PWM.n13039 ),
            .carryout(\PWM.n13040 ),
            .clk(N__56256),
            .ce(),
            .sr(N__48693));
    defparam \PWM.pwm_counter_664__i19_LC_14_30_3 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i19_LC_14_30_3 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i19_LC_14_30_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i19_LC_14_30_3  (
            .in0(_gnd_net_),
            .in1(N__48527),
            .in2(_gnd_net_),
            .in3(N__48507),
            .lcout(pwm_counter_19),
            .ltout(),
            .carryin(\PWM.n13040 ),
            .carryout(\PWM.n13041 ),
            .clk(N__56256),
            .ce(),
            .sr(N__48693));
    defparam \PWM.pwm_counter_664__i20_LC_14_30_4 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i20_LC_14_30_4 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i20_LC_14_30_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i20_LC_14_30_4  (
            .in0(_gnd_net_),
            .in1(N__48500),
            .in2(_gnd_net_),
            .in3(N__48480),
            .lcout(pwm_counter_20),
            .ltout(),
            .carryin(\PWM.n13041 ),
            .carryout(\PWM.n13042 ),
            .clk(N__56256),
            .ce(),
            .sr(N__48693));
    defparam \PWM.pwm_counter_664__i21_LC_14_30_5 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i21_LC_14_30_5 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i21_LC_14_30_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i21_LC_14_30_5  (
            .in0(_gnd_net_),
            .in1(N__48463),
            .in2(_gnd_net_),
            .in3(N__48435),
            .lcout(pwm_counter_21),
            .ltout(),
            .carryin(\PWM.n13042 ),
            .carryout(\PWM.n13043 ),
            .clk(N__56256),
            .ce(),
            .sr(N__48693));
    defparam \PWM.pwm_counter_664__i22_LC_14_30_6 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i22_LC_14_30_6 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i22_LC_14_30_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i22_LC_14_30_6  (
            .in0(_gnd_net_),
            .in1(N__48428),
            .in2(_gnd_net_),
            .in3(N__48408),
            .lcout(pwm_counter_22),
            .ltout(),
            .carryin(\PWM.n13043 ),
            .carryout(\PWM.n13044 ),
            .clk(N__56256),
            .ce(),
            .sr(N__48693));
    defparam \PWM.pwm_counter_664__i23_LC_14_30_7 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i23_LC_14_30_7 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i23_LC_14_30_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i23_LC_14_30_7  (
            .in0(_gnd_net_),
            .in1(N__50981),
            .in2(_gnd_net_),
            .in3(N__48405),
            .lcout(pwm_counter_23),
            .ltout(),
            .carryin(\PWM.n13044 ),
            .carryout(\PWM.n13045 ),
            .clk(N__56256),
            .ce(),
            .sr(N__48693));
    defparam \PWM.pwm_counter_664__i24_LC_14_31_0 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i24_LC_14_31_0 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i24_LC_14_31_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i24_LC_14_31_0  (
            .in0(_gnd_net_),
            .in1(N__48672),
            .in2(_gnd_net_),
            .in3(N__48402),
            .lcout(pwm_counter_24),
            .ltout(),
            .carryin(bfn_14_31_0_),
            .carryout(\PWM.n13046 ),
            .clk(N__56257),
            .ce(),
            .sr(N__48695));
    defparam \PWM.pwm_counter_664__i25_LC_14_31_1 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i25_LC_14_31_1 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i25_LC_14_31_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i25_LC_14_31_1  (
            .in0(_gnd_net_),
            .in1(N__48609),
            .in2(_gnd_net_),
            .in3(N__48399),
            .lcout(pwm_counter_25),
            .ltout(),
            .carryin(\PWM.n13046 ),
            .carryout(\PWM.n13047 ),
            .clk(N__56257),
            .ce(),
            .sr(N__48695));
    defparam \PWM.pwm_counter_664__i26_LC_14_31_2 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i26_LC_14_31_2 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i26_LC_14_31_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i26_LC_14_31_2  (
            .in0(_gnd_net_),
            .in1(N__48633),
            .in2(_gnd_net_),
            .in3(N__48720),
            .lcout(pwm_counter_26),
            .ltout(),
            .carryin(\PWM.n13047 ),
            .carryout(\PWM.n13048 ),
            .clk(N__56257),
            .ce(),
            .sr(N__48695));
    defparam \PWM.pwm_counter_664__i27_LC_14_31_3 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i27_LC_14_31_3 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i27_LC_14_31_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i27_LC_14_31_3  (
            .in0(_gnd_net_),
            .in1(N__48647),
            .in2(_gnd_net_),
            .in3(N__48717),
            .lcout(pwm_counter_27),
            .ltout(),
            .carryin(\PWM.n13048 ),
            .carryout(\PWM.n13049 ),
            .clk(N__56257),
            .ce(),
            .sr(N__48695));
    defparam \PWM.pwm_counter_664__i28_LC_14_31_4 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i28_LC_14_31_4 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i28_LC_14_31_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i28_LC_14_31_4  (
            .in0(_gnd_net_),
            .in1(N__48594),
            .in2(_gnd_net_),
            .in3(N__48714),
            .lcout(pwm_counter_28),
            .ltout(),
            .carryin(\PWM.n13049 ),
            .carryout(\PWM.n13050 ),
            .clk(N__56257),
            .ce(),
            .sr(N__48695));
    defparam \PWM.pwm_counter_664__i29_LC_14_31_5 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i29_LC_14_31_5 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i29_LC_14_31_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i29_LC_14_31_5  (
            .in0(_gnd_net_),
            .in1(N__48660),
            .in2(_gnd_net_),
            .in3(N__48711),
            .lcout(pwm_counter_29),
            .ltout(),
            .carryin(\PWM.n13050 ),
            .carryout(\PWM.n13051 ),
            .clk(N__56257),
            .ce(),
            .sr(N__48695));
    defparam \PWM.pwm_counter_664__i30_LC_14_31_6 .C_ON=1'b1;
    defparam \PWM.pwm_counter_664__i30_LC_14_31_6 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i30_LC_14_31_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i30_LC_14_31_6  (
            .in0(_gnd_net_),
            .in1(N__48621),
            .in2(_gnd_net_),
            .in3(N__48708),
            .lcout(pwm_counter_30),
            .ltout(),
            .carryin(\PWM.n13051 ),
            .carryout(\PWM.n13052 ),
            .clk(N__56257),
            .ce(),
            .sr(N__48695));
    defparam \PWM.pwm_counter_664__i31_LC_14_31_7 .C_ON=1'b0;
    defparam \PWM.pwm_counter_664__i31_LC_14_31_7 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_counter_664__i31_LC_14_31_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \PWM.pwm_counter_664__i31_LC_14_31_7  (
            .in0(_gnd_net_),
            .in1(N__50952),
            .in2(_gnd_net_),
            .in3(N__48705),
            .lcout(pwm_counter_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56257),
            .ce(),
            .sr(N__48695));
    defparam i5_4_lut_LC_14_32_5.C_ON=1'b0;
    defparam i5_4_lut_LC_14_32_5.SEQ_MODE=4'b0000;
    defparam i5_4_lut_LC_14_32_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i5_4_lut_LC_14_32_5 (
            .in0(N__48671),
            .in1(N__48659),
            .in2(N__48648),
            .in3(N__48632),
            .lcout(),
            .ltout(n12_adj_615_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_LC_14_32_6.C_ON=1'b0;
    defparam i6_4_lut_LC_14_32_6.SEQ_MODE=4'b0000;
    defparam i6_4_lut_LC_14_32_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_LC_14_32_6 (
            .in0(N__48620),
            .in1(N__48608),
            .in2(N__48597),
            .in3(N__48593),
            .lcout(n5180),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1047_3_lut_LC_15_17_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1047_3_lut_LC_15_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1047_3_lut_LC_15_17_1.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i1047_3_lut_LC_15_17_1 (
            .in0(_gnd_net_),
            .in1(N__51606),
            .in2(N__48885),
            .in3(N__51626),
            .lcout(n1631_adj_611),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i973_3_lut_LC_15_17_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i973_3_lut_LC_15_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i973_3_lut_LC_15_17_2.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i973_3_lut_LC_15_17_2 (
            .in0(_gnd_net_),
            .in1(N__51333),
            .in2(N__49007),
            .in3(N__51309),
            .lcout(n1525),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i1048_3_lut_LC_15_17_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i1048_3_lut_LC_15_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i1048_3_lut_LC_15_17_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i1048_3_lut_LC_15_17_4 (
            .in0(_gnd_net_),
            .in1(N__51662),
            .in2(N__51642),
            .in3(N__48866),
            .lcout(n1632_adj_612),
            .ltout(n1632_adj_612_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9943_3_lut_LC_15_17_5.C_ON=1'b0;
    defparam i9943_3_lut_LC_15_17_5.SEQ_MODE=4'b0000;
    defparam i9943_3_lut_LC_15_17_5.LUT_INIT=16'b1111000011000000;
    LogicCell40 i9943_3_lut_LC_15_17_5 (
            .in0(_gnd_net_),
            .in1(N__48787),
            .in2(N__48759),
            .in3(N__48742),
            .lcout(n11919),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i981_3_lut_LC_15_18_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i981_3_lut_LC_15_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i981_3_lut_LC_15_18_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 encoder0_position_31__I_0_i981_3_lut_LC_15_18_0 (
            .in0(N__50754),
            .in1(N__50718),
            .in2(_gnd_net_),
            .in3(N__48976),
            .lcout(n1533),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i972_3_lut_LC_15_18_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i972_3_lut_LC_15_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i972_3_lut_LC_15_18_1.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i972_3_lut_LC_15_18_1 (
            .in0(N__51855),
            .in1(_gnd_net_),
            .in2(N__48999),
            .in3(N__51843),
            .lcout(n1524),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i970_3_lut_LC_15_18_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i970_3_lut_LC_15_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i970_3_lut_LC_15_18_2.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i970_3_lut_LC_15_18_2 (
            .in0(_gnd_net_),
            .in1(N__51791),
            .in2(N__51765),
            .in3(N__48987),
            .lcout(n1522),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i978_3_lut_LC_15_18_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i978_3_lut_LC_15_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i978_3_lut_LC_15_18_3.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i978_3_lut_LC_15_18_3 (
            .in0(_gnd_net_),
            .in1(N__51476),
            .in2(N__49000),
            .in3(N__51450),
            .lcout(n1530),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i976_rep_49_3_lut_LC_15_18_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i976_rep_49_3_lut_LC_15_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i976_rep_49_3_lut_LC_15_18_4.LUT_INIT=16'b1111001111000000;
    LogicCell40 encoder0_position_31__I_0_i976_rep_49_3_lut_LC_15_18_4 (
            .in0(_gnd_net_),
            .in1(N__48972),
            .in2(N__52281),
            .in3(N__51408),
            .lcout(n1528),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i974_3_lut_LC_15_18_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i974_3_lut_LC_15_18_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i974_3_lut_LC_15_18_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i974_3_lut_LC_15_18_5 (
            .in0(N__51356),
            .in1(_gnd_net_),
            .in2(N__48998),
            .in3(N__51342),
            .lcout(n1526),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i980_3_lut_LC_15_18_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i980_3_lut_LC_15_18_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i980_3_lut_LC_15_18_6.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i980_3_lut_LC_15_18_6 (
            .in0(N__51519),
            .in1(_gnd_net_),
            .in2(N__51557),
            .in3(N__48980),
            .lcout(n1532),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i975_3_lut_LC_15_18_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i975_3_lut_LC_15_18_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i975_3_lut_LC_15_18_7.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i975_3_lut_LC_15_18_7 (
            .in0(_gnd_net_),
            .in1(N__51392),
            .in2(N__48997),
            .in3(N__51372),
            .lcout(n1527),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12842_1_lut_LC_15_19_0.C_ON=1'b0;
    defparam i12842_1_lut_LC_15_19_0.SEQ_MODE=4'b0000;
    defparam i12842_1_lut_LC_15_19_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12842_1_lut_LC_15_19_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48991),
            .lcout(n15572),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i905_3_lut_LC_15_19_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i905_3_lut_LC_15_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i905_3_lut_LC_15_19_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i905_3_lut_LC_15_19_1 (
            .in0(_gnd_net_),
            .in1(N__49050),
            .in2(N__49380),
            .in3(N__52343),
            .lcout(n1425),
            .ltout(n1425_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_110_LC_15_19_2.C_ON=1'b0;
    defparam i1_4_lut_adj_110_LC_15_19_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_110_LC_15_19_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_110_LC_15_19_2 (
            .in0(N__51325),
            .in1(N__51815),
            .in2(N__49041),
            .in3(N__49038),
            .lcout(),
            .ltout(n14490_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12845_4_lut_LC_15_19_3.C_ON=1'b0;
    defparam i12845_4_lut_LC_15_19_3.SEQ_MODE=4'b0000;
    defparam i12845_4_lut_LC_15_19_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12845_4_lut_LC_15_19_3 (
            .in0(N__51728),
            .in1(N__51781),
            .in2(N__49032),
            .in3(N__49101),
            .lcout(n1455),
            .ltout(n1455_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i979_3_lut_LC_15_19_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i979_3_lut_LC_15_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i979_3_lut_LC_15_19_4.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i979_3_lut_LC_15_19_4 (
            .in0(N__51489),
            .in1(_gnd_net_),
            .in2(N__49029),
            .in3(N__51503),
            .lcout(n1531),
            .ltout(n1531_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10020_4_lut_LC_15_19_5.C_ON=1'b0;
    defparam i10020_4_lut_LC_15_19_5.SEQ_MODE=4'b0000;
    defparam i10020_4_lut_LC_15_19_5.LUT_INIT=16'b1111111011110000;
    LogicCell40 i10020_4_lut_LC_15_19_5 (
            .in0(N__51658),
            .in1(N__51706),
            .in2(N__49026),
            .in3(N__51622),
            .lcout(n11997),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i977_3_lut_LC_15_19_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i977_3_lut_LC_15_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i977_3_lut_LC_15_19_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i977_3_lut_LC_15_19_6 (
            .in0(_gnd_net_),
            .in1(N__51420),
            .in2(N__51440),
            .in3(N__48992),
            .lcout(n1529),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i906_3_lut_LC_15_19_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i906_3_lut_LC_15_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i906_3_lut_LC_15_19_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i906_3_lut_LC_15_19_7 (
            .in0(_gnd_net_),
            .in1(N__49152),
            .in2(N__49260),
            .in3(N__52342),
            .lcout(n1426),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i903_3_lut_LC_15_20_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i903_3_lut_LC_15_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i903_3_lut_LC_15_20_0.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i903_3_lut_LC_15_20_0 (
            .in0(_gnd_net_),
            .in1(N__50000),
            .in2(N__52349),
            .in3(N__49146),
            .lcout(n1423),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9949_3_lut_LC_15_20_1.C_ON=1'b0;
    defparam i9949_3_lut_LC_15_20_1.SEQ_MODE=4'b0000;
    defparam i9949_3_lut_LC_15_20_1.LUT_INIT=16'b1111110000000000;
    LogicCell40 i9949_3_lut_LC_15_20_1 (
            .in0(_gnd_net_),
            .in1(N__49140),
            .in2(N__49079),
            .in3(N__49208),
            .lcout(),
            .ltout(n11925_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_106_LC_15_20_2.C_ON=1'b0;
    defparam i1_4_lut_adj_106_LC_15_20_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_106_LC_15_20_2.LUT_INIT=16'b1010100000000000;
    LogicCell40 i1_4_lut_adj_106_LC_15_20_2 (
            .in0(N__53113),
            .in1(N__49225),
            .in2(N__49113),
            .in3(N__49177),
            .lcout(n13720),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i910_3_lut_LC_15_20_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i910_3_lut_LC_15_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i910_3_lut_LC_15_20_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i910_3_lut_LC_15_20_3 (
            .in0(_gnd_net_),
            .in1(N__49110),
            .in2(N__49232),
            .in3(N__52338),
            .lcout(n1430),
            .ltout(n1430_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_108_LC_15_20_4.C_ON=1'b0;
    defparam i1_4_lut_adj_108_LC_15_20_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_108_LC_15_20_4.LUT_INIT=16'b1010000010000000;
    LogicCell40 i1_4_lut_adj_108_LC_15_20_4 (
            .in0(N__52276),
            .in1(N__51466),
            .in2(N__49104),
            .in3(N__49056),
            .lcout(n13739),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12826_4_lut_LC_15_20_5.C_ON=1'b0;
    defparam i12826_4_lut_LC_15_20_5.SEQ_MODE=4'b0000;
    defparam i12826_4_lut_LC_15_20_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12826_4_lut_LC_15_20_5 (
            .in0(N__49999),
            .in1(N__49266),
            .in2(N__52577),
            .in3(N__49095),
            .lcout(n1356),
            .ltout(n1356_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i912_3_lut_LC_15_20_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i912_3_lut_LC_15_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i912_3_lut_LC_15_20_6.LUT_INIT=16'b1111110000001100;
    LogicCell40 encoder0_position_31__I_0_i912_3_lut_LC_15_20_6 (
            .in0(_gnd_net_),
            .in1(N__49089),
            .in2(N__49083),
            .in3(N__49075),
            .lcout(n1432),
            .ltout(n1432_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9947_3_lut_LC_15_20_7.C_ON=1'b0;
    defparam i9947_3_lut_LC_15_20_7.SEQ_MODE=4'b0000;
    defparam i9947_3_lut_LC_15_20_7.LUT_INIT=16'b1111000011000000;
    LogicCell40 i9947_3_lut_LC_15_20_7 (
            .in0(_gnd_net_),
            .in1(N__50743),
            .in2(N__49059),
            .in3(N__51538),
            .lcout(n11923),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i840_3_lut_LC_15_21_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i840_3_lut_LC_15_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i840_3_lut_LC_15_21_0.LUT_INIT=16'b1111101000001010;
    LogicCell40 encoder0_position_31__I_0_i840_3_lut_LC_15_21_0 (
            .in0(N__52755),
            .in1(_gnd_net_),
            .in2(N__53180),
            .in3(N__52781),
            .lcout(n1328),
            .ltout(n1328_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_105_LC_15_21_1.C_ON=1'b0;
    defparam i1_4_lut_adj_105_LC_15_21_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_105_LC_15_21_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_4_lut_adj_105_LC_15_21_1 (
            .in0(N__49249),
            .in1(N__49369),
            .in2(N__49269),
            .in3(N__49657),
            .lcout(n14414),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i839_3_lut_LC_15_21_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i839_3_lut_LC_15_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i839_3_lut_LC_15_21_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i839_3_lut_LC_15_21_3 (
            .in0(_gnd_net_),
            .in1(N__52719),
            .in2(N__52746),
            .in3(N__53166),
            .lcout(n1327),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i843_3_lut_LC_15_21_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i843_3_lut_LC_15_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i843_3_lut_LC_15_21_4.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i843_3_lut_LC_15_21_4 (
            .in0(_gnd_net_),
            .in1(N__52178),
            .in2(N__53179),
            .in3(N__52158),
            .lcout(n1331),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i844_3_lut_LC_15_21_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i844_3_lut_LC_15_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i844_3_lut_LC_15_21_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i844_3_lut_LC_15_21_5 (
            .in0(_gnd_net_),
            .in1(N__52194),
            .in2(N__52214),
            .in3(N__53162),
            .lcout(n1332),
            .ltout(n1332_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i911_3_lut_LC_15_21_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i911_3_lut_LC_15_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i911_3_lut_LC_15_21_6.LUT_INIT=16'b1111000010101010;
    LogicCell40 encoder0_position_31__I_0_i911_3_lut_LC_15_21_6 (
            .in0(N__49197),
            .in1(_gnd_net_),
            .in2(N__49191),
            .in3(N__52331),
            .lcout(n1431),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i841_3_lut_LC_15_21_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i841_3_lut_LC_15_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i841_3_lut_LC_15_21_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i841_3_lut_LC_15_21_7 (
            .in0(_gnd_net_),
            .in1(N__52794),
            .in2(N__52821),
            .in3(N__53167),
            .lcout(n1329),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_101_LC_15_22_0.C_ON=1'b0;
    defparam i1_4_lut_adj_101_LC_15_22_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_101_LC_15_22_0.LUT_INIT=16'b1000100010000000;
    LogicCell40 i1_4_lut_adj_101_LC_15_22_0 (
            .in0(N__52813),
            .in1(N__52774),
            .in2(N__53221),
            .in3(N__49161),
            .lcout(),
            .ltout(n13723_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12810_4_lut_LC_15_22_1.C_ON=1'b0;
    defparam i12810_4_lut_LC_15_22_1.SEQ_MODE=4'b0000;
    defparam i12810_4_lut_LC_15_22_1.LUT_INIT=16'b0000000000000001;
    LogicCell40 i12810_4_lut_LC_15_22_1 (
            .in0(N__52652),
            .in1(N__49344),
            .in2(N__49155),
            .in3(N__52601),
            .lcout(n1257),
            .ltout(n1257_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i837_3_lut_LC_15_22_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i837_3_lut_LC_15_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i837_3_lut_LC_15_22_2.LUT_INIT=16'b1010111110100000;
    LogicCell40 encoder0_position_31__I_0_i837_3_lut_LC_15_22_2 (
            .in0(N__52679),
            .in1(_gnd_net_),
            .in2(N__49671),
            .in3(N__52665),
            .lcout(n1325),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12807_1_lut_LC_15_22_3.C_ON=1'b0;
    defparam i12807_1_lut_LC_15_22_3.SEQ_MODE=4'b0000;
    defparam i12807_1_lut_LC_15_22_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 i12807_1_lut_LC_15_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53171),
            .lcout(n15537),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_mux_3_i22_3_lut_LC_15_22_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_mux_3_i22_3_lut_LC_15_22_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_mux_3_i22_3_lut_LC_15_22_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 encoder0_position_31__I_0_mux_3_i22_3_lut_LC_15_22_4 (
            .in0(N__49641),
            .in1(N__49622),
            .in2(_gnd_net_),
            .in3(N__52416),
            .lcout(n298),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i838_3_lut_LC_15_22_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i838_3_lut_LC_15_22_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i838_3_lut_LC_15_22_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i838_3_lut_LC_15_22_5 (
            .in0(_gnd_net_),
            .in1(N__52692),
            .in2(N__52710),
            .in3(N__53172),
            .lcout(n1326),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i771_3_lut_LC_15_22_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i771_3_lut_LC_15_22_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i771_3_lut_LC_15_22_6.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i771_3_lut_LC_15_22_6 (
            .in0(_gnd_net_),
            .in1(N__49806),
            .in2(N__49943),
            .in3(N__49353),
            .lcout(n1227),
            .ltout(n1227_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_100_LC_15_22_7.C_ON=1'b0;
    defparam i1_3_lut_adj_100_LC_15_22_7.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_100_LC_15_22_7.LUT_INIT=16'b1111111111111100;
    LogicCell40 i1_3_lut_adj_100_LC_15_22_7 (
            .in0(_gnd_net_),
            .in1(N__52732),
            .in2(N__49347),
            .in3(N__52678),
            .lcout(n14476),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i775_3_lut_LC_15_23_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i775_3_lut_LC_15_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i775_3_lut_LC_15_23_0.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i775_3_lut_LC_15_23_0 (
            .in0(_gnd_net_),
            .in1(N__49338),
            .in2(N__49332),
            .in3(N__49928),
            .lcout(n1231),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i703_3_lut_LC_15_23_1.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i703_3_lut_LC_15_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i703_3_lut_LC_15_23_1.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i703_3_lut_LC_15_23_1 (
            .in0(_gnd_net_),
            .in1(N__52859),
            .in2(N__49876),
            .in3(N__52833),
            .lcout(n1127),
            .ltout(n1127_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i770_3_lut_LC_15_23_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i770_3_lut_LC_15_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i770_3_lut_LC_15_23_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i770_3_lut_LC_15_23_2 (
            .in0(_gnd_net_),
            .in1(N__49296),
            .in2(N__49290),
            .in3(N__49929),
            .lcout(n1226),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i769_3_lut_LC_15_23_3.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i769_3_lut_LC_15_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i769_3_lut_LC_15_23_3.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i769_3_lut_LC_15_23_3 (
            .in0(_gnd_net_),
            .in1(N__50034),
            .in2(N__49942),
            .in3(N__50010),
            .lcout(n1225),
            .ltout(n1225_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i836_3_lut_LC_15_23_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i836_3_lut_LC_15_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i836_3_lut_LC_15_23_4.LUT_INIT=16'b1110010011100100;
    LogicCell40 encoder0_position_31__I_0_i836_3_lut_LC_15_23_4 (
            .in0(N__53175),
            .in1(N__52641),
            .in2(N__50004),
            .in3(_gnd_net_),
            .lcout(n1324),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i772_3_lut_LC_15_23_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i772_3_lut_LC_15_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i772_3_lut_LC_15_23_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i772_3_lut_LC_15_23_6 (
            .in0(_gnd_net_),
            .in1(N__49983),
            .in2(N__49962),
            .in3(N__49930),
            .lcout(n1228),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i704_3_lut_LC_15_23_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i704_3_lut_LC_15_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i704_3_lut_LC_15_23_7.LUT_INIT=16'b1100111111000000;
    LogicCell40 encoder0_position_31__I_0_i704_3_lut_LC_15_23_7 (
            .in0(_gnd_net_),
            .in1(N__52895),
            .in2(N__49875),
            .in3(N__52869),
            .lcout(n1128),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_305_1_LC_15_25_0.C_ON=1'b1;
    defparam add_305_1_LC_15_25_0.SEQ_MODE=4'b0000;
    defparam add_305_1_LC_15_25_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_305_1_LC_15_25_0 (
            .in0(_gnd_net_),
            .in1(N__51118),
            .in2(N__51164),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_25_0_),
            .carryout(n12449),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i0_LC_15_25_1.C_ON=1'b1;
    defparam encoder0_position_target_i0_i0_LC_15_25_1.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i0_LC_15_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i0_LC_15_25_1 (
            .in0(_gnd_net_),
            .in1(N__49762),
            .in2(N__49782),
            .in3(N__49743),
            .lcout(encoder0_position_target_0),
            .ltout(),
            .carryin(n12449),
            .carryout(n12450),
            .clk(N__56234),
            .ce(N__55881),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i1_LC_15_25_2.C_ON=1'b1;
    defparam encoder0_position_target_i0_i1_LC_15_25_2.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i1_LC_15_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i1_LC_15_25_2 (
            .in0(_gnd_net_),
            .in1(N__51119),
            .in2(N__49735),
            .in3(N__49707),
            .lcout(encoder0_position_target_1),
            .ltout(),
            .carryin(n12450),
            .carryout(n12451),
            .clk(N__56234),
            .ce(N__55881),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i2_LC_15_25_3.C_ON=1'b1;
    defparam encoder0_position_target_i0_i2_LC_15_25_3.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i2_LC_15_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i2_LC_15_25_3 (
            .in0(_gnd_net_),
            .in1(N__51125),
            .in2(N__49703),
            .in3(N__49674),
            .lcout(encoder0_position_target_2),
            .ltout(),
            .carryin(n12451),
            .carryout(n12452),
            .clk(N__56234),
            .ce(N__55881),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i3_LC_15_25_4.C_ON=1'b1;
    defparam encoder0_position_target_i0_i3_LC_15_25_4.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i3_LC_15_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i3_LC_15_25_4 (
            .in0(_gnd_net_),
            .in1(N__51120),
            .in2(N__50351),
            .in3(N__50322),
            .lcout(encoder0_position_target_3),
            .ltout(),
            .carryin(n12452),
            .carryout(n12453),
            .clk(N__56234),
            .ce(N__55881),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i4_LC_15_25_5.C_ON=1'b1;
    defparam encoder0_position_target_i0_i4_LC_15_25_5.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i4_LC_15_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i4_LC_15_25_5 (
            .in0(_gnd_net_),
            .in1(N__51126),
            .in2(N__50317),
            .in3(N__50277),
            .lcout(encoder0_position_target_4),
            .ltout(),
            .carryin(n12453),
            .carryout(n12454),
            .clk(N__56234),
            .ce(N__55881),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i5_LC_15_25_6.C_ON=1'b1;
    defparam encoder0_position_target_i0_i5_LC_15_25_6.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i5_LC_15_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i5_LC_15_25_6 (
            .in0(_gnd_net_),
            .in1(N__51121),
            .in2(N__50270),
            .in3(N__50241),
            .lcout(encoder0_position_target_5),
            .ltout(),
            .carryin(n12454),
            .carryout(n12455),
            .clk(N__56234),
            .ce(N__55881),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i6_LC_15_25_7.C_ON=1'b1;
    defparam encoder0_position_target_i0_i6_LC_15_25_7.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i6_LC_15_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i6_LC_15_25_7 (
            .in0(_gnd_net_),
            .in1(N__51127),
            .in2(N__50237),
            .in3(N__50205),
            .lcout(encoder0_position_target_6),
            .ltout(),
            .carryin(n12455),
            .carryout(n12456),
            .clk(N__56234),
            .ce(N__55881),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i7_LC_15_26_0.C_ON=1'b1;
    defparam encoder0_position_target_i0_i7_LC_15_26_0.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i7_LC_15_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i7_LC_15_26_0 (
            .in0(_gnd_net_),
            .in1(N__50181),
            .in2(N__51165),
            .in3(N__50160),
            .lcout(encoder0_position_target_7),
            .ltout(),
            .carryin(bfn_15_26_0_),
            .carryout(n12457),
            .clk(N__56239),
            .ce(N__55916),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i8_LC_15_26_1.C_ON=1'b1;
    defparam encoder0_position_target_i0_i8_LC_15_26_1.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i8_LC_15_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i8_LC_15_26_1 (
            .in0(_gnd_net_),
            .in1(N__51131),
            .in2(N__50152),
            .in3(N__50121),
            .lcout(encoder0_position_target_8),
            .ltout(),
            .carryin(n12457),
            .carryout(n12458),
            .clk(N__56239),
            .ce(N__55916),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i9_LC_15_26_2.C_ON=1'b1;
    defparam encoder0_position_target_i0_i9_LC_15_26_2.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i9_LC_15_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i9_LC_15_26_2 (
            .in0(_gnd_net_),
            .in1(N__50106),
            .in2(N__51166),
            .in3(N__50079),
            .lcout(encoder0_position_target_9),
            .ltout(),
            .carryin(n12458),
            .carryout(n12459),
            .clk(N__56239),
            .ce(N__55916),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i10_LC_15_26_3.C_ON=1'b1;
    defparam encoder0_position_target_i0_i10_LC_15_26_3.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i10_LC_15_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i10_LC_15_26_3 (
            .in0(_gnd_net_),
            .in1(N__51135),
            .in2(N__50070),
            .in3(N__50037),
            .lcout(encoder0_position_target_10),
            .ltout(),
            .carryin(n12459),
            .carryout(n12460),
            .clk(N__56239),
            .ce(N__55916),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i11_LC_15_26_4.C_ON=1'b1;
    defparam encoder0_position_target_i0_i11_LC_15_26_4.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i11_LC_15_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i11_LC_15_26_4 (
            .in0(_gnd_net_),
            .in1(N__50704),
            .in2(N__51167),
            .in3(N__50679),
            .lcout(encoder0_position_target_11),
            .ltout(),
            .carryin(n12460),
            .carryout(n12461),
            .clk(N__56239),
            .ce(N__55916),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i12_LC_15_26_5.C_ON=1'b1;
    defparam encoder0_position_target_i0_i12_LC_15_26_5.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i12_LC_15_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i12_LC_15_26_5 (
            .in0(_gnd_net_),
            .in1(N__51139),
            .in2(N__50675),
            .in3(N__50640),
            .lcout(encoder0_position_target_12),
            .ltout(),
            .carryin(n12461),
            .carryout(n12462),
            .clk(N__56239),
            .ce(N__55916),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i13_LC_15_26_6.C_ON=1'b1;
    defparam encoder0_position_target_i0_i13_LC_15_26_6.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i13_LC_15_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i13_LC_15_26_6 (
            .in0(_gnd_net_),
            .in1(N__50629),
            .in2(N__51168),
            .in3(N__50601),
            .lcout(encoder0_position_target_13),
            .ltout(),
            .carryin(n12462),
            .carryout(n12463),
            .clk(N__56239),
            .ce(N__55916),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i14_LC_15_26_7.C_ON=1'b1;
    defparam encoder0_position_target_i0_i14_LC_15_26_7.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i14_LC_15_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i14_LC_15_26_7 (
            .in0(_gnd_net_),
            .in1(N__51143),
            .in2(N__50597),
            .in3(N__50568),
            .lcout(encoder0_position_target_14),
            .ltout(),
            .carryin(n12463),
            .carryout(n12464),
            .clk(N__56239),
            .ce(N__55916),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i15_LC_15_27_0.C_ON=1'b1;
    defparam encoder0_position_target_i0_i15_LC_15_27_0.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i15_LC_15_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i15_LC_15_27_0 (
            .in0(_gnd_net_),
            .in1(N__51169),
            .in2(N__50558),
            .in3(N__50520),
            .lcout(encoder0_position_target_15),
            .ltout(),
            .carryin(bfn_15_27_0_),
            .carryout(n12465),
            .clk(N__56247),
            .ce(N__55898),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i16_LC_15_27_1.C_ON=1'b1;
    defparam encoder0_position_target_i0_i16_LC_15_27_1.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i16_LC_15_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i16_LC_15_27_1 (
            .in0(_gnd_net_),
            .in1(N__50509),
            .in2(N__51186),
            .in3(N__50484),
            .lcout(encoder0_position_target_16),
            .ltout(),
            .carryin(n12465),
            .carryout(n12466),
            .clk(N__56247),
            .ce(N__55898),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i17_LC_15_27_2.C_ON=1'b1;
    defparam encoder0_position_target_i0_i17_LC_15_27_2.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i17_LC_15_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i17_LC_15_27_2 (
            .in0(_gnd_net_),
            .in1(N__51173),
            .in2(N__50477),
            .in3(N__50439),
            .lcout(encoder0_position_target_17),
            .ltout(),
            .carryin(n12466),
            .carryout(n12467),
            .clk(N__56247),
            .ce(N__55898),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i18_LC_15_27_3.C_ON=1'b1;
    defparam encoder0_position_target_i0_i18_LC_15_27_3.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i18_LC_15_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i18_LC_15_27_3 (
            .in0(_gnd_net_),
            .in1(N__50429),
            .in2(N__51187),
            .in3(N__50400),
            .lcout(encoder0_position_target_18),
            .ltout(),
            .carryin(n12467),
            .carryout(n12468),
            .clk(N__56247),
            .ce(N__55898),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i19_LC_15_27_4.C_ON=1'b1;
    defparam encoder0_position_target_i0_i19_LC_15_27_4.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i19_LC_15_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i19_LC_15_27_4 (
            .in0(_gnd_net_),
            .in1(N__51177),
            .in2(N__50391),
            .in3(N__50355),
            .lcout(encoder0_position_target_19),
            .ltout(),
            .carryin(n12468),
            .carryout(n12469),
            .clk(N__56247),
            .ce(N__55898),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i20_LC_15_27_5.C_ON=1'b1;
    defparam encoder0_position_target_i0_i20_LC_15_27_5.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i20_LC_15_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i20_LC_15_27_5 (
            .in0(_gnd_net_),
            .in1(N__51296),
            .in2(N__51188),
            .in3(N__51273),
            .lcout(encoder0_position_target_20),
            .ltout(),
            .carryin(n12469),
            .carryout(n12470),
            .clk(N__56247),
            .ce(N__55898),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i21_LC_15_27_6.C_ON=1'b1;
    defparam encoder0_position_target_i0_i21_LC_15_27_6.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i21_LC_15_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i21_LC_15_27_6 (
            .in0(_gnd_net_),
            .in1(N__51181),
            .in2(N__51264),
            .in3(N__51231),
            .lcout(encoder0_position_target_21),
            .ltout(),
            .carryin(n12470),
            .carryout(n12471),
            .clk(N__56247),
            .ce(N__55898),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i22_LC_15_27_7.C_ON=1'b1;
    defparam encoder0_position_target_i0_i22_LC_15_27_7.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i22_LC_15_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_target_i0_i22_LC_15_27_7 (
            .in0(_gnd_net_),
            .in1(N__51220),
            .in2(N__51189),
            .in3(N__51192),
            .lcout(encoder0_position_target_22),
            .ltout(),
            .carryin(n12471),
            .carryout(n12472),
            .clk(N__56247),
            .ce(N__55898),
            .sr(_gnd_net_));
    defparam encoder0_position_target_i0_i23_LC_15_28_0.C_ON=1'b0;
    defparam encoder0_position_target_i0_i23_LC_15_28_0.SEQ_MODE=4'b1000;
    defparam encoder0_position_target_i0_i23_LC_15_28_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 encoder0_position_target_i0_i23_LC_15_28_0 (
            .in0(N__51185),
            .in1(N__51037),
            .in2(_gnd_net_),
            .in3(N__51057),
            .lcout(encoder0_position_target_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56253),
            .ce(N__55911),
            .sr(_gnd_net_));
    defparam \PWM.pwm_out_12_LC_15_30_6 .C_ON=1'b0;
    defparam \PWM.pwm_out_12_LC_15_30_6 .SEQ_MODE=4'b1000;
    defparam \PWM.pwm_out_12_LC_15_30_6 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \PWM.pwm_out_12_LC_15_30_6  (
            .in0(N__50997),
            .in1(N__50982),
            .in2(_gnd_net_),
            .in3(N__50964),
            .lcout(pwm_out),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56258),
            .ce(),
            .sr(N__50919));
    defparam i1_2_lut_adj_44_LC_15_31_1.C_ON=1'b0;
    defparam i1_2_lut_adj_44_LC_15_31_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_44_LC_15_31_1.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1_2_lut_adj_44_LC_15_31_1 (
            .in0(_gnd_net_),
            .in1(N__50950),
            .in2(_gnd_net_),
            .in3(N__50933),
            .lcout(n5182),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dir_160_LC_15_31_7.C_ON=1'b0;
    defparam dir_160_LC_15_31_7.SEQ_MODE=4'b1000;
    defparam dir_160_LC_15_31_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 dir_160_LC_15_31_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50909),
            .lcout(dir),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56259),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_2_lut_LC_16_17_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_2_lut_LC_16_17_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_2_lut_LC_16_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_2_lut_LC_16_17_0 (
            .in0(_gnd_net_),
            .in1(N__50750),
            .in2(_gnd_net_),
            .in3(N__50712),
            .lcout(n1501),
            .ltout(),
            .carryin(bfn_16_17_0_),
            .carryout(n12552),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_3_lut_LC_16_17_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_3_lut_LC_16_17_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_3_lut_LC_16_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_3_lut_LC_16_17_1 (
            .in0(_gnd_net_),
            .in1(N__55128),
            .in2(N__51558),
            .in3(N__51513),
            .lcout(n1500),
            .ltout(),
            .carryin(n12552),
            .carryout(n12553),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_4_lut_LC_16_17_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_4_lut_LC_16_17_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_4_lut_LC_16_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_4_lut_LC_16_17_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51510),
            .in3(N__51480),
            .lcout(n1499),
            .ltout(),
            .carryin(n12553),
            .carryout(n12554),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_5_lut_LC_16_17_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_5_lut_LC_16_17_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_5_lut_LC_16_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_5_lut_LC_16_17_3 (
            .in0(_gnd_net_),
            .in1(N__55129),
            .in2(N__51477),
            .in3(N__51444),
            .lcout(n1498),
            .ltout(),
            .carryin(n12554),
            .carryout(n12555),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_6_lut_LC_16_17_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_6_lut_LC_16_17_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_6_lut_LC_16_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_6_lut_LC_16_17_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51441),
            .in3(N__51411),
            .lcout(n1497),
            .ltout(),
            .carryin(n12555),
            .carryout(n12556),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_7_lut_LC_16_17_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_7_lut_LC_16_17_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_7_lut_LC_16_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_7_lut_LC_16_17_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__52280),
            .in3(N__51402),
            .lcout(n1496),
            .ltout(),
            .carryin(n12556),
            .carryout(n12557),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_8_lut_LC_16_17_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_8_lut_LC_16_17_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_8_lut_LC_16_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_8_lut_LC_16_17_6 (
            .in0(_gnd_net_),
            .in1(N__55131),
            .in2(N__51399),
            .in3(N__51366),
            .lcout(n1495),
            .ltout(),
            .carryin(n12557),
            .carryout(n12558),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_9_lut_LC_16_17_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_9_lut_LC_16_17_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_9_lut_LC_16_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_9_lut_LC_16_17_7 (
            .in0(_gnd_net_),
            .in1(N__55130),
            .in2(N__51363),
            .in3(N__51336),
            .lcout(n1494),
            .ltout(),
            .carryin(n12558),
            .carryout(n12559),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_10_lut_LC_16_18_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_10_lut_LC_16_18_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_10_lut_LC_16_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_10_lut_LC_16_18_0 (
            .in0(_gnd_net_),
            .in1(N__55121),
            .in2(N__51332),
            .in3(N__51303),
            .lcout(n1493),
            .ltout(),
            .carryin(bfn_16_18_0_),
            .carryout(n12560),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_11_lut_LC_16_18_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_11_lut_LC_16_18_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_11_lut_LC_16_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_11_lut_LC_16_18_1 (
            .in0(_gnd_net_),
            .in1(N__51854),
            .in2(N__55288),
            .in3(N__51837),
            .lcout(n1492),
            .ltout(),
            .carryin(n12560),
            .carryout(n12561),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_12_lut_LC_16_18_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_12_lut_LC_16_18_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_12_lut_LC_16_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_12_lut_LC_16_18_2 (
            .in0(_gnd_net_),
            .in1(N__55125),
            .in2(N__51833),
            .in3(N__51795),
            .lcout(n1491),
            .ltout(),
            .carryin(n12561),
            .carryout(n12562),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_13_lut_LC_16_18_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_967_13_lut_LC_16_18_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_13_lut_LC_16_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_967_13_lut_LC_16_18_3 (
            .in0(_gnd_net_),
            .in1(N__55126),
            .in2(N__51792),
            .in3(N__51756),
            .lcout(n1490),
            .ltout(),
            .carryin(n12562),
            .carryout(n12563),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_967_14_lut_LC_16_18_4.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_967_14_lut_LC_16_18_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_967_14_lut_LC_16_18_4.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_967_14_lut_LC_16_18_4 (
            .in0(N__55127),
            .in1(N__51746),
            .in2(N__51735),
            .in3(N__51714),
            .lcout(n1521),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_2_lut_LC_16_19_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_2_lut_LC_16_19_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_2_lut_LC_16_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_2_lut_LC_16_19_0 (
            .in0(_gnd_net_),
            .in1(N__51711),
            .in2(_gnd_net_),
            .in3(N__51666),
            .lcout(n1601),
            .ltout(),
            .carryin(bfn_16_19_0_),
            .carryout(n12564),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_3_lut_LC_16_19_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_3_lut_LC_16_19_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_3_lut_LC_16_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_3_lut_LC_16_19_1 (
            .in0(_gnd_net_),
            .in1(N__55117),
            .in2(N__51663),
            .in3(N__51630),
            .lcout(n1600),
            .ltout(),
            .carryin(n12564),
            .carryout(n12565),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_4_lut_LC_16_19_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_4_lut_LC_16_19_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_4_lut_LC_16_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_4_lut_LC_16_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__51627),
            .in3(N__51597),
            .lcout(n1599),
            .ltout(),
            .carryin(n12565),
            .carryout(n12566),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_5_lut_LC_16_19_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_5_lut_LC_16_19_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_5_lut_LC_16_19_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_5_lut_LC_16_19_3 (
            .in0(_gnd_net_),
            .in1(N__55118),
            .in2(N__51590),
            .in3(N__51561),
            .lcout(n1598),
            .ltout(),
            .carryin(n12566),
            .carryout(n12567),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_6_lut_LC_16_19_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_6_lut_LC_16_19_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_6_lut_LC_16_19_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_6_lut_LC_16_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__52148),
            .in3(N__52113),
            .lcout(n1597),
            .ltout(),
            .carryin(n12567),
            .carryout(n12568),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_7_lut_LC_16_19_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_7_lut_LC_16_19_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_7_lut_LC_16_19_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_7_lut_LC_16_19_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__52110),
            .in3(N__52080),
            .lcout(n1596),
            .ltout(),
            .carryin(n12568),
            .carryout(n12569),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_8_lut_LC_16_19_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_8_lut_LC_16_19_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_8_lut_LC_16_19_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_8_lut_LC_16_19_6 (
            .in0(_gnd_net_),
            .in1(N__55120),
            .in2(N__52076),
            .in3(N__52038),
            .lcout(n1595),
            .ltout(),
            .carryin(n12569),
            .carryout(n12570),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_9_lut_LC_16_19_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_9_lut_LC_16_19_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_9_lut_LC_16_19_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_9_lut_LC_16_19_7 (
            .in0(_gnd_net_),
            .in1(N__55119),
            .in2(N__52034),
            .in3(N__52002),
            .lcout(n1594),
            .ltout(),
            .carryin(n12570),
            .carryout(n12571),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_10_lut_LC_16_20_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_10_lut_LC_16_20_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_10_lut_LC_16_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_10_lut_LC_16_20_0 (
            .in0(_gnd_net_),
            .in1(N__51992),
            .in2(N__55278),
            .in3(N__51957),
            .lcout(n1593),
            .ltout(),
            .carryin(bfn_16_20_0_),
            .carryout(n12572),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_11_lut_LC_16_20_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_11_lut_LC_16_20_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_11_lut_LC_16_20_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_11_lut_LC_16_20_1 (
            .in0(_gnd_net_),
            .in1(N__55091),
            .in2(N__51954),
            .in3(N__51915),
            .lcout(n1592),
            .ltout(),
            .carryin(n12572),
            .carryout(n12573),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_12_lut_LC_16_20_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_12_lut_LC_16_20_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_12_lut_LC_16_20_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_12_lut_LC_16_20_2 (
            .in0(_gnd_net_),
            .in1(N__55096),
            .in2(N__51912),
            .in3(N__51879),
            .lcout(n1591),
            .ltout(),
            .carryin(n12573),
            .carryout(n12574),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_13_lut_LC_16_20_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_13_lut_LC_16_20_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_13_lut_LC_16_20_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_13_lut_LC_16_20_3 (
            .in0(_gnd_net_),
            .in1(N__55092),
            .in2(N__51876),
            .in3(N__52539),
            .lcout(n1590),
            .ltout(),
            .carryin(n12574),
            .carryout(n12575),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_14_lut_LC_16_20_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_1034_14_lut_LC_16_20_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_14_lut_LC_16_20_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_1034_14_lut_LC_16_20_4 (
            .in0(_gnd_net_),
            .in1(N__52532),
            .in2(N__55279),
            .in3(N__52500),
            .lcout(n1589),
            .ltout(),
            .carryin(n12575),
            .carryout(n12576),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_1034_15_lut_LC_16_20_5.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_1034_15_lut_LC_16_20_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_1034_15_lut_LC_16_20_5.LUT_INIT=16'b1001000001100000;
    LogicCell40 encoder0_position_31__I_0_add_1034_15_lut_LC_16_20_5 (
            .in0(N__55097),
            .in1(N__52497),
            .in2(N__52475),
            .in3(N__52446),
            .lcout(n1620_adj_600),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut_LC_16_20_6.C_ON=1'b0;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut_LC_16_20_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut_LC_16_20_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut_LC_16_20_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52409),
            .lcout(n12_adj_630),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i909_3_lut_LC_16_20_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i909_3_lut_LC_16_20_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i909_3_lut_LC_16_20_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 encoder0_position_31__I_0_i909_3_lut_LC_16_20_7 (
            .in0(_gnd_net_),
            .in1(N__53114),
            .in2(N__52371),
            .in3(N__52337),
            .lcout(n1429),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_2_lut_LC_16_21_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_2_lut_LC_16_21_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_2_lut_LC_16_21_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_2_lut_LC_16_21_0 (
            .in0(_gnd_net_),
            .in1(N__52247),
            .in2(_gnd_net_),
            .in3(N__52221),
            .lcout(n1301),
            .ltout(),
            .carryin(bfn_16_21_0_),
            .carryout(n12531),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_3_lut_LC_16_21_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_3_lut_LC_16_21_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_3_lut_LC_16_21_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_3_lut_LC_16_21_1 (
            .in0(_gnd_net_),
            .in1(N__54650),
            .in2(N__52218),
            .in3(N__52188),
            .lcout(n1300),
            .ltout(),
            .carryin(n12531),
            .carryout(n12532),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_4_lut_LC_16_21_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_4_lut_LC_16_21_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_4_lut_LC_16_21_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_4_lut_LC_16_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__52185),
            .in3(N__52152),
            .lcout(n1299),
            .ltout(),
            .carryin(n12532),
            .carryout(n12533),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_5_lut_LC_16_21_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_5_lut_LC_16_21_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_5_lut_LC_16_21_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_5_lut_LC_16_21_3 (
            .in0(_gnd_net_),
            .in1(N__54651),
            .in2(N__53223),
            .in3(N__52824),
            .lcout(n1298),
            .ltout(),
            .carryin(n12533),
            .carryout(n12534),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_6_lut_LC_16_21_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_6_lut_LC_16_21_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_6_lut_LC_16_21_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_6_lut_LC_16_21_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__52820),
            .in3(N__52788),
            .lcout(n1297),
            .ltout(),
            .carryin(n12534),
            .carryout(n12535),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_7_lut_LC_16_21_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_7_lut_LC_16_21_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_7_lut_LC_16_21_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_7_lut_LC_16_21_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__52785),
            .in3(N__52749),
            .lcout(n1296),
            .ltout(),
            .carryin(n12535),
            .carryout(n12536),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_8_lut_LC_16_21_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_8_lut_LC_16_21_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_8_lut_LC_16_21_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_8_lut_LC_16_21_6 (
            .in0(_gnd_net_),
            .in1(N__54653),
            .in2(N__52745),
            .in3(N__52713),
            .lcout(n1295),
            .ltout(),
            .carryin(n12536),
            .carryout(n12537),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_9_lut_LC_16_21_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_9_lut_LC_16_21_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_9_lut_LC_16_21_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_9_lut_LC_16_21_7 (
            .in0(_gnd_net_),
            .in1(N__54652),
            .in2(N__52709),
            .in3(N__52686),
            .lcout(n1294),
            .ltout(),
            .carryin(n12537),
            .carryout(n12538),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_10_lut_LC_16_22_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_10_lut_LC_16_22_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_10_lut_LC_16_22_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_10_lut_LC_16_22_0 (
            .in0(_gnd_net_),
            .in1(N__54647),
            .in2(N__52683),
            .in3(N__52659),
            .lcout(n1293),
            .ltout(),
            .carryin(bfn_16_22_0_),
            .carryout(n12539),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_11_lut_LC_16_22_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_833_11_lut_LC_16_22_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_11_lut_LC_16_22_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_833_11_lut_LC_16_22_1 (
            .in0(_gnd_net_),
            .in1(N__54648),
            .in2(N__52656),
            .in3(N__52635),
            .lcout(n1292),
            .ltout(),
            .carryin(n12539),
            .carryout(n12540),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_833_12_lut_LC_16_22_2.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_833_12_lut_LC_16_22_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_833_12_lut_LC_16_22_2.LUT_INIT=16'b1000010001001000;
    LogicCell40 encoder0_position_31__I_0_add_833_12_lut_LC_16_22_2 (
            .in0(N__54649),
            .in1(N__52619),
            .in2(N__52608),
            .in3(N__52584),
            .lcout(n1323),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_i842_3_lut_LC_16_22_7.C_ON=1'b0;
    defparam encoder0_position_31__I_0_i842_3_lut_LC_16_22_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_i842_3_lut_LC_16_22_7.LUT_INIT=16'b1111000011001100;
    LogicCell40 encoder0_position_31__I_0_i842_3_lut_LC_16_22_7 (
            .in0(_gnd_net_),
            .in1(N__53229),
            .in2(N__53222),
            .in3(N__53173),
            .lcout(n1330),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_2_lut_LC_16_23_0.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_2_lut_LC_16_23_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_2_lut_LC_16_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_2_lut_LC_16_23_0 (
            .in0(_gnd_net_),
            .in1(N__53091),
            .in2(_gnd_net_),
            .in3(N__53058),
            .lcout(n1101),
            .ltout(),
            .carryin(bfn_16_23_0_),
            .carryout(n12514),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_3_lut_LC_16_23_1.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_3_lut_LC_16_23_1.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_3_lut_LC_16_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_3_lut_LC_16_23_1 (
            .in0(_gnd_net_),
            .in1(N__54643),
            .in2(N__53055),
            .in3(N__53025),
            .lcout(n1100),
            .ltout(),
            .carryin(n12514),
            .carryout(n12515),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_4_lut_LC_16_23_2.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_4_lut_LC_16_23_2.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_4_lut_LC_16_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_4_lut_LC_16_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__53022),
            .in3(N__52983),
            .lcout(n1099),
            .ltout(),
            .carryin(n12515),
            .carryout(n12516),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_5_lut_LC_16_23_3.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_5_lut_LC_16_23_3.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_5_lut_LC_16_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_5_lut_LC_16_23_3 (
            .in0(_gnd_net_),
            .in1(N__54644),
            .in2(N__52980),
            .in3(N__52941),
            .lcout(n1098),
            .ltout(),
            .carryin(n12516),
            .carryout(n12517),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_6_lut_LC_16_23_4.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_6_lut_LC_16_23_4.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_6_lut_LC_16_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_6_lut_LC_16_23_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__52938),
            .in3(N__52899),
            .lcout(n1097),
            .ltout(),
            .carryin(n12517),
            .carryout(n12518),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_7_lut_LC_16_23_5.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_7_lut_LC_16_23_5.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_7_lut_LC_16_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_7_lut_LC_16_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__52896),
            .in3(N__52863),
            .lcout(n1096),
            .ltout(),
            .carryin(n12518),
            .carryout(n12519),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_8_lut_LC_16_23_6.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_8_lut_LC_16_23_6.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_8_lut_LC_16_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_8_lut_LC_16_23_6 (
            .in0(_gnd_net_),
            .in1(N__54646),
            .in2(N__52860),
            .in3(N__52827),
            .lcout(n1095),
            .ltout(),
            .carryin(n12519),
            .carryout(n12520),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_9_lut_LC_16_23_7.C_ON=1'b1;
    defparam encoder0_position_31__I_0_add_699_9_lut_LC_16_23_7.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_9_lut_LC_16_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_9_lut_LC_16_23_7 (
            .in0(_gnd_net_),
            .in1(N__54645),
            .in2(N__55599),
            .in3(N__55566),
            .lcout(n1094),
            .ltout(),
            .carryin(n12520),
            .carryout(n12521),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam encoder0_position_31__I_0_add_699_10_lut_LC_16_24_0.C_ON=1'b0;
    defparam encoder0_position_31__I_0_add_699_10_lut_LC_16_24_0.SEQ_MODE=4'b0000;
    defparam encoder0_position_31__I_0_add_699_10_lut_LC_16_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 encoder0_position_31__I_0_add_699_10_lut_LC_16_24_0 (
            .in0(_gnd_net_),
            .in1(N__53791),
            .in2(N__53385),
            .in3(N__53358),
            .lcout(n1093),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam sweep_counter_660_661__i1_LC_16_25_0.C_ON=1'b1;
    defparam sweep_counter_660_661__i1_LC_16_25_0.SEQ_MODE=4'b1000;
    defparam sweep_counter_660_661__i1_LC_16_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_660_661__i1_LC_16_25_0 (
            .in0(_gnd_net_),
            .in1(N__53345),
            .in2(_gnd_net_),
            .in3(N__53331),
            .lcout(sweep_counter_0),
            .ltout(),
            .carryin(bfn_16_25_0_),
            .carryout(n13053),
            .clk(N__56240),
            .ce(),
            .sr(N__55897));
    defparam sweep_counter_660_661__i2_LC_16_25_1.C_ON=1'b1;
    defparam sweep_counter_660_661__i2_LC_16_25_1.SEQ_MODE=4'b1000;
    defparam sweep_counter_660_661__i2_LC_16_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_660_661__i2_LC_16_25_1 (
            .in0(_gnd_net_),
            .in1(N__53327),
            .in2(_gnd_net_),
            .in3(N__53313),
            .lcout(sweep_counter_1),
            .ltout(),
            .carryin(n13053),
            .carryout(n13054),
            .clk(N__56240),
            .ce(),
            .sr(N__55897));
    defparam sweep_counter_660_661__i3_LC_16_25_2.C_ON=1'b1;
    defparam sweep_counter_660_661__i3_LC_16_25_2.SEQ_MODE=4'b1000;
    defparam sweep_counter_660_661__i3_LC_16_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_660_661__i3_LC_16_25_2 (
            .in0(_gnd_net_),
            .in1(N__53309),
            .in2(_gnd_net_),
            .in3(N__53292),
            .lcout(sweep_counter_2),
            .ltout(),
            .carryin(n13054),
            .carryout(n13055),
            .clk(N__56240),
            .ce(),
            .sr(N__55897));
    defparam sweep_counter_660_661__i4_LC_16_25_3.C_ON=1'b1;
    defparam sweep_counter_660_661__i4_LC_16_25_3.SEQ_MODE=4'b1000;
    defparam sweep_counter_660_661__i4_LC_16_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_660_661__i4_LC_16_25_3 (
            .in0(_gnd_net_),
            .in1(N__53285),
            .in2(_gnd_net_),
            .in3(N__53271),
            .lcout(sweep_counter_3),
            .ltout(),
            .carryin(n13055),
            .carryout(n13056),
            .clk(N__56240),
            .ce(),
            .sr(N__55897));
    defparam sweep_counter_660_661__i5_LC_16_25_4.C_ON=1'b1;
    defparam sweep_counter_660_661__i5_LC_16_25_4.SEQ_MODE=4'b1000;
    defparam sweep_counter_660_661__i5_LC_16_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_660_661__i5_LC_16_25_4 (
            .in0(_gnd_net_),
            .in1(N__53264),
            .in2(_gnd_net_),
            .in3(N__53250),
            .lcout(sweep_counter_4),
            .ltout(),
            .carryin(n13056),
            .carryout(n13057),
            .clk(N__56240),
            .ce(),
            .sr(N__55897));
    defparam sweep_counter_660_661__i6_LC_16_25_5.C_ON=1'b1;
    defparam sweep_counter_660_661__i6_LC_16_25_5.SEQ_MODE=4'b1000;
    defparam sweep_counter_660_661__i6_LC_16_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_660_661__i6_LC_16_25_5 (
            .in0(_gnd_net_),
            .in1(N__53246),
            .in2(_gnd_net_),
            .in3(N__53232),
            .lcout(sweep_counter_5),
            .ltout(),
            .carryin(n13057),
            .carryout(n13058),
            .clk(N__56240),
            .ce(),
            .sr(N__55897));
    defparam sweep_counter_660_661__i7_LC_16_25_6.C_ON=1'b1;
    defparam sweep_counter_660_661__i7_LC_16_25_6.SEQ_MODE=4'b1000;
    defparam sweep_counter_660_661__i7_LC_16_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_660_661__i7_LC_16_25_6 (
            .in0(_gnd_net_),
            .in1(N__55715),
            .in2(_gnd_net_),
            .in3(N__55701),
            .lcout(sweep_counter_6),
            .ltout(),
            .carryin(n13058),
            .carryout(n13059),
            .clk(N__56240),
            .ce(),
            .sr(N__55897));
    defparam sweep_counter_660_661__i8_LC_16_25_7.C_ON=1'b1;
    defparam sweep_counter_660_661__i8_LC_16_25_7.SEQ_MODE=4'b1000;
    defparam sweep_counter_660_661__i8_LC_16_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_660_661__i8_LC_16_25_7 (
            .in0(_gnd_net_),
            .in1(N__55694),
            .in2(_gnd_net_),
            .in3(N__55680),
            .lcout(sweep_counter_7),
            .ltout(),
            .carryin(n13059),
            .carryout(n13060),
            .clk(N__56240),
            .ce(),
            .sr(N__55897));
    defparam sweep_counter_660_661__i9_LC_16_26_0.C_ON=1'b1;
    defparam sweep_counter_660_661__i9_LC_16_26_0.SEQ_MODE=4'b1000;
    defparam sweep_counter_660_661__i9_LC_16_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_660_661__i9_LC_16_26_0 (
            .in0(_gnd_net_),
            .in1(N__55835),
            .in2(_gnd_net_),
            .in3(N__55677),
            .lcout(sweep_counter_8),
            .ltout(),
            .carryin(bfn_16_26_0_),
            .carryout(n13061),
            .clk(N__56248),
            .ce(),
            .sr(N__55912));
    defparam sweep_counter_660_661__i10_LC_16_26_1.C_ON=1'b1;
    defparam sweep_counter_660_661__i10_LC_16_26_1.SEQ_MODE=4'b1000;
    defparam sweep_counter_660_661__i10_LC_16_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_660_661__i10_LC_16_26_1 (
            .in0(_gnd_net_),
            .in1(N__55667),
            .in2(_gnd_net_),
            .in3(N__55653),
            .lcout(sweep_counter_9),
            .ltout(),
            .carryin(n13061),
            .carryout(n13062),
            .clk(N__56248),
            .ce(),
            .sr(N__55912));
    defparam sweep_counter_660_661__i11_LC_16_26_2.C_ON=1'b1;
    defparam sweep_counter_660_661__i11_LC_16_26_2.SEQ_MODE=4'b1000;
    defparam sweep_counter_660_661__i11_LC_16_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_660_661__i11_LC_16_26_2 (
            .in0(_gnd_net_),
            .in1(N__55646),
            .in2(_gnd_net_),
            .in3(N__55632),
            .lcout(sweep_counter_10),
            .ltout(),
            .carryin(n13062),
            .carryout(n13063),
            .clk(N__56248),
            .ce(),
            .sr(N__55912));
    defparam sweep_counter_660_661__i12_LC_16_26_3.C_ON=1'b1;
    defparam sweep_counter_660_661__i12_LC_16_26_3.SEQ_MODE=4'b1000;
    defparam sweep_counter_660_661__i12_LC_16_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_660_661__i12_LC_16_26_3 (
            .in0(_gnd_net_),
            .in1(N__55625),
            .in2(_gnd_net_),
            .in3(N__55611),
            .lcout(sweep_counter_11),
            .ltout(),
            .carryin(n13063),
            .carryout(n13064),
            .clk(N__56248),
            .ce(),
            .sr(N__55912));
    defparam sweep_counter_660_661__i13_LC_16_26_4.C_ON=1'b1;
    defparam sweep_counter_660_661__i13_LC_16_26_4.SEQ_MODE=4'b1000;
    defparam sweep_counter_660_661__i13_LC_16_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_660_661__i13_LC_16_26_4 (
            .in0(_gnd_net_),
            .in1(N__55775),
            .in2(_gnd_net_),
            .in3(N__55608),
            .lcout(sweep_counter_12),
            .ltout(),
            .carryin(n13064),
            .carryout(n13065),
            .clk(N__56248),
            .ce(),
            .sr(N__55912));
    defparam sweep_counter_660_661__i14_LC_16_26_5.C_ON=1'b1;
    defparam sweep_counter_660_661__i14_LC_16_26_5.SEQ_MODE=4'b1000;
    defparam sweep_counter_660_661__i14_LC_16_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_660_661__i14_LC_16_26_5 (
            .in0(_gnd_net_),
            .in1(N__55805),
            .in2(_gnd_net_),
            .in3(N__55605),
            .lcout(sweep_counter_13),
            .ltout(),
            .carryin(n13065),
            .carryout(n13066),
            .clk(N__56248),
            .ce(),
            .sr(N__55912));
    defparam sweep_counter_660_661__i15_LC_16_26_6.C_ON=1'b1;
    defparam sweep_counter_660_661__i15_LC_16_26_6.SEQ_MODE=4'b1000;
    defparam sweep_counter_660_661__i15_LC_16_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_660_661__i15_LC_16_26_6 (
            .in0(_gnd_net_),
            .in1(N__55820),
            .in2(_gnd_net_),
            .in3(N__55602),
            .lcout(sweep_counter_14),
            .ltout(),
            .carryin(n13066),
            .carryout(n13067),
            .clk(N__56248),
            .ce(),
            .sr(N__55912));
    defparam sweep_counter_660_661__i16_LC_16_26_7.C_ON=1'b1;
    defparam sweep_counter_660_661__i16_LC_16_26_7.SEQ_MODE=4'b1000;
    defparam sweep_counter_660_661__i16_LC_16_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_660_661__i16_LC_16_26_7 (
            .in0(_gnd_net_),
            .in1(N__55955),
            .in2(_gnd_net_),
            .in3(N__55941),
            .lcout(sweep_counter_15),
            .ltout(),
            .carryin(n13067),
            .carryout(n13068),
            .clk(N__56248),
            .ce(),
            .sr(N__55912));
    defparam sweep_counter_660_661__i17_LC_16_27_0.C_ON=1'b1;
    defparam sweep_counter_660_661__i17_LC_16_27_0.SEQ_MODE=4'b1000;
    defparam sweep_counter_660_661__i17_LC_16_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_660_661__i17_LC_16_27_0 (
            .in0(_gnd_net_),
            .in1(N__55937),
            .in2(_gnd_net_),
            .in3(N__55923),
            .lcout(sweep_counter_16),
            .ltout(),
            .carryin(bfn_16_27_0_),
            .carryout(n13069),
            .clk(N__56254),
            .ce(),
            .sr(N__55917));
    defparam sweep_counter_660_661__i18_LC_16_27_1.C_ON=1'b0;
    defparam sweep_counter_660_661__i18_LC_16_27_1.SEQ_MODE=4'b1000;
    defparam sweep_counter_660_661__i18_LC_16_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 sweep_counter_660_661__i18_LC_16_27_1 (
            .in0(_gnd_net_),
            .in1(N__55791),
            .in2(_gnd_net_),
            .in3(N__55920),
            .lcout(sweep_counter_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56254),
            .ce(),
            .sr(N__55917));
    defparam i1_2_lut_adj_74_LC_16_28_5.C_ON=1'b0;
    defparam i1_2_lut_adj_74_LC_16_28_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_74_LC_16_28_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 i1_2_lut_adj_74_LC_16_28_5 (
            .in0(_gnd_net_),
            .in1(N__55836),
            .in2(_gnd_net_),
            .in3(N__55821),
            .lcout(),
            .ltout(n6_adj_712_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_adj_75_LC_16_28_6.C_ON=1'b0;
    defparam i4_4_lut_adj_75_LC_16_28_6.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_75_LC_16_28_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 i4_4_lut_adj_75_LC_16_28_6 (
            .in0(N__55806),
            .in1(N__55790),
            .in2(N__55779),
            .in3(N__55776),
            .lcout(n13968),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GHC_174_LC_16_31_6.C_ON=1'b0;
    defparam GHC_174_LC_16_31_6.SEQ_MODE=4'b1000;
    defparam GHC_174_LC_16_31_6.LUT_INIT=16'b0101010110000010;
    LogicCell40 GHC_174_LC_16_31_6 (
            .in0(N__56353),
            .in1(N__56516),
            .in2(N__56439),
            .in3(N__56328),
            .lcout(GHC),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56260),
            .ce(N__56056),
            .sr(N__56029));
    defparam GHB_172_LC_17_31_4.C_ON=1'b0;
    defparam GHB_172_LC_17_31_4.SEQ_MODE=4'b1000;
    defparam GHB_172_LC_17_31_4.LUT_INIT=16'b1001100000000011;
    LogicCell40 GHB_172_LC_17_31_4 (
            .in0(N__56515),
            .in1(N__56323),
            .in2(N__56440),
            .in3(N__56354),
            .lcout(GHB),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56261),
            .ce(N__56063),
            .sr(N__56030));
    defparam i9546_2_lut_LC_17_32_5.C_ON=1'b0;
    defparam i9546_2_lut_LC_17_32_5.SEQ_MODE=4'b0000;
    defparam i9546_2_lut_LC_17_32_5.LUT_INIT=16'b1010101000000000;
    LogicCell40 i9546_2_lut_LC_17_32_5 (
            .in0(N__55994),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55734),
            .lcout(INHC_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9545_2_lut_LC_17_32_6.C_ON=1'b0;
    defparam i9545_2_lut_LC_17_32_6.SEQ_MODE=4'b0000;
    defparam i9545_2_lut_LC_17_32_6.LUT_INIT=16'b1100110000000000;
    LogicCell40 i9545_2_lut_LC_17_32_6 (
            .in0(_gnd_net_),
            .in1(N__55993),
            .in2(_gnd_net_),
            .in3(N__56571),
            .lcout(INHB_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GHA_170_LC_18_31_2.C_ON=1'b0;
    defparam GHA_170_LC_18_31_2.SEQ_MODE=4'b1000;
    defparam GHA_170_LC_18_31_2.LUT_INIT=16'b0001010010011000;
    LogicCell40 GHA_170_LC_18_31_2 (
            .in0(N__56324),
            .in1(N__56355),
            .in2(N__56441),
            .in3(N__56513),
            .lcout(GHA),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56262),
            .ce(N__56064),
            .sr(N__56034));
    defparam GLA_171_LC_18_31_5.C_ON=1'b0;
    defparam GLA_171_LC_18_31_5.SEQ_MODE=4'b1000;
    defparam GLA_171_LC_18_31_5.LUT_INIT=16'b0000010111000010;
    LogicCell40 GLA_171_LC_18_31_5 (
            .in0(N__56512),
            .in1(N__56431),
            .in2(N__56363),
            .in3(N__56326),
            .lcout(INLA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56262),
            .ce(N__56064),
            .sr(N__56034));
    defparam GLB_173_LC_18_31_6.C_ON=1'b0;
    defparam GLB_173_LC_18_31_6.SEQ_MODE=4'b1000;
    defparam GLB_173_LC_18_31_6.LUT_INIT=16'b0010011000010100;
    LogicCell40 GLB_173_LC_18_31_6 (
            .in0(N__56325),
            .in1(N__56359),
            .in2(N__56442),
            .in3(N__56514),
            .lcout(INLB_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56262),
            .ce(N__56064),
            .sr(N__56034));
    defparam GLC_175_LC_18_31_7.C_ON=1'b0;
    defparam GLC_175_LC_18_31_7.SEQ_MODE=4'b1000;
    defparam GLC_175_LC_18_31_7.LUT_INIT=16'b1111000000001001;
    LogicCell40 GLC_175_LC_18_31_7 (
            .in0(N__56511),
            .in1(N__56432),
            .in2(N__56364),
            .in3(N__56327),
            .lcout(INLC_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56262),
            .ce(N__56064),
            .sr(N__56034));
    defparam i9544_2_lut_LC_18_32_0.C_ON=1'b0;
    defparam i9544_2_lut_LC_18_32_0.SEQ_MODE=4'b0000;
    defparam i9544_2_lut_LC_18_32_0.LUT_INIT=16'b1010101000000000;
    LogicCell40 i9544_2_lut_LC_18_32_0 (
            .in0(N__56001),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55995),
            .lcout(INHA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
