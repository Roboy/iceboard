// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Mon Feb  3 22:48:23 2020
//
// Verilog Description of module TinyFPGA_B
//

module TinyFPGA_B (CLK, LED, USBPU, ENCODER0_A, ENCODER0_B, ENCODER1_A, 
            ENCODER1_B, HALL1, HALL2, HALL3, FAULT_N, NEOPXL, DE, 
            TX, RX, CS_CLK, CS, CS_MISO, SCL, SDA, INLC, INHC, 
            INLB, INHB, INLA, INHA) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(2[8:18])
    input CLK;   // verilog/TinyFPGA_B.v(3[9:12])
    output LED;   // verilog/TinyFPGA_B.v(4[10:13])
    output USBPU;   // verilog/TinyFPGA_B.v(5[10:15])
    input ENCODER0_A;   // verilog/TinyFPGA_B.v(6[9:19])
    input ENCODER0_B;   // verilog/TinyFPGA_B.v(7[9:19])
    input ENCODER1_A;   // verilog/TinyFPGA_B.v(8[9:19])
    input ENCODER1_B;   // verilog/TinyFPGA_B.v(9[9:19])
    input HALL1 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(10[9:14])
    input HALL2 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(11[9:14])
    input HALL3 /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(12[9:14])
    input FAULT_N;   // verilog/TinyFPGA_B.v(13[9:16])
    output NEOPXL;   // verilog/TinyFPGA_B.v(14[10:16])
    output DE;   // verilog/TinyFPGA_B.v(15[10:12])
    output TX /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(16[10:12])
    input RX;   // verilog/TinyFPGA_B.v(17[9:11])
    output CS_CLK;   // verilog/TinyFPGA_B.v(18[10:16])
    output CS;   // verilog/TinyFPGA_B.v(19[10:12])
    input CS_MISO;   // verilog/TinyFPGA_B.v(20[9:16])
    inout SCL /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(21[9:12])
    inout SDA /* synthesis black_box_pad_pin=1 */ ;   // verilog/TinyFPGA_B.v(22[9:12])
    output INLC;   // verilog/TinyFPGA_B.v(23[10:14])
    output INHC;   // verilog/TinyFPGA_B.v(24[10:14])
    output INLB;   // verilog/TinyFPGA_B.v(25[10:14])
    output INHB;   // verilog/TinyFPGA_B.v(26[10:14])
    output INLA;   // verilog/TinyFPGA_B.v(27[10:14])
    output INHA;   // verilog/TinyFPGA_B.v(28[10:14])
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    wire GND_net, VCC_net, LED_c, ENCODER0_A_N, ENCODER0_B_N, ENCODER1_A_N, 
        ENCODER1_B_N, NEOPXL_c, DE_c, RX_c, INHC_c, INLB_c, INHB_c, 
        INLA_c, INHA_c;
    wire [7:0]ID;   // verilog/TinyFPGA_B.v(39[11:13])
    wire [23:0]neopxl_color;   // verilog/TinyFPGA_B.v(41[13:25])
    
    wire hall1, hall2, hall3;
    wire [22:0]pwm_setpoint;   // verilog/TinyFPGA_B.v(87[13:25])
    wire [23:0]duty;   // verilog/TinyFPGA_B.v(88[21:25])
    
    wire tx_o, tx_enable;
    wire [23:0]encoder0_position_scaled;   // verilog/TinyFPGA_B.v(125[21:45])
    wire [23:0]encoder1_position_scaled;   // verilog/TinyFPGA_B.v(127[21:45])
    wire [23:0]displacement;   // verilog/TinyFPGA_B.v(128[21:33])
    wire [23:0]setpoint;   // verilog/TinyFPGA_B.v(129[22:30])
    wire [23:0]Kp;   // verilog/TinyFPGA_B.v(130[22:24])
    wire [23:0]Ki;   // verilog/TinyFPGA_B.v(131[22:24])
    
    wire n39778;
    wire [7:0]control_mode;   // verilog/TinyFPGA_B.v(133[14:26])
    wire [23:0]PWMLimit;   // verilog/TinyFPGA_B.v(134[22:30])
    wire [23:0]IntegralLimit;   // verilog/TinyFPGA_B.v(135[22:35])
    
    wire n40209, n39777, n39776;
    wire [23:0]motor_state;   // verilog/TinyFPGA_B.v(165[22:33])
    
    wire n516;
    wire [7:0]data;   // verilog/TinyFPGA_B.v(228[14:18])
    
    wire data_ready, sda_out, sda_enable, scl, scl_enable;
    wire [31:0]delay_counter;   // verilog/TinyFPGA_B.v(252[11:24])
    
    wire read;
    wire [2:0]\ID_READOUT_FSM.state ;   // verilog/TinyFPGA_B.v(260[15:20])
    wire [22:0]pwm_setpoint_22__N_11;
    
    wire RX_N_10;
    wire [31:0]encoder0_position;   // verilog/TinyFPGA_B.v(124[11:28])
    
    wire n1152;
    wire [31:0]motor_state_23__N_106;
    wire [32:0]encoder0_position_scaled_23__N_34;
    
    wire encoder1_position_scaled_23__N_231;
    wire [31:0]encoder1_position_scaled_23__N_58;
    wire [23:0]displacement_23__N_82;
    
    wire n659, n660, n661, n662, n663, n664, n665, n666, n667, 
        n668, n669, n670, n671, n672, n673, n674, n675, n676, 
        n677, n678, n679, n680, n681, n682, n683, n684, n685, 
        n686, n687, n688, n689, n690, read_N_321, n7, n777, 
        n43797, n39775, n39774, n39773, n40208, n40207, n40206, 
        n40205, n39772, n1193;
    wire [31:0]encoder1_position;   // verilog/TinyFPGA_B.v(126[11:28])
    wire [31:0]timer;   // verilog/neopixel.v(9[12:17])
    wire [3:0]state;   // verilog/neopixel.v(16[20:25])
    
    wire start, \neo_pixel_transmitter.done ;
    wire [31:0]\neo_pixel_transmitter.t0 ;   // verilog/neopixel.v(28[14:16])
    
    wire n39771, n39770, n28315, n28314, n28313, n28312, n28311, 
        n28310, n28309, n28308, n28307, n39769, n40204;
    wire [3:0]state_3__N_428;
    
    wire n40203, n39768, n40202, n40201, n39767, n39766, n39765, 
        n40200, n40199, n40198, n40197, n4227, n39764, n40196, 
        n40195, n26645, n40194, n39763, n39762, n2, n40193, n15, 
        n40192, n46363, n5728, n28306, n28305, n40191, n40190, 
        n39761, n39760, n28304, n28303;
    wire [31:0]pwm_counter;   // verilog/pwm.v(11[9:20])
    
    wire n15_adj_4885, n28302, n40189, n28301, n3, n4, n5, n6, 
        n7_adj_4886, n8, n9, n10, n11, n12, n13, n14, n15_adj_4887, 
        n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, 
        n33765, rx_data_ready;
    wire [7:0]rx_data;   // verilog/coms.v(91[13:20])
    wire [7:0]\data_in[3] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[2] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[1] ;   // verilog/coms.v(95[12:19])
    wire [7:0]\data_in[0] ;   // verilog/coms.v(95[12:19])
    
    wire n40188;
    wire [7:0]\data_in_frame[13] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[12] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[11] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[10] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[9] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[8] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[6] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[5] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[4] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[3] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[2] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[1] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_out_frame[25] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[24] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[23] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[20] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[19] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[18] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[17] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[16] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[15] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[14] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[13] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[12] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[11] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[10] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[9] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[8] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[7] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[6] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[5] ;   // verilog/coms.v(97[12:26])
    wire [7:0]\data_out_frame[4] ;   // verilog/coms.v(97[12:26])
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(102[12:33])
    wire [31:0]\FRAME_MATCHER.state ;   // verilog/coms.v(112[11:16])
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(115[11:12])
    
    wire n12_adj_4888, n40187, n40186, n39759, n39758, n39757, n50224, 
        n25_adj_4889, n17_adj_4890, n45174, n44839, n45531, n43285, 
        n50222, n39756, n50509, n28300, n39755, n40185, n39754, 
        n40184, n39753, n39752, n771, n40183, n33298, n33302, 
        n46360, n33308, n5_adj_4891, n6_adj_4892, n7_adj_4893, n8_adj_4894, 
        n9_adj_4895, n10_adj_4896, n11_adj_4897, n12_adj_4898, n13_adj_4899, 
        n14_adj_4900, n15_adj_4901, n16_adj_4902, n17_adj_4903, n18_adj_4904, 
        n19_adj_4905, n20_adj_4906, n21_adj_4907, n22_adj_4908, n23_adj_4909, 
        n24_adj_4910, n25_adj_4911, n40182, n40181, n40180, n39751, 
        n39750, n39749, n40179, n40178, n40177, n39748, n40176, 
        n39747, n39013, n40175, n39746, n39012, n45105, n40174, 
        n40173, n40172, n40171, n39745, n39744, n39743, n34801, 
        n40170, n39742, n39380, n39741, n39740, n39379, n40169, 
        n39739, n40168, n39738, n39378, n38997, n39377, n39011, 
        n40167, n40166, n40165, n39737, n40164, n40163, n40162, 
        n39376, n39736, n39735, n51302, n38996, n39010, n39724, 
        n39539, n39538, n39723, n39537, n40152, n39722, n39536, 
        n39535, n34735, n40151, n39534, n39721, n39720, n40150, 
        n45026, n39719, n39009, n38995, n40149, n40148, n39718, 
        n40147, n39717, n40146, n39920, n39919, n39716, n39715, 
        n34707, n39714, n40145, n39918, n40144, n40143, n39713, 
        n40142, n39917, n39916, n39915, n39712, n39711, n45088, 
        n39710, n45047, n40141, n40140, n39914, n39709, n39708, 
        n40139, n39707, n40138, n39913, n39912, n39706, n39705, 
        n40137, n39008, n40136, n39911, n40135, n40134, n39704, 
        n51056, n39703, n40133, n39910, n39702, n39701, n39909, 
        n40132, n39908, n40131, n39700, n39699, n39907, n39906, 
        n39905, n39007, n39698, n39697, n40130, n39696, n39904, 
        n40129, tx_transmit_N_3413, n39903, n40128, n34693, n28299, 
        n40127, n50593, n39902, n39695, n39694, n3303, n39693, 
        n40126, n50933, n40, n51237, n39901, n40125, n40124, n39692, 
        n39691, n26480, n40123, n39690, n40122, n4452, n40121, 
        n38994, n39689, n39688, n40120, n40119, n5_adj_4912, n15_adj_4913, 
        n44805, n40118, n40117, n39043, n39042, n39687, n40116, 
        n40115, n40114, n39686, n29985, n76, n73, n74, n61, 
        n40113, n34457, n34677, n39685, n40112, n39041, n39040, 
        n40111, n40110, n39684, n39683, n39682, n51904, n44120, 
        n45377, n43085, n40109, n39681, n4_adj_4914, n4_adj_4915, 
        \FRAME_MATCHER.i_31__N_2524 , \FRAME_MATCHER.i_31__N_2526 , n40534, 
        n40108, n40107, n40533, n40532, n40531, n40530, n40106, 
        n40529, n40528, n40527, n40105, n40526, n40525, n40325, 
        n40104, n40524, n40324, n40523, n40522, n40323, n34475, 
        n34471, n34461, n34459, n34641, n34334, n34393, n34671, 
        n28771, n28770, n28769, n28768, n28767, n28766, n28765, 
        n40521, n40103, n40322, n40321, n40320, n40520, n40102, 
        n40519, n40101, n40319, n40100, n28759, n28758, n28757, 
        n28756, n28755, n28754, n28753, n28752, n28751, n28750, 
        n28749, n28748, n28747, n28746, n28745, n28744, n28743, 
        n28742, n28741, n28740, n28739, n28738, n28737, n28736, 
        n28735, n28734, n28733, n28732, n4_adj_4916, n28731, n28730, 
        n40518, n40517, n39680, n39679, n40318, n33, n32, n31, 
        n30, n29, n28, n27, n26, n25_adj_4917, n24_adj_4918, n23_adj_4919, 
        n22_adj_4920, n21_adj_4921, n20_adj_4922, n19_adj_4923, n18_adj_4924, 
        n17_adj_4925, n16_adj_4926, n15_adj_4927, n14_adj_4928, n13_adj_4929, 
        n12_adj_4930, n11_adj_4931, n10_adj_4932, n9_adj_4933, n8_adj_4934, 
        n28729, n28728, n28727, n40317, n40099, n40516, n10_adj_4935, 
        n40515, n28726, n28725, n28724, n28723, n40514, n28722, 
        n28721, n28720, n40098, n40316, n40097, n3_adj_4936, n4_adj_4937, 
        n28719, n28718, n28717, n28716, n28715, n28714, n28713, 
        n5722, n28712, n28298, n28297, n28296, n28295, n28294, 
        n28293, n28292, n28291, n28290, n28289, n28288, n28287, 
        n28286, n28285, n28284, n28283, n28282, n28281, n28280, 
        n28279, n28278, n28277, n28276, n28275, n28274, n28273, 
        n28272, n28271, n28270, n28269, n28268, n28267, n28266, 
        n28711, n28710, n28709, n28708, n28707, n28706, n28705, 
        n28704, n28703, n28702, n28701, n28700, n28699, n28698, 
        n28697, n40315, n28696, n40314, n40313, n28695, n28694, 
        n28693, n28692, n28691, n28690, n28689, n28688, n28687, 
        n28686, n28685, n28684, n28683, n28682, n28681, n28680, 
        n28679, n28678, n28677, n28676, n28675, n28674, n28673, 
        n28672, n28671, n28670, n28669, n28668, n28667, n28666, 
        n28665, n28664, n28663, n28662, n28661, n28660, n28659, 
        n28658, n28657, n28656, n28655, n28654, n28653, n40312, 
        n40096, n40095, n40513, n40512, n40311, n40094, n39678, 
        n40310, n40093, n40511, n40309, n40308, n40092, n40091, 
        n39039, n39038, n40090, n39677, n39676, n39675, n39674, 
        n40089, n40307, n39673, n40510, n40306, n40088, n39672, 
        n40305, n40087, n40086, n28652, n28651, n28650, n28649, 
        n28648, n28647, n28646, n28645, n40085, n28644, n28643, 
        n28642, n28641, n28640, n28639, n28638, n28637, n40509, 
        n40508, n39671, n40304, n28636, n28635, n4_adj_4938, n28634, 
        n28633, n28632, n39670, n28631, n28630, n28629, n28628;
    wire [1:0]a_new;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire b_prev, n28627, n28626, n28625, n28624, n28623, n28622, 
        n28621, n28620, n28619, n28618, n28617, n34637, n28616, 
        n28615, n28614, n1476, n28613, n28612, n28611, n28610, 
        n28609, n28608, n39669, n28607, n28606, direction_N_3807, 
        n28605, n28604, n28603, n28602, n28601, n28600, n28599, 
        n28598, n28597, n28596, n28595, n28594, n28593, n28592, 
        n28591, n28590, n28589, n28588, n28587, n28586, n39323, 
        n28585, n40507, n28584, n28583, n39668, n40084, n40303, 
        n28265, n39322, n28264, n39667, n40302, n28582, n39666, 
        n40506, n28263, n28262, n28261, n28260, n28259, n28258, 
        n28257, n28256, n28255, n28581, n40505, n28580, n39321, 
        n40083, n40504, n40082, n28579;
    wire [1:0]a_new_adj_5076;   // vhdl/quadrature_decoder.vhd(40[9:14])
    
    wire b_prev_adj_4940, n28578, n28577, n28576, n28575, n28574, 
        n28573, n28572, n28571, n39665, n2482, n40081, n1419, 
        n39320, n28570, n28569, n28568, n40301, n28567, direction_N_3807_adj_4941, 
        n44092, n28566, n28565, n4_adj_4942, n28564, n28563, n28561, 
        n28560, n28559, n28558, n28557, n28556, n28555, n40080, 
        n40300, n40299, n40298, n5855, n28554, n28553, n40079, 
        n40078, n40297, n40296, n40295, n40294, n40293, n40292, 
        n6014, n40291, n28552, n40290, n28551, n40077, n39319, 
        n40289, n39318, n40076, n40075, n40288, n40074, n28550, 
        n28549, n28548, n28547, n28250, n28246, n28241, n40073, 
        n43685, n28234, n28546, n40072, n40287, rw;
    wire [7:0]state_adj_5100;   // verilog/eeprom.v(23[11:16])
    
    wire n15_adj_4945, n14_adj_4946, n40071, n40286, n40070, n40285, 
        n40284, n28545, n28544, n28543, n28542, n28541, n28540, 
        n39317, n5_adj_4947, n28539, n28538, n28537, n28536, n28535, 
        n28534, n28533, n28532, n39316, n28531, n28530, n7_adj_4948, 
        n6_adj_4949, n5_adj_4950, n4_adj_4951, n3_adj_4952, n2_adj_4953, 
        r_Rx_Data;
    wire [2:0]r_Bit_Index;   // verilog/uart_rx.v(33[17:28])
    wire [2:0]r_SM_Main;   // verilog/uart_rx.v(36[17:26])
    
    wire n28529, n28528, n28527;
    wire [2:0]r_SM_Main_2__N_3442;
    
    wire n28526, n28525, n28524, n28523, n28522, n28521, n28520, 
        n28519, n28518, n28517, n28516, n28515, n28514, n28513, 
        n28512, n40069, n40283, n40068, n28511, n28510, n28509, 
        n28508, n40282, n28507, n28506, n28505, n28504, n28503, 
        n28502, n28501, n40067, n39315, n28500, n28499, n28498, 
        n28497, n28496, n28495, n28494, n28493, n40281;
    wire [7:0]state_adj_5116;   // verilog/i2c_controller.v(33[12:17])
    
    wire n10_adj_4955;
    wire [7:0]saved_addr;   // verilog/i2c_controller.v(34[12:22])
    
    wire n40066, enable_slow_N_4090, n40280, n39314, n40065, n40279, 
        n40278, n40064, n39313, n39312, n39311;
    wire [7:0]state_7__N_3987;
    
    wire n39654, n40063, n40062, n39653, n28230, n5538, n40277, 
        n40061, n40060, n45439;
    wire [7:0]state_7__N_4003;
    
    wire n34629, n26489, n40276, n42985, n39652, n40275, n34657, 
        n39651, n39650, n40274, n28225, n28224, n28223, n28222, 
        n40273, n39649, n40272, n39648, n45178, n621, n622, n623, 
        n625, n652, n40059, n39647, n731, n6539, n6538, n6537, 
        n6536, n6535, n6534, n828, n829, n830, n831, n832, n833, 
        n834, n51203, n27916, n861, n896, n897, n898, n899, 
        n900, n901, n927, n928, n929, n930, n931, n932, n933, 
        n934, n935, n936, n937, n938, n939, n940, n941, n942, 
        n943, n944, n945, n946, n947, n948, n949, n950, n951, 
        n952, n953, n954, n955, n956, n957, n960, n995, n996, 
        n997, n998, n999, n1000, n1001, n1026, n1027, n1028, 
        n1029, n1030, n1031, n1032, n1033, n1059, n1093, n1094, 
        n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1125, 
        n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, 
        n1158, n1193_adj_4956, n1194, n1195, n1196, n1197, n1198, 
        n1199, n1200, n1201, n1224, n1225, n1226, n1227, n1228, 
        n1229, n1230, n1231, n1232, n1233, n1257, n1292, n1293, 
        n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, 
        n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, 
        n1331, n1332, n1333, n1356, n1391, n1392, n1393, n1394, 
        n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1422, 
        n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, 
        n1431, n1432, n1433, n1455, n1490, n1491, n1492, n1493, 
        n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, 
        n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, 
        n1529, n1530, n1531, n1532, n1533, n1554, n12_adj_4957, 
        n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
        n1597, n1598, n1599, n1600, n1601, n43693, n1620, n1621, 
        n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, 
        n1630, n1631, n1632, n1633, n28044, n1653, n40058, n1688, 
        n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
        n1697, n1698, n1699, n1700, n1701, n40271, n47577, n40057, 
        n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
        n1727, n1728, n1729, n1730, n1731, n1732, n1733, n47571, 
        n40270, n1752, n47565, n40056, n1787, n1788, n1789, n1790, 
        n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, 
        n1799, n1800, n1801, n50798, n44859, n1818, n1819, n1820, 
        n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, 
        n1829, n1830, n1831, n1832, n1833, n8_adj_4958, n47559, 
        n1851, n1886, n1887, n1888, n1889, n1890, n1891, n1892, 
        n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, 
        n1901, n27846, n1917, n1918, n1919, n1920, n1921, n1922, 
        n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, 
        n1931, n1932, n1933, n47553, n1950, n47549, n1985, n1986, 
        n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, 
        n1995, n1996, n1997, n1998, n1999, n2000, n2001, n39646, 
        n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, 
        n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, 
        n2032, n2033, n2049, n47547, n50465, n2084, n2085, n2086, 
        n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, 
        n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2115, 
        n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, 
        n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, 
        n2132, n2133, n39310, n39645, n2148, n39309, n39308, n2183, 
        n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, 
        n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, 
        n2200, n2201, n39644, n39307, n2214, n2215, n2216, n2217, 
        n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, 
        n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, 
        n39306, n2247, n40055, n2281, n2282, n2283, n2284, n2285, 
        n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, 
        n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, 
        n47537, n2313, n2314, n2315, n2316, n2317, n2318, n2319, 
        n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, 
        n2328, n2329, n2330, n2331, n2332, n2333, n50672, n2346, 
        n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, 
        n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, 
        n2397, n2398, n2399, n2400, n2401, n2412, n2413, n2414, 
        n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
        n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, 
        n2431, n2432, n2433, n2445, n27803, n2480, n2481, n2482_adj_4959, 
        n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, 
        n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, 
        n2499, n2500, n2501, n2511, n2512, n2513, n2514, n2515, 
        n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, 
        n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, 
        n2532, n2533, n2544, n47525, n2579, n2580, n2581, n2582, 
        n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, 
        n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, 
        n2599, n2600, n2601, n2610, n2611, n2612, n2613, n2614, 
        n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, 
        n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, 
        n2631, n2632, n2633, n2643, n43659, n2678, n2679, n2680, 
        n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, 
        n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, 
        n2697, n2698, n2699, n2700, n2701, n2709, n2710, n2711, 
        n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, 
        n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, 
        n2728, n2729, n2730, n2731, n2732, n2733, n2742, n2777, 
        n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, 
        n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, 
        n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, 
        n49819, n2808, n2809, n2810, n2811, n2812, n2813, n2814, 
        n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, 
        n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, 
        n2831, n2832, n2833, n49818, n2841, n49817, n47519, n2876, 
        n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, 
        n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, 
        n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, 
        n2901, n2907, n2908, n2909, n2910, n2911, n2912, n2913, 
        n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, 
        n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, 
        n2930, n2931, n2932, n2933, n2940, n2975, n2976, n2977, 
        n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, 
        n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, 
        n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, 
        n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, 
        n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, 
        n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, 
        n3030, n3031, n3032, n3033, n51169, n3039, n3074, n3075, 
        n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, 
        n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, 
        n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, 
        n3100, n3101, n3105, n3106, n3107, n3108, n3109, n3110, 
        n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, 
        n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, 
        n3127, n3128, n3129, n3130, n3131, n3132, n3133, n51241, 
        n3138, n44058, n3173, n3174, n3175, n3176, n3177, n3178, 
        n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, 
        n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, 
        n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3204, 
        n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, 
        n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, 
        n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, 
        n3229, n3230, n3231, n3232, n3233, n51275, n3237, n3272, 
        n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, 
        n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, 
        n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, 
        n3298, n3299, n3300, n3301, n47513, n51546, n27771, n24_adj_4960, 
        n50024, n62, n47507, n39006, n26505, n26508, n39305, n26492, 
        n7_adj_4961, n47501, n47499, n47497, n28221, n47477, n63, 
        n47471, n39304, n39643, n28219, n51137, n4_adj_4962, n6_adj_4963, 
        n7_adj_4964, n8_adj_4965, n9_adj_4966, n10_adj_4967, n11_adj_4968, 
        n12_adj_4969, n13_adj_4970, n15_adj_4971, n17_adj_4972, n19_adj_4973, 
        n21_adj_4974, n50508, n23_adj_4975, n50533, n25_adj_4976, 
        n27_adj_4977, n29_adj_4978, n30_adj_4979, n31_adj_4980, n33_adj_4981, 
        n35, n26490, n40269, n40054, n39642, n39303, n47465, n47463, 
        n28218, n28217, n40053, n47457, n28214, n28213, n47453, 
        n47451, n39641, n50904, n50018, n50783, n50641, n26687, 
        n39302, n47437, n47431, n40052, n49785, n50507, n50013, 
        n50594, n47425, n51102, n47419, n50674, n47415, n39640, 
        n39639, n40051, n40268, n40050, n40049, n50417, n47411, 
        n39638, n50419, n40267, n39301, n5_adj_4982, n7_adj_4983, 
        n45116, n46759, n39637, n47397, n45051, n47391, n45031, 
        n6_adj_4984, n49984, n49982, n4_adj_4985, n47385, n14_adj_4986, 
        n34723, n34617, n47379, n10_adj_4987, n40048, n28211, n8_adj_4988, 
        n28210, n28209, n28208, n28207, n28206, n28205, n28204, 
        n28203, n39636, n47377, n28202, n28200, n28199, n28198, 
        n28194, n39037, n34615, n51637, n61_adj_4989, n65, n39, 
        n47363, n6_adj_4990, n51636, n2_adj_4991, n3_adj_4992, n4_adj_4993, 
        n5_adj_4994, n6_adj_4995, n7_adj_4996, n8_adj_4997, n9_adj_4998, 
        n10_adj_4999, n11_adj_5000, n12_adj_5001, n13_adj_5002, n14_adj_5003, 
        n15_adj_5004, n16_adj_5005, n17_adj_5006, n18_adj_5007, n19_adj_5008, 
        n20_adj_5009, n21_adj_5010, n22_adj_5011, n23_adj_5012, n24_adj_5013, 
        n25_adj_5014, n26_adj_5015, n27_adj_5016, n28_adj_5017, n29_adj_5018, 
        n30_adj_5019, n31_adj_5020, n32_adj_5021, n33_adj_5022, n45073, 
        n39635, n47357, n39300, n39634, n39633, n8_adj_5023, n45111, 
        n7_adj_5024, n39632, n34611, n39299, n47351, n40266, n39298, 
        n39297, n39296, n45134, n47345, n39036, n39005, n34607, 
        n4_adj_5025, n34603, n40047, n39295, n39294, n34599, n40265, 
        n39035, n47333, n45109, n39631, n40046, n39004, n39034, 
        n40264, n40263, n40045, n39003, n44436, n34593, n40044, 
        n40043, n40262, n34591, n45125, n40042, n40261, n40041, 
        n40040, n39293, n44035, n39033, n39292, n40039, n40038, 
        n39291, n40260, n44685, n34631, n47327, n40259, n34583, 
        n40258, n40257, n39002, n39290, n39032, n39031, n40256, 
        n43485, n40255, n47321, n39030, n38993, n34675, n47317, 
        n38992, n39289, n39029, n6_adj_5026, n39288, n40254, n39287, 
        n40253, n39819, n39818, n39286, n40252, n39817, n40251, 
        n39816, n39285, n40250, n40249, n39284, n39815, n39814, 
        n40248, n40247, n40246, n39028, n39813, n39812, n39811, 
        n38991, n39283, n39282, n39810, n39809, n39027, n39808, 
        n39281, n39280, n39279, n40245, n15_adj_5027, n17_adj_5028, 
        n19_adj_5029, n39026, n27_adj_5030, n29_adj_5031, n39025, 
        n33_adj_5032, n39024, n37, n41, n39023, n39022, n59, n61_adj_5033, 
        n40244, n50506, n47311, n44048, n47297, n47291, n47287, 
        n51390, n48793, n47269, n47263, n8_adj_5034, n7_adj_5035, 
        n40_adj_5036, n51356, n8_adj_5037, n51327, n40243, n47253, 
        n5_adj_5038, n39807, n39806, n47247, n39805, n40242, n50531, 
        n10_adj_5039, n47239, n26624, n40241, n47229, n40240, n40239, 
        n50273, n50283, n39804, n40238, n50832, n47219, n23831, 
        n26603, n26881, n47213, n40237, n51045, n40236, n10_adj_5040, 
        n50673, n47203, n46246, n39803, n49758, n47197, n40235, 
        n40234, n39802, n39021, n47191, n47185, n47181, n51019, 
        n47179, n47167, n40233, n46845, n47159, n47157, n34541, 
        n48729, n47151, n40232, n39020, n47145, n47139, n39019, 
        n50740, n47133, n39018, n47127, n47121, n47119, n50998, 
        n45131, n45146, n40231, n44240, n40230, n47105, n28189, 
        n34531, n40229, n39801, n49734, n6_adj_5041, n39800, n40228, 
        n40227, n39799, n40226, n39798, n39797, n47099, n50505, 
        n40225, n39796, n39795, n47093, n47087, n47081, n40224, 
        n47079, n47077, n39794, n34525, n39001, n5_adj_5042, n39793, 
        n39792, n38990, n39791, n39017, n47059, n46808, n39000, 
        n47053, n47051, n39016, n40223, n47045, n47043, n40222, 
        n40221, n47033, n39015, n39790, n38999, n26629, n26502, 
        n47027, n28188, n47025, n40220, n40219, n39789, n39788, 
        n40218, n14_adj_5043, n50817, n44813, n44811, n44809, n47019, 
        n44807, n50560, n40217, n39787, n39786, n44804, n39785, 
        n47017, n39784, n26650, n47003, n40216, n39783, n47001, 
        n45435, n46999, n40215, n46997, n49726, n46995, n39014, 
        n46993, n23935, n50974, n46991, n38998, n46989, n46987, 
        n40214, n40213, n46983, n46981, n46977, n46969, n46967, 
        n46965, n39782, n49724, n39781, n46963, n46961, n10_adj_5044, 
        n40212, n46959, n46953, n46943, n33769, n39780, n46937, 
        n46931, n46929, n46921, n40211, n46915, n43968, n51409, 
        n46909, n27546, n46903, n45042, n40210, n45023, n46899, 
        n39779, n46895, n26484, n26483, n49714, n50955;
    
    VCC i2 (.Y(VCC_net));
    SB_DFF encoder0_position_scaled_i0 (.Q(encoder0_position_scaled[0]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[0]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_IO hall2_input (.PACKAGE_PIN(HALL2), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall2)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall2_input.PIN_TYPE = 6'b000001;
    defparam hall2_input.PULLUP = 1'b1;
    defparam hall2_input.NEG_TRIGGER = 1'b0;
    defparam hall2_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO hall3_input (.PACKAGE_PIN(HALL3), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall3)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall3_input.PIN_TYPE = 6'b000001;
    defparam hall3_input.PULLUP = 1'b1;
    defparam hall3_input.NEG_TRIGGER = 1'b0;
    defparam hall3_input.IO_STANDARD = "SB_LVCMOS";
    SB_IO tx_output (.PACKAGE_PIN(TX), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(tx_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(tx_o)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam tx_output.PIN_TYPE = 6'b101001;
    defparam tx_output.PULLUP = 1'b1;
    defparam tx_output.NEG_TRIGGER = 1'b0;
    defparam tx_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF h3_58 (.Q(INLB_c), .C(CLK_c), .D(hall3));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 encoder0_position_31__I_0_add_833_11_lut (.I0(GND_net), .I1(n1225), 
            .I2(VCC_net), .I3(n39673), .O(n1292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_11_lut.LUT_INIT = 16'hC33C;
    SB_DFF encoder1_position_scaled_i0 (.Q(encoder1_position_scaled[0]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[0]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_IO sda_output (.PACKAGE_PIN(SDA), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(sda_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(sda_out), .D_IN_0(state_7__N_4003[3])) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam sda_output.PIN_TYPE = 6'b101001;
    defparam sda_output.PULLUP = 1'b1;
    defparam sda_output.NEG_TRIGGER = 1'b0;
    defparam sda_output.IO_STANDARD = "SB_LVCMOS";
    SB_DFF displacement_i0 (.Q(displacement[0]), .C(CLK_c), .D(displacement_23__N_82[0]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_IO CS_pad (.PACKAGE_PIN(CS), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_pad.PIN_TYPE = 6'b011001;
    defparam CS_pad.PULLUP = 1'b0;
    defparam CS_pad.NEG_TRIGGER = 1'b0;
    defparam CS_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 i36066_1_lut (.I0(n1950), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51019));
    defparam i36066_1_lut.LUT_INIT = 16'h5555;
    SB_IO scl_output (.PACKAGE_PIN(SCL), .LATCH_INPUT_VALUE(GND_net), .INPUT_CLK(GND_net), 
          .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(scl_enable), .D_OUT_1(GND_net), 
          .D_OUT_0(scl)) /* synthesis syn_instantiated=1 */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam scl_output.PIN_TYPE = 6'b101001;
    defparam scl_output.PULLUP = 1'b1;
    defparam scl_output.NEG_TRIGGER = 1'b0;
    defparam scl_output.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_31__I_0_add_833_11 (.CI(n39673), .I0(n1225), 
            .I1(VCC_net), .CO(n39674));
    SB_DFF h2_57 (.Q(INHB_c), .C(CLK_c), .D(hall2));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_IO hall1_input (.PACKAGE_PIN(HALL1), .LATCH_INPUT_VALUE(GND_net), 
          .INPUT_CLK(GND_net), .OUTPUT_CLK(GND_net), .OUTPUT_ENABLE(GND_net), 
          .D_OUT_1(GND_net), .D_OUT_0(GND_net), .D_IN_0(hall1)) /* synthesis syn_instantiated=1, IO_FF_IN=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam hall1_input.PIN_TYPE = 6'b000001;
    defparam hall1_input.PULLUP = 1'b1;
    defparam hall1_input.NEG_TRIGGER = 1'b0;
    defparam hall1_input.IO_STANDARD = "SB_LVCMOS";
    \neopixel(CLOCK_SPEED_HZ=16000000)  nx (.n28315(n28315), .\neo_pixel_transmitter.t0 ({\neo_pixel_transmitter.t0 }), 
            .CLK_c(CLK_c), .n28314(n28314), .n28313(n28313), .n28312(n28312), 
            .VCC_net(VCC_net), .GND_net(GND_net), .\neo_pixel_transmitter.done (\neo_pixel_transmitter.done ), 
            .n28311(n28311), .n28310(n28310), .n28309(n28309), .\state[0] (state[0]), 
            .n34525(n34525), .\state[1] (state[1]), .n28308(n28308), .timer({timer}), 
            .n28307(n28307), .n28306(n28306), .n28305(n28305), .n28304(n28304), 
            .n28303(n28303), .n28302(n28302), .n28301(n28301), .n28300(n28300), 
            .n28299(n28299), .n28298(n28298), .n28297(n28297), .n28296(n28296), 
            .n28295(n28295), .n28294(n28294), .n28293(n28293), .n28292(n28292), 
            .n28291(n28291), .n28290(n28290), .n28289(n28289), .n28288(n28288), 
            .n28287(n28287), .n28286(n28286), .n28285(n28285), .\state_3__N_428[1] (state_3__N_428[1]), 
            .LED_c(LED_c), .n34629(n34629), .n44839(n44839), .n27916(n27916), 
            .neopxl_color({neopxl_color}), .start(start), .n43085(n43085), 
            .n42985(n42985), .n28194(n28194), .n28188(n28188), .NEOPXL_c(NEOPXL_c)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(43[24] 49[2])
    SB_CARRY encoder0_position_31__I_0_add_1302_9 (.CI(n39772), .I0(n1927), 
            .I1(VCC_net), .CO(n39773));
    SB_LUT4 encoder0_position_31__I_0_add_1302_8_lut (.I0(GND_net), .I1(n1928), 
            .I2(VCC_net), .I3(n39771), .O(n1995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_833_10_lut (.I0(GND_net), .I1(n1226), 
            .I2(VCC_net), .I3(n39672), .O(n1293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_10_lut.LUT_INIT = 16'hC33C;
    SB_DFF dir_62 (.Q(INHC_c), .C(CLK_c), .D(duty[23]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 i35879_1_lut (.I0(n1356), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50832));
    defparam i35879_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_83_i19_4_lut (.I0(encoder1_position_scaled[18]), .I1(displacement[18]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[18]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i19_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i20_1_lut (.I0(encoder1_position_scaled[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4892));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_83_i20_4_lut (.I0(encoder1_position_scaled[19]), .I1(displacement[19]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[19]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i20_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_31__I_0_add_833_10 (.CI(n39672), .I0(n1226), 
            .I1(VCC_net), .CO(n39673));
    SB_LUT4 encoder0_position_31__I_0_i1249_3_lut (.I0(n1830), .I1(n1897), 
            .I2(n1851), .I3(GND_net), .O(n1929));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36092_1_lut (.I0(n2049), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51045));
    defparam i36092_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1302_8 (.CI(n39771), .I0(n1928), 
            .I1(VCC_net), .CO(n39772));
    SB_LUT4 encoder0_position_31__I_0_add_1302_7_lut (.I0(GND_net), .I1(n1929), 
            .I2(GND_net), .I3(n39770), .O(n1996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_833_9_lut (.I0(GND_net), .I1(n1227), 
            .I2(VCC_net), .I3(n39671), .O(n1294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35951_1_lut (.I0(n1455), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50904));
    defparam i35951_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1302_7 (.CI(n39770), .I0(n1929), 
            .I1(GND_net), .CO(n39771));
    SB_LUT4 encoder0_position_31__I_0_add_1302_6_lut (.I0(GND_net), .I1(n1930), 
            .I2(GND_net), .I3(n39769), .O(n1997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n62), .I2(delay_counter[31]), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n46845));
    defparam i3_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i15167_4_lut (.I0(state_7__N_4003[3]), .I1(data[0]), .I2(n10_adj_5039), 
            .I3(n26645), .O(n28230));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15167_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15245_3_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(timer[8]), 
            .I2(n43085), .I3(GND_net), .O(n28308));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15245_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i21_1_lut (.I0(encoder1_position_scaled[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4891));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36374_1_lut (.I0(n2346), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51327));
    defparam i36374_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_833_9 (.CI(n39671), .I0(n1227), 
            .I1(VCC_net), .CO(n39672));
    SB_LUT4 encoder0_position_31__I_0_add_833_8_lut (.I0(GND_net), .I1(n1228), 
            .I2(VCC_net), .I3(n39670), .O(n1295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_6 (.CI(n39769), .I0(n1930), 
            .I1(GND_net), .CO(n39770));
    SB_LUT4 mux_83_i21_4_lut (.I0(encoder1_position_scaled[20]), .I1(displacement[20]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[20]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i21_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY encoder0_position_31__I_0_add_833_8 (.CI(n39670), .I0(n1228), 
            .I1(VCC_net), .CO(n39671));
    SB_LUT4 mux_83_i22_4_lut (.I0(encoder1_position_scaled[21]), .I1(displacement[21]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[21]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i22_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i22_1_lut (.I0(encoder1_position_scaled[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4937));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_83_i23_4_lut (.I0(encoder1_position_scaled[22]), .I1(displacement[22]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[22]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i23_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_add_833_7_lut (.I0(GND_net), .I1(n1229), 
            .I2(GND_net), .I3(n39669), .O(n1296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut (.I0(control_mode[3]), .I1(control_mode[5]), .I2(control_mode[4]), 
            .I3(control_mode[7]), .O(n10_adj_5040));   // verilog/TinyFPGA_B.v(169[5:22])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut (.I0(control_mode[6]), .I1(n10_adj_5040), .I2(control_mode[2]), 
            .I3(GND_net), .O(n26603));   // verilog/TinyFPGA_B.v(169[5:22])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut (.I0(n26480), .I1(control_mode[1]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4885));   // verilog/TinyFPGA_B.v(170[5:22])
    defparam i1_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_3_lut (.I0(control_mode[0]), .I1(control_mode[1]), .I2(n26603), 
            .I3(GND_net), .O(n15));   // verilog/TinyFPGA_B.v(169[5:22])
    defparam i2_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 mux_83_i24_4_lut (.I0(encoder1_position_scaled[23]), .I1(displacement[23]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[23]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i24_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i23_1_lut (.I0(encoder1_position_scaled[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4936));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1302_5_lut (.I0(GND_net), .I1(n1931), 
            .I2(VCC_net), .I3(n39768), .O(n1998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_833_7 (.CI(n39669), .I0(n1229), 
            .I1(GND_net), .CO(n39670));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i24_3_lut (.I0(encoder0_position[23]), 
            .I1(n10_adj_4932), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n935));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i24_1_lut (.I0(encoder1_position_scaled[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR delay_counter_i0_i31 (.Q(delay_counter[31]), .C(CLK_c), .E(n5722), 
            .D(n659), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 i36403_1_lut (.I0(n2445), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51356));
    defparam i36403_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i25_3_lut (.I0(encoder0_position[24]), 
            .I1(n9_adj_4933), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n934));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i25_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i641_3_lut (.I0(n934), .I1(n1001), 
            .I2(n960), .I3(GND_net), .O(n1033));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i573_3_lut (.I0(n834), .I1(n901), 
            .I2(n861), .I3(GND_net), .O(n933));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i573_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i640_3_lut (.I0(n933), .I1(n1000), 
            .I2(n960), .I3(GND_net), .O(n1032));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_833_6_lut (.I0(GND_net), .I1(n1230), 
            .I2(GND_net), .I3(n39668), .O(n1297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut (.I0(n34334), .I1(n44120), .I2(state_adj_5100[0]), 
            .I3(read), .O(n43685));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut.LUT_INIT = 16'h8280;
    SB_CARRY encoder0_position_31__I_0_add_1302_5 (.CI(n39768), .I0(n1931), 
            .I1(VCC_net), .CO(n39769));
    SB_LUT4 encoder0_position_31__I_0_add_1302_4_lut (.I0(GND_net), .I1(n1932), 
            .I2(GND_net), .I3(n39767), .O(n1999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15430_3_lut (.I0(neopxl_color[23]), .I1(\data_in_frame[4] [7]), 
            .I2(n46360), .I3(GND_net), .O(n28493));   // verilog/coms.v(127[12] 300[6])
    defparam i15430_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15431_3_lut (.I0(neopxl_color[22]), .I1(\data_in_frame[4] [6]), 
            .I2(n46360), .I3(GND_net), .O(n28494));   // verilog/coms.v(127[12] 300[6])
    defparam i15431_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_833_6 (.CI(n39668), .I0(n1230), 
            .I1(GND_net), .CO(n39669));
    SB_LUT4 i15432_3_lut (.I0(neopxl_color[21]), .I1(\data_in_frame[4] [5]), 
            .I2(n46360), .I3(GND_net), .O(n28495));   // verilog/coms.v(127[12] 300[6])
    defparam i15432_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i30 (.Q(delay_counter[30]), .C(CLK_c), .E(n5722), 
            .D(n660), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 i15433_3_lut (.I0(neopxl_color[20]), .I1(\data_in_frame[4] [4]), 
            .I2(n46360), .I3(GND_net), .O(n28496));   // verilog/coms.v(127[12] 300[6])
    defparam i15433_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_833_5_lut (.I0(GND_net), .I1(n1231), 
            .I2(VCC_net), .I3(n39667), .O(n1298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15434_3_lut (.I0(neopxl_color[19]), .I1(\data_in_frame[4] [3]), 
            .I2(n46360), .I3(GND_net), .O(n28497));   // verilog/coms.v(127[12] 300[6])
    defparam i15434_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15435_3_lut (.I0(neopxl_color[18]), .I1(\data_in_frame[4] [2]), 
            .I2(n46360), .I3(GND_net), .O(n28498));   // verilog/coms.v(127[12] 300[6])
    defparam i15435_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15436_3_lut (.I0(neopxl_color[17]), .I1(\data_in_frame[4] [1]), 
            .I2(n46360), .I3(GND_net), .O(n28499));   // verilog/coms.v(127[12] 300[6])
    defparam i15436_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1302_4 (.CI(n39767), .I0(n1932), 
            .I1(GND_net), .CO(n39768));
    SB_LUT4 i15437_3_lut (.I0(neopxl_color[16]), .I1(\data_in_frame[4] [0]), 
            .I2(n46360), .I3(GND_net), .O(n28500));   // verilog/coms.v(127[12] 300[6])
    defparam i15437_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15438_3_lut (.I0(neopxl_color[15]), .I1(\data_in_frame[5] [7]), 
            .I2(n46360), .I3(GND_net), .O(n28501));   // verilog/coms.v(127[12] 300[6])
    defparam i15438_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15439_3_lut (.I0(neopxl_color[14]), .I1(\data_in_frame[5] [6]), 
            .I2(n46360), .I3(GND_net), .O(n28502));   // verilog/coms.v(127[12] 300[6])
    defparam i15439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15440_3_lut (.I0(neopxl_color[13]), .I1(\data_in_frame[5] [5]), 
            .I2(n46360), .I3(GND_net), .O(n28503));   // verilog/coms.v(127[12] 300[6])
    defparam i15440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15441_3_lut (.I0(neopxl_color[12]), .I1(\data_in_frame[5] [4]), 
            .I2(n46360), .I3(GND_net), .O(n28504));   // verilog/coms.v(127[12] 300[6])
    defparam i15441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15442_3_lut (.I0(neopxl_color[11]), .I1(\data_in_frame[5] [3]), 
            .I2(n46360), .I3(GND_net), .O(n28505));   // verilog/coms.v(127[12] 300[6])
    defparam i15442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15443_3_lut (.I0(neopxl_color[10]), .I1(\data_in_frame[5] [2]), 
            .I2(n46360), .I3(GND_net), .O(n28506));   // verilog/coms.v(127[12] 300[6])
    defparam i15443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15444_3_lut (.I0(neopxl_color[9]), .I1(\data_in_frame[5] [1]), 
            .I2(n46360), .I3(GND_net), .O(n28507));   // verilog/coms.v(127[12] 300[6])
    defparam i15444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15445_3_lut (.I0(neopxl_color[8]), .I1(\data_in_frame[5] [0]), 
            .I2(n46360), .I3(GND_net), .O(n28508));   // verilog/coms.v(127[12] 300[6])
    defparam i15445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15446_3_lut (.I0(neopxl_color[7]), .I1(\data_in_frame[6] [7]), 
            .I2(n46360), .I3(GND_net), .O(n28509));   // verilog/coms.v(127[12] 300[6])
    defparam i15446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15447_3_lut (.I0(neopxl_color[6]), .I1(\data_in_frame[6] [6]), 
            .I2(n46360), .I3(GND_net), .O(n28510));   // verilog/coms.v(127[12] 300[6])
    defparam i15447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15448_3_lut (.I0(neopxl_color[5]), .I1(\data_in_frame[6] [5]), 
            .I2(n46360), .I3(GND_net), .O(n28511));   // verilog/coms.v(127[12] 300[6])
    defparam i15448_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15449_3_lut (.I0(neopxl_color[4]), .I1(\data_in_frame[6] [4]), 
            .I2(n46360), .I3(GND_net), .O(n28512));   // verilog/coms.v(127[12] 300[6])
    defparam i15449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15450_3_lut (.I0(neopxl_color[3]), .I1(\data_in_frame[6] [3]), 
            .I2(n46360), .I3(GND_net), .O(n28513));   // verilog/coms.v(127[12] 300[6])
    defparam i15450_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15451_3_lut (.I0(neopxl_color[2]), .I1(\data_in_frame[6] [2]), 
            .I2(n46360), .I3(GND_net), .O(n28514));   // verilog/coms.v(127[12] 300[6])
    defparam i15451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15452_3_lut (.I0(neopxl_color[1]), .I1(\data_in_frame[6] [1]), 
            .I2(n46360), .I3(GND_net), .O(n28515));   // verilog/coms.v(127[12] 300[6])
    defparam i15452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i26_3_lut (.I0(encoder0_position[25]), 
            .I1(n8_adj_4934), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n834));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i26_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15453_3_lut (.I0(\data_out_frame[25] [7]), .I1(neopxl_color[7]), 
            .I2(n23935), .I3(GND_net), .O(n28516));   // verilog/coms.v(127[12] 300[6])
    defparam i15453_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15454_3_lut (.I0(\data_out_frame[25] [6]), .I1(neopxl_color[6]), 
            .I2(n23935), .I3(GND_net), .O(n28517));   // verilog/coms.v(127[12] 300[6])
    defparam i15454_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15455_3_lut (.I0(\data_out_frame[25] [5]), .I1(neopxl_color[5]), 
            .I2(n23935), .I3(GND_net), .O(n28518));   // verilog/coms.v(127[12] 300[6])
    defparam i15455_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15456_3_lut (.I0(\data_out_frame[25] [4]), .I1(neopxl_color[4]), 
            .I2(n23935), .I3(GND_net), .O(n28519));   // verilog/coms.v(127[12] 300[6])
    defparam i15456_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15457_3_lut (.I0(\data_out_frame[25] [3]), .I1(neopxl_color[3]), 
            .I2(n23935), .I3(GND_net), .O(n28520));   // verilog/coms.v(127[12] 300[6])
    defparam i15457_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15458_3_lut (.I0(\data_out_frame[25] [2]), .I1(neopxl_color[2]), 
            .I2(n23935), .I3(GND_net), .O(n28521));   // verilog/coms.v(127[12] 300[6])
    defparam i15458_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15125_3_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(timer[0]), 
            .I2(n43085), .I3(GND_net), .O(n28188));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15125_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15126_3_lut (.I0(IntegralLimit[0]), .I1(\data_in_frame[13] [0]), 
            .I2(n27771), .I3(GND_net), .O(n28189));   // verilog/coms.v(127[12] 300[6])
    defparam i15126_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15131_4_lut (.I0(n44839), .I1(state[1]), .I2(state_3__N_428[1]), 
            .I3(n27916), .O(n28194));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15131_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i15459_3_lut (.I0(\data_out_frame[25] [1]), .I1(neopxl_color[1]), 
            .I2(n23935), .I3(GND_net), .O(n28522));   // verilog/coms.v(127[12] 300[6])
    defparam i15459_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15460_3_lut (.I0(\data_out_frame[25] [0]), .I1(neopxl_color[0]), 
            .I2(n23935), .I3(GND_net), .O(n28523));   // verilog/coms.v(127[12] 300[6])
    defparam i15460_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15461_3_lut (.I0(\data_out_frame[24] [7]), .I1(neopxl_color[15]), 
            .I2(n23935), .I3(GND_net), .O(n28524));   // verilog/coms.v(127[12] 300[6])
    defparam i15461_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15462_3_lut (.I0(\data_out_frame[24] [6]), .I1(neopxl_color[14]), 
            .I2(n23935), .I3(GND_net), .O(n28525));   // verilog/coms.v(127[12] 300[6])
    defparam i15462_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15463_3_lut (.I0(\data_out_frame[24] [5]), .I1(neopxl_color[13]), 
            .I2(n23935), .I3(GND_net), .O(n28526));   // verilog/coms.v(127[12] 300[6])
    defparam i15463_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15464_3_lut (.I0(\data_out_frame[24] [4]), .I1(neopxl_color[12]), 
            .I2(n23935), .I3(GND_net), .O(n28527));   // verilog/coms.v(127[12] 300[6])
    defparam i15464_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15465_3_lut (.I0(\data_out_frame[24] [3]), .I1(neopxl_color[11]), 
            .I2(n23935), .I3(GND_net), .O(n28528));   // verilog/coms.v(127[12] 300[6])
    defparam i15465_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15135_4_lut (.I0(state_7__N_4003[3]), .I1(data[7]), .I2(n33769), 
            .I3(n26650), .O(n28198));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15135_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15136_4_lut (.I0(state_7__N_4003[3]), .I1(data[6]), .I2(n33769), 
            .I3(n26645), .O(n28199));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15136_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15137_4_lut (.I0(state_7__N_4003[3]), .I1(data[5]), .I2(n4_adj_4915), 
            .I3(n26650), .O(n28200));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15137_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15139_4_lut (.I0(r_Rx_Data), .I1(rx_data[1]), .I2(n4_adj_4938), 
            .I3(n26624), .O(n28202));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15139_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15466_3_lut (.I0(\data_out_frame[24] [2]), .I1(neopxl_color[10]), 
            .I2(n23935), .I3(GND_net), .O(n28529));   // verilog/coms.v(127[12] 300[6])
    defparam i15466_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15467_3_lut (.I0(\data_out_frame[24] [1]), .I1(neopxl_color[9]), 
            .I2(n23935), .I3(GND_net), .O(n28530));   // verilog/coms.v(127[12] 300[6])
    defparam i15467_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15468_3_lut (.I0(\data_out_frame[24] [0]), .I1(neopxl_color[8]), 
            .I2(n23935), .I3(GND_net), .O(n28531));   // verilog/coms.v(127[12] 300[6])
    defparam i15468_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15469_3_lut (.I0(\data_out_frame[23] [7]), .I1(neopxl_color[23]), 
            .I2(n23935), .I3(GND_net), .O(n28532));   // verilog/coms.v(127[12] 300[6])
    defparam i15469_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15470_3_lut (.I0(\data_out_frame[23] [6]), .I1(neopxl_color[22]), 
            .I2(n23935), .I3(GND_net), .O(n28533));   // verilog/coms.v(127[12] 300[6])
    defparam i15470_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15471_3_lut (.I0(\data_out_frame[23] [5]), .I1(neopxl_color[21]), 
            .I2(n23935), .I3(GND_net), .O(n28534));   // verilog/coms.v(127[12] 300[6])
    defparam i15471_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15472_3_lut (.I0(\data_out_frame[23] [4]), .I1(neopxl_color[20]), 
            .I2(n23935), .I3(GND_net), .O(n28535));   // verilog/coms.v(127[12] 300[6])
    defparam i15472_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15473_3_lut (.I0(\data_out_frame[23] [3]), .I1(neopxl_color[19]), 
            .I2(n23935), .I3(GND_net), .O(n28536));   // verilog/coms.v(127[12] 300[6])
    defparam i15473_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15187_4_lut (.I0(r_Rx_Data), .I1(rx_data[0]), .I2(n4_adj_4938), 
            .I3(n26629), .O(n28250));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15187_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15474_3_lut (.I0(\data_out_frame[23] [2]), .I1(neopxl_color[18]), 
            .I2(n23935), .I3(GND_net), .O(n28537));   // verilog/coms.v(127[12] 300[6])
    defparam i15474_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15475_3_lut (.I0(\data_out_frame[23] [1]), .I1(neopxl_color[17]), 
            .I2(n23935), .I3(GND_net), .O(n28538));   // verilog/coms.v(127[12] 300[6])
    defparam i15475_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15476_3_lut (.I0(\data_out_frame[23] [0]), .I1(neopxl_color[16]), 
            .I2(n23935), .I3(GND_net), .O(n28539));   // verilog/coms.v(127[12] 300[6])
    defparam i15476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15477_3_lut (.I0(\data_out_frame[20] [7]), .I1(displacement[7]), 
            .I2(n23935), .I3(GND_net), .O(n28540));   // verilog/coms.v(127[12] 300[6])
    defparam i15477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15478_3_lut (.I0(\data_out_frame[20] [6]), .I1(displacement[6]), 
            .I2(n23935), .I3(GND_net), .O(n28541));   // verilog/coms.v(127[12] 300[6])
    defparam i15478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15479_3_lut (.I0(\data_out_frame[20] [5]), .I1(displacement[5]), 
            .I2(n23935), .I3(GND_net), .O(n28542));   // verilog/coms.v(127[12] 300[6])
    defparam i15479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15480_3_lut (.I0(\data_out_frame[20] [4]), .I1(displacement[4]), 
            .I2(n23935), .I3(GND_net), .O(n28543));   // verilog/coms.v(127[12] 300[6])
    defparam i15480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15183_4_lut (.I0(n27846), .I1(r_Bit_Index[0]), .I2(n43968), 
            .I3(r_SM_Main[1]), .O(n28246));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15183_4_lut.LUT_INIT = 16'h4644;
    SB_LUT4 i15481_3_lut (.I0(\data_out_frame[20] [3]), .I1(displacement[3]), 
            .I2(n23935), .I3(GND_net), .O(n28544));   // verilog/coms.v(127[12] 300[6])
    defparam i15481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15482_3_lut (.I0(\data_out_frame[20] [2]), .I1(displacement[2]), 
            .I2(n23935), .I3(GND_net), .O(n28545));   // verilog/coms.v(127[12] 300[6])
    defparam i15482_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15483_3_lut (.I0(\data_out_frame[20] [1]), .I1(displacement[1]), 
            .I2(n23935), .I3(GND_net), .O(n28546));   // verilog/coms.v(127[12] 300[6])
    defparam i15483_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17199_3_lut (.I0(\data_out_frame[20] [0]), .I1(displacement[0]), 
            .I2(n23935), .I3(GND_net), .O(n28547));
    defparam i17199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1674 (.I0(n771), .I1(n63), .I2(n74), .I3(n8_adj_5037), 
            .O(n5_adj_5038));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1674.LUT_INIT = 16'hcc04;
    SB_LUT4 i3_4_lut_adj_1675 (.I0(n7_adj_4983), .I1(n5_adj_4982), .I2(n51904), 
            .I3(n46759), .O(n8_adj_4988));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1675.LUT_INIT = 16'heefe;
    SB_LUT4 i4_4_lut_adj_1676 (.I0(n29985), .I1(n8_adj_4988), .I2(n76), 
            .I3(n5_adj_5038), .O(n51637));   // verilog/coms.v(127[12] 300[6])
    defparam i4_4_lut_adj_1676.LUT_INIT = 16'hefcf;
    SB_LUT4 i15485_3_lut (.I0(\data_out_frame[19] [7]), .I1(displacement[15]), 
            .I2(n23935), .I3(GND_net), .O(n28548));   // verilog/coms.v(127[12] 300[6])
    defparam i15485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15486_3_lut (.I0(\data_out_frame[19] [6]), .I1(displacement[14]), 
            .I2(n23935), .I3(GND_net), .O(n28549));   // verilog/coms.v(127[12] 300[6])
    defparam i15486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15487_3_lut (.I0(\data_out_frame[19] [5]), .I1(displacement[13]), 
            .I2(n23935), .I3(GND_net), .O(n28550));   // verilog/coms.v(127[12] 300[6])
    defparam i15487_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_833_5 (.CI(n39667), .I0(n1231), 
            .I1(VCC_net), .CO(n39668));
    SB_LUT4 i15488_3_lut (.I0(\data_out_frame[19] [4]), .I1(displacement[12]), 
            .I2(n23935), .I3(GND_net), .O(n28551));   // verilog/coms.v(127[12] 300[6])
    defparam i15488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15489_3_lut (.I0(\data_out_frame[19] [3]), .I1(displacement[11]), 
            .I2(n23935), .I3(GND_net), .O(n28552));   // verilog/coms.v(127[12] 300[6])
    defparam i15489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15490_3_lut (.I0(\data_out_frame[19] [2]), .I1(displacement[10]), 
            .I2(n23935), .I3(GND_net), .O(n28553));   // verilog/coms.v(127[12] 300[6])
    defparam i15490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15491_3_lut (.I0(\data_out_frame[19] [1]), .I1(displacement[9]), 
            .I2(n23935), .I3(GND_net), .O(n28554));   // verilog/coms.v(127[12] 300[6])
    defparam i15491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15492_3_lut (.I0(\data_out_frame[19] [0]), .I1(displacement[8]), 
            .I2(n23935), .I3(GND_net), .O(n28555));   // verilog/coms.v(127[12] 300[6])
    defparam i15492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1677 (.I0(n44092), .I1(\FRAME_MATCHER.i_31__N_2526 ), 
            .I2(n26687), .I3(\FRAME_MATCHER.i [31]), .O(n4_adj_5025));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1677.LUT_INIT = 16'heeae;
    SB_LUT4 i70_4_lut (.I0(n2482), .I1(n1476), .I2(n33302), .I3(n44058), 
            .O(n65));   // verilog/coms.v(127[12] 300[6])
    defparam i70_4_lut.LUT_INIT = 16'h5c0c;
    SB_LUT4 i1_4_lut_adj_1678 (.I0(n65), .I1(n39), .I2(n4_adj_5025), .I3(n63), 
            .O(n61_adj_4989));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1678.LUT_INIT = 16'hc8fa;
    SB_LUT4 i2_4_lut (.I0(n61_adj_4989), .I1(\FRAME_MATCHER.i [31]), .I2(n26489), 
            .I3(\FRAME_MATCHER.i_31__N_2524 ), .O(n6_adj_4990));   // verilog/coms.v(127[12] 300[6])
    defparam i2_4_lut.LUT_INIT = 16'hbaaa;
    SB_LUT4 i3_4_lut_adj_1679 (.I0(n76), .I1(n6_adj_4990), .I2(n74), .I3(n771), 
            .O(n51636));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1679.LUT_INIT = 16'hdfdd;
    SB_LUT4 i15192_3_lut (.I0(PWMLimit[23]), .I1(\data_in_frame[8] [7]), 
            .I2(n27771), .I3(GND_net), .O(n28255));   // verilog/coms.v(127[12] 300[6])
    defparam i15192_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15193_3_lut (.I0(PWMLimit[22]), .I1(\data_in_frame[8] [6]), 
            .I2(n27771), .I3(GND_net), .O(n28256));   // verilog/coms.v(127[12] 300[6])
    defparam i15193_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15194_3_lut (.I0(PWMLimit[21]), .I1(\data_in_frame[8] [5]), 
            .I2(n27771), .I3(GND_net), .O(n28257));   // verilog/coms.v(127[12] 300[6])
    defparam i15194_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15195_3_lut (.I0(PWMLimit[20]), .I1(\data_in_frame[8] [4]), 
            .I2(n27771), .I3(GND_net), .O(n28258));   // verilog/coms.v(127[12] 300[6])
    defparam i15195_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15196_3_lut (.I0(PWMLimit[19]), .I1(\data_in_frame[8] [3]), 
            .I2(n27771), .I3(GND_net), .O(n28259));   // verilog/coms.v(127[12] 300[6])
    defparam i15196_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15197_3_lut (.I0(PWMLimit[18]), .I1(\data_in_frame[8] [2]), 
            .I2(n27771), .I3(GND_net), .O(n28260));   // verilog/coms.v(127[12] 300[6])
    defparam i15197_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15198_3_lut (.I0(PWMLimit[17]), .I1(\data_in_frame[8] [1]), 
            .I2(n27771), .I3(GND_net), .O(n28261));   // verilog/coms.v(127[12] 300[6])
    defparam i15198_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15199_3_lut (.I0(PWMLimit[16]), .I1(\data_in_frame[8] [0]), 
            .I2(n27771), .I3(GND_net), .O(n28262));   // verilog/coms.v(127[12] 300[6])
    defparam i15199_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15493_3_lut (.I0(\data_out_frame[18] [7]), .I1(displacement[23]), 
            .I2(n23935), .I3(GND_net), .O(n28556));   // verilog/coms.v(127[12] 300[6])
    defparam i15493_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15494_3_lut (.I0(\data_out_frame[18] [6]), .I1(displacement[22]), 
            .I2(n23935), .I3(GND_net), .O(n28557));   // verilog/coms.v(127[12] 300[6])
    defparam i15494_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15200_3_lut (.I0(PWMLimit[15]), .I1(\data_in_frame[9] [7]), 
            .I2(n27771), .I3(GND_net), .O(n28263));   // verilog/coms.v(127[12] 300[6])
    defparam i15200_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15201_3_lut (.I0(PWMLimit[14]), .I1(\data_in_frame[9] [6]), 
            .I2(n27771), .I3(GND_net), .O(n28264));   // verilog/coms.v(127[12] 300[6])
    defparam i15201_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15202_3_lut (.I0(PWMLimit[13]), .I1(\data_in_frame[9] [5]), 
            .I2(n27771), .I3(GND_net), .O(n28265));   // verilog/coms.v(127[12] 300[6])
    defparam i15202_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15203_3_lut (.I0(PWMLimit[12]), .I1(\data_in_frame[9] [4]), 
            .I2(n27771), .I3(GND_net), .O(n28266));   // verilog/coms.v(127[12] 300[6])
    defparam i15203_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15495_3_lut (.I0(\data_out_frame[18] [5]), .I1(displacement[21]), 
            .I2(n23935), .I3(GND_net), .O(n28558));   // verilog/coms.v(127[12] 300[6])
    defparam i15495_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15496_3_lut (.I0(\data_out_frame[18] [4]), .I1(displacement[20]), 
            .I2(n23935), .I3(GND_net), .O(n28559));   // verilog/coms.v(127[12] 300[6])
    defparam i15496_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15497_3_lut (.I0(\data_out_frame[18] [3]), .I1(displacement[19]), 
            .I2(n23935), .I3(GND_net), .O(n28560));   // verilog/coms.v(127[12] 300[6])
    defparam i15497_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15498_3_lut (.I0(\data_out_frame[18] [2]), .I1(displacement[18]), 
            .I2(n23935), .I3(GND_net), .O(n28561));   // verilog/coms.v(127[12] 300[6])
    defparam i15498_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15500_3_lut (.I0(\data_out_frame[18] [0]), .I1(displacement[16]), 
            .I2(n23935), .I3(GND_net), .O(n28563));   // verilog/coms.v(127[12] 300[6])
    defparam i15500_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15204_3_lut (.I0(PWMLimit[11]), .I1(\data_in_frame[9] [3]), 
            .I2(n27771), .I3(GND_net), .O(n28267));   // verilog/coms.v(127[12] 300[6])
    defparam i15204_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15501_3_lut (.I0(\data_out_frame[17] [7]), .I1(duty[7]), .I2(n23935), 
            .I3(GND_net), .O(n28564));   // verilog/coms.v(127[12] 300[6])
    defparam i15501_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15205_3_lut (.I0(PWMLimit[10]), .I1(\data_in_frame[9] [2]), 
            .I2(n27771), .I3(GND_net), .O(n28268));   // verilog/coms.v(127[12] 300[6])
    defparam i15205_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15206_3_lut (.I0(PWMLimit[9]), .I1(\data_in_frame[9] [1]), 
            .I2(n27771), .I3(GND_net), .O(n28269));   // verilog/coms.v(127[12] 300[6])
    defparam i15206_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15207_3_lut (.I0(PWMLimit[8]), .I1(\data_in_frame[9] [0]), 
            .I2(n27771), .I3(GND_net), .O(n28270));   // verilog/coms.v(127[12] 300[6])
    defparam i15207_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15502_3_lut (.I0(\data_out_frame[17] [6]), .I1(duty[6]), .I2(n23935), 
            .I3(GND_net), .O(n28565));   // verilog/coms.v(127[12] 300[6])
    defparam i15502_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15503_3_lut (.I0(\data_out_frame[17] [5]), .I1(duty[5]), .I2(n23935), 
            .I3(GND_net), .O(n28566));   // verilog/coms.v(127[12] 300[6])
    defparam i15503_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15504_3_lut (.I0(\data_out_frame[17] [4]), .I1(duty[4]), .I2(n23935), 
            .I3(GND_net), .O(n28567));   // verilog/coms.v(127[12] 300[6])
    defparam i15504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15505_3_lut (.I0(\data_out_frame[17] [3]), .I1(duty[3]), .I2(n23935), 
            .I3(GND_net), .O(n28568));   // verilog/coms.v(127[12] 300[6])
    defparam i15505_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15506_3_lut (.I0(\data_out_frame[17] [2]), .I1(duty[2]), .I2(n23935), 
            .I3(GND_net), .O(n28569));   // verilog/coms.v(127[12] 300[6])
    defparam i15506_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15507_3_lut (.I0(\data_out_frame[17] [1]), .I1(duty[1]), .I2(n23935), 
            .I3(GND_net), .O(n28570));   // verilog/coms.v(127[12] 300[6])
    defparam i15507_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i570_3_lut (.I0(n831), .I1(n898), 
            .I2(n861), .I3(GND_net), .O(n930));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i637_3_lut (.I0(n930), .I1(n997), 
            .I2(n960), .I3(GND_net), .O(n1029));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15508_3_lut (.I0(\data_out_frame[17] [0]), .I1(duty[0]), .I2(n23935), 
            .I3(GND_net), .O(n28571));   // verilog/coms.v(127[12] 300[6])
    defparam i15508_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29926_3_lut (.I0(n5_adj_4950), .I1(n6537), .I2(n44804), .I3(GND_net), 
            .O(n44809));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i29926_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17189_3_lut (.I0(\data_out_frame[16] [7]), .I1(duty[15]), .I2(n23935), 
            .I3(GND_net), .O(n28572));
    defparam i17189_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15510_3_lut (.I0(\data_out_frame[16] [6]), .I1(duty[14]), .I2(n23935), 
            .I3(GND_net), .O(n28573));   // verilog/coms.v(127[12] 300[6])
    defparam i15510_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15511_3_lut (.I0(\data_out_frame[16] [5]), .I1(duty[13]), .I2(n23935), 
            .I3(GND_net), .O(n28574));   // verilog/coms.v(127[12] 300[6])
    defparam i15511_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29927_3_lut (.I0(encoder0_position[28]), .I1(n44809), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n831));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i29927_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15512_3_lut (.I0(\data_out_frame[16] [4]), .I1(duty[12]), .I2(n23935), 
            .I3(GND_net), .O(n28575));   // verilog/coms.v(127[12] 300[6])
    defparam i15512_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15513_3_lut (.I0(\data_out_frame[16] [3]), .I1(duty[11]), .I2(n23935), 
            .I3(GND_net), .O(n28576));   // verilog/coms.v(127[12] 300[6])
    defparam i15513_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_833_4_lut (.I0(GND_net), .I1(n1232), 
            .I2(GND_net), .I3(n39666), .O(n1299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15514_3_lut (.I0(\data_out_frame[16] [2]), .I1(duty[10]), .I2(n23935), 
            .I3(GND_net), .O(n28577));   // verilog/coms.v(127[12] 300[6])
    defparam i15514_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15515_3_lut (.I0(\data_out_frame[16] [1]), .I1(duty[9]), .I2(n23935), 
            .I3(GND_net), .O(n28578));   // verilog/coms.v(127[12] 300[6])
    defparam i15515_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15516_3_lut (.I0(\data_out_frame[16] [0]), .I1(duty[8]), .I2(n23935), 
            .I3(GND_net), .O(n28579));   // verilog/coms.v(127[12] 300[6])
    defparam i15516_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15517_3_lut (.I0(\data_out_frame[15] [7]), .I1(duty[23]), .I2(n23935), 
            .I3(GND_net), .O(n28580));   // verilog/coms.v(127[12] 300[6])
    defparam i15517_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15518_3_lut (.I0(\data_out_frame[15] [6]), .I1(duty[22]), .I2(n23935), 
            .I3(GND_net), .O(n28581));   // verilog/coms.v(127[12] 300[6])
    defparam i15518_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15519_3_lut (.I0(\data_out_frame[15] [5]), .I1(duty[21]), .I2(n23935), 
            .I3(GND_net), .O(n28582));   // verilog/coms.v(127[12] 300[6])
    defparam i15519_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15520_3_lut (.I0(\data_out_frame[15] [4]), .I1(duty[20]), .I2(n23935), 
            .I3(GND_net), .O(n28583));   // verilog/coms.v(127[12] 300[6])
    defparam i15520_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15521_3_lut (.I0(\data_out_frame[15] [3]), .I1(duty[19]), .I2(n23935), 
            .I3(GND_net), .O(n28584));   // verilog/coms.v(127[12] 300[6])
    defparam i15521_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15522_3_lut (.I0(\data_out_frame[15] [2]), .I1(duty[18]), .I2(n23935), 
            .I3(GND_net), .O(n28585));   // verilog/coms.v(127[12] 300[6])
    defparam i15522_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1040_3_lut (.I0(n1525), .I1(n1592), 
            .I2(n1554), .I3(GND_net), .O(n1624));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1040_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15523_3_lut (.I0(\data_out_frame[15] [1]), .I1(duty[17]), .I2(n23935), 
            .I3(GND_net), .O(n28586));   // verilog/coms.v(127[12] 300[6])
    defparam i15523_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15524_3_lut (.I0(\data_out_frame[15] [0]), .I1(duty[16]), .I2(n23935), 
            .I3(GND_net), .O(n28587));   // verilog/coms.v(127[12] 300[6])
    defparam i15524_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15525_3_lut (.I0(\data_out_frame[14] [7]), .I1(setpoint[7]), 
            .I2(n23935), .I3(GND_net), .O(n28588));   // verilog/coms.v(127[12] 300[6])
    defparam i15525_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15526_3_lut (.I0(\data_out_frame[14] [6]), .I1(setpoint[6]), 
            .I2(n23935), .I3(GND_net), .O(n28589));   // verilog/coms.v(127[12] 300[6])
    defparam i15526_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15527_3_lut (.I0(\data_out_frame[14] [5]), .I1(setpoint[5]), 
            .I2(n23935), .I3(GND_net), .O(n28590));   // verilog/coms.v(127[12] 300[6])
    defparam i15527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15528_3_lut (.I0(\data_out_frame[14] [4]), .I1(setpoint[4]), 
            .I2(n23935), .I3(GND_net), .O(n28591));   // verilog/coms.v(127[12] 300[6])
    defparam i15528_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15529_3_lut (.I0(\data_out_frame[14] [3]), .I1(setpoint[3]), 
            .I2(n23935), .I3(GND_net), .O(n28592));   // verilog/coms.v(127[12] 300[6])
    defparam i15529_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15530_3_lut (.I0(\data_out_frame[14] [2]), .I1(setpoint[2]), 
            .I2(n23935), .I3(GND_net), .O(n28593));   // verilog/coms.v(127[12] 300[6])
    defparam i15530_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15531_3_lut (.I0(\data_out_frame[14] [1]), .I1(setpoint[1]), 
            .I2(n23935), .I3(GND_net), .O(n28594));   // verilog/coms.v(127[12] 300[6])
    defparam i15531_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n5722), 
            .D(n680), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 i15532_3_lut (.I0(\data_out_frame[14] [0]), .I1(setpoint[0]), 
            .I2(n23935), .I3(GND_net), .O(n28595));   // verilog/coms.v(127[12] 300[6])
    defparam i15532_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i29 (.Q(delay_counter[29]), .C(CLK_c), .E(n5722), 
            .D(n661), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 i15533_3_lut (.I0(\data_out_frame[13] [7]), .I1(setpoint[15]), 
            .I2(n23935), .I3(GND_net), .O(n28596));   // verilog/coms.v(127[12] 300[6])
    defparam i15533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15534_3_lut (.I0(\data_out_frame[13] [6]), .I1(setpoint[14]), 
            .I2(n23935), .I3(GND_net), .O(n28597));   // verilog/coms.v(127[12] 300[6])
    defparam i15534_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15535_3_lut (.I0(\data_out_frame[13] [5]), .I1(setpoint[13]), 
            .I2(n23935), .I3(GND_net), .O(n28598));   // verilog/coms.v(127[12] 300[6])
    defparam i15535_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15536_3_lut (.I0(\data_out_frame[13] [4]), .I1(setpoint[12]), 
            .I2(n23935), .I3(GND_net), .O(n28599));   // verilog/coms.v(127[12] 300[6])
    defparam i15536_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15537_3_lut (.I0(\data_out_frame[13] [3]), .I1(setpoint[11]), 
            .I2(n23935), .I3(GND_net), .O(n28600));   // verilog/coms.v(127[12] 300[6])
    defparam i15537_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15538_3_lut (.I0(\data_out_frame[13] [2]), .I1(setpoint[10]), 
            .I2(n23935), .I3(GND_net), .O(n28601));   // verilog/coms.v(127[12] 300[6])
    defparam i15538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15539_3_lut (.I0(\data_out_frame[13] [1]), .I1(setpoint[9]), 
            .I2(n23935), .I3(GND_net), .O(n28602));   // verilog/coms.v(127[12] 300[6])
    defparam i15539_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n5722), 
            .D(n681), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 i15540_3_lut (.I0(\data_out_frame[13] [0]), .I1(setpoint[8]), 
            .I2(n23935), .I3(GND_net), .O(n28603));   // verilog/coms.v(127[12] 300[6])
    defparam i15540_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15541_3_lut (.I0(\data_out_frame[12] [7]), .I1(setpoint[23]), 
            .I2(n23935), .I3(GND_net), .O(n28604));   // verilog/coms.v(127[12] 300[6])
    defparam i15541_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_833_4 (.CI(n39666), .I0(n1232), 
            .I1(GND_net), .CO(n39667));
    SB_LUT4 i15542_3_lut (.I0(\data_out_frame[12] [6]), .I1(setpoint[22]), 
            .I2(n23935), .I3(GND_net), .O(n28605));   // verilog/coms.v(127[12] 300[6])
    defparam i15542_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_3_lut (.I0(n5_adj_4912), .I1(n3_adj_4952), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n47311));
    defparam i1_3_lut.LUT_INIT = 16'h8080;
    SB_DFF pwm_setpoint_i0 (.Q(pwm_setpoint[0]), .C(CLK_c), .D(pwm_setpoint_22__N_11[0]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 encoder0_position_31__I_0_i500_4_lut (.I0(n2_adj_4953), .I1(n6534), 
            .I2(n47311), .I3(encoder0_position[31]), .O(n828));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i500_4_lut.LUT_INIT = 16'h8a80;
    SB_LUT4 i15543_3_lut (.I0(\data_out_frame[12] [5]), .I1(setpoint[21]), 
            .I2(n23935), .I3(GND_net), .O(n28606));   // verilog/coms.v(127[12] 300[6])
    defparam i15543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15544_3_lut (.I0(\data_out_frame[12] [4]), .I1(setpoint[20]), 
            .I2(n23935), .I3(GND_net), .O(n28607));   // verilog/coms.v(127[12] 300[6])
    defparam i15544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i28_3_lut (.I0(encoder0_position[27]), 
            .I1(n6_adj_4949), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n625));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i28_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i29_3_lut (.I0(encoder0_position[28]), 
            .I1(n5_adj_4950), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n516));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i29_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1302_3_lut (.I0(GND_net), .I1(n1933), 
            .I2(VCC_net), .I3(n39766), .O(n2000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_833_3_lut (.I0(GND_net), .I1(n1233), 
            .I2(VCC_net), .I3(n39665), .O(n1300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36021_1_lut (.I0(n1752), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50974));
    defparam i36021_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i1_1_lut (.I0(duty[0]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n25));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i30_3_lut (.I0(encoder0_position[29]), 
            .I1(n4_adj_4951), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n623));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_833_3 (.CI(n39665), .I0(n1233), 
            .I1(VCC_net), .CO(n39666));
    SB_LUT4 unary_minus_4_inv_0_i2_1_lut (.I0(duty[1]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n24));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i31_3_lut (.I0(encoder0_position[30]), 
            .I1(n3_adj_4952), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n622));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i31_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4091_2_lut (.I0(n2_adj_4953), .I1(encoder0_position[31]), .I2(GND_net), 
            .I3(GND_net), .O(n621));
    defparam i4091_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15545_3_lut (.I0(\data_out_frame[12] [3]), .I1(setpoint[19]), 
            .I2(n23935), .I3(GND_net), .O(n28608));   // verilog/coms.v(127[12] 300[6])
    defparam i15545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_4_inv_0_i3_1_lut (.I0(duty[2]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n23));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15140_4_lut (.I0(r_Rx_Data), .I1(rx_data[2]), .I2(n4_adj_4916), 
            .I3(n26629), .O(n28203));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15140_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_4_inv_0_i4_1_lut (.I0(duty[3]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n22));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i5_1_lut (.I0(duty[4]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n21));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1302_3 (.CI(n39766), .I0(n1933), 
            .I1(VCC_net), .CO(n39767));
    SB_LUT4 encoder0_position_31__I_0_add_833_2_lut (.I0(GND_net), .I1(n937), 
            .I2(GND_net), .I3(VCC_net), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15141_4_lut (.I0(state_7__N_4003[3]), .I1(data[4]), .I2(n4_adj_4915), 
            .I3(n26645), .O(n28204));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15141_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_31__I_0_add_833_2 (.CI(VCC_net), .I0(n937), 
            .I1(GND_net), .CO(n39665));
    SB_LUT4 encoder0_position_31__I_0_add_1302_2_lut (.I0(GND_net), .I1(n944), 
            .I2(GND_net), .I3(VCC_net), .O(n2001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_2 (.CI(VCC_net), .I0(n944), 
            .I1(GND_net), .CO(n39766));
    SB_LUT4 encoder0_position_31__I_0_i1043_3_lut (.I0(n1528), .I1(n1595), 
            .I2(n1554), .I3(GND_net), .O(n1627));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1235_18_lut (.I0(n50998), .I1(n1818), 
            .I2(VCC_net), .I3(n39765), .O(n1917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_i1041_3_lut (.I0(n1526), .I1(n1593), 
            .I2(n1554), .I3(GND_net), .O(n1625));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1041_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i971_3_lut (.I0(n1424), .I1(n1491), 
            .I2(n1455), .I3(GND_net), .O(n1523));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i971_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36437_1_lut (.I0(n2544), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51390));
    defparam i36437_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i6_1_lut (.I0(duty[5]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n20));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35787_1_lut (.I0(n2643), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50740));
    defparam i35787_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i7_1_lut (.I0(duty[6]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n19));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR delay_counter_i0_i28 (.Q(delay_counter[28]), .C(CLK_c), .E(n5722), 
            .D(n662), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 i15142_4_lut (.I0(state_7__N_4003[3]), .I1(data[3]), .I2(n4_adj_4914), 
            .I3(n26650), .O(n28205));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15142_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15546_3_lut (.I0(\data_out_frame[12] [2]), .I1(setpoint[18]), 
            .I2(n23935), .I3(GND_net), .O(n28609));   // verilog/coms.v(127[12] 300[6])
    defparam i15546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15547_3_lut (.I0(\data_out_frame[12] [1]), .I1(setpoint[17]), 
            .I2(n23935), .I3(GND_net), .O(n28610));   // verilog/coms.v(127[12] 300[6])
    defparam i15547_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i27 (.Q(delay_counter[27]), .C(CLK_c), .E(n5722), 
            .D(n663), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 i15548_3_lut (.I0(\data_out_frame[12] [0]), .I1(setpoint[16]), 
            .I2(n23935), .I3(GND_net), .O(n28611));   // verilog/coms.v(127[12] 300[6])
    defparam i15548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15549_3_lut (.I0(\data_out_frame[11] [7]), .I1(encoder1_position_scaled[7]), 
            .I2(n23935), .I3(GND_net), .O(n28612));   // verilog/coms.v(127[12] 300[6])
    defparam i15549_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n5722), 
            .D(n687), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 i15550_3_lut (.I0(\data_out_frame[11] [6]), .I1(encoder1_position_scaled[6]), 
            .I2(n23935), .I3(GND_net), .O(n28613));   // verilog/coms.v(127[12] 300[6])
    defparam i15550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15551_3_lut (.I0(\data_out_frame[11] [5]), .I1(encoder1_position_scaled[5]), 
            .I2(n23935), .I3(GND_net), .O(n28614));   // verilog/coms.v(127[12] 300[6])
    defparam i15551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1235_17_lut (.I0(GND_net), .I1(n1819), 
            .I2(VCC_net), .I3(n39764), .O(n1886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15552_3_lut (.I0(\data_out_frame[11] [4]), .I1(encoder1_position_scaled[4]), 
            .I2(n23935), .I3(GND_net), .O(n28615));   // verilog/coms.v(127[12] 300[6])
    defparam i15552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15553_3_lut (.I0(\data_out_frame[11] [3]), .I1(encoder1_position_scaled[3]), 
            .I2(n23935), .I3(GND_net), .O(n28616));   // verilog/coms.v(127[12] 300[6])
    defparam i15553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15554_3_lut (.I0(\data_out_frame[11] [2]), .I1(encoder1_position_scaled[2]), 
            .I2(n23935), .I3(GND_net), .O(n28617));   // verilog/coms.v(127[12] 300[6])
    defparam i15554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15555_3_lut (.I0(\data_out_frame[11] [1]), .I1(encoder1_position_scaled[1]), 
            .I2(n23935), .I3(GND_net), .O(n28618));   // verilog/coms.v(127[12] 300[6])
    defparam i15555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_33_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n2_adj_4991), .I3(n40534), .O(n2_adj_4953)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_32_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n3_adj_4992), .I3(n40533), .O(n3_adj_4952)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15556_3_lut (.I0(\data_out_frame[11] [0]), .I1(encoder1_position_scaled[0]), 
            .I2(n23935), .I3(GND_net), .O(n28619));   // verilog/coms.v(127[12] 300[6])
    defparam i15556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15557_3_lut (.I0(\data_out_frame[10] [7]), .I1(encoder1_position_scaled[15]), 
            .I2(n23935), .I3(GND_net), .O(n28620));   // verilog/coms.v(127[12] 300[6])
    defparam i15557_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_32 (.CI(n40533), 
            .I0(GND_net), .I1(n3_adj_4992), .CO(n40534));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_31_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n4_adj_4993), .I3(n40532), .O(n4_adj_4951)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_31 (.CI(n40532), 
            .I0(GND_net), .I1(n4_adj_4993), .CO(n40533));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_30_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n5_adj_4994), .I3(n40531), .O(n5_adj_4950)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15558_3_lut (.I0(\data_out_frame[10] [6]), .I1(encoder1_position_scaled[14]), 
            .I2(n23935), .I3(GND_net), .O(n28621));   // verilog/coms.v(127[12] 300[6])
    defparam i15558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15559_3_lut (.I0(\data_out_frame[10] [5]), .I1(encoder1_position_scaled[13]), 
            .I2(n23935), .I3(GND_net), .O(n28622));   // verilog/coms.v(127[12] 300[6])
    defparam i15559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15560_3_lut (.I0(\data_out_frame[10] [4]), .I1(encoder1_position_scaled[12]), 
            .I2(n23935), .I3(GND_net), .O(n28623));   // verilog/coms.v(127[12] 300[6])
    defparam i15560_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15561_3_lut (.I0(\data_out_frame[10] [3]), .I1(encoder1_position_scaled[11]), 
            .I2(n23935), .I3(GND_net), .O(n28624));   // verilog/coms.v(127[12] 300[6])
    defparam i15561_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1235_17 (.CI(n39764), .I0(n1819), 
            .I1(VCC_net), .CO(n39765));
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_30 (.CI(n40531), 
            .I0(GND_net), .I1(n5_adj_4994), .CO(n40532));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_29_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n6_adj_4995), .I3(n40530), .O(n6_adj_4949)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_29 (.CI(n40530), 
            .I0(GND_net), .I1(n6_adj_4995), .CO(n40531));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_28_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n7_adj_4996), .I3(n40529), .O(n7_adj_4948)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_28 (.CI(n40529), 
            .I0(GND_net), .I1(n7_adj_4996), .CO(n40530));
    SB_LUT4 i15562_3_lut (.I0(\data_out_frame[10] [2]), .I1(encoder1_position_scaled[10]), 
            .I2(n23935), .I3(GND_net), .O(n28625));   // verilog/coms.v(127[12] 300[6])
    defparam i15562_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_27_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n8_adj_4997), .I3(n40528), .O(n8_adj_4934)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_27_lut.LUT_INIT = 16'hC33C;
    SB_IO INLC_pad (.PACKAGE_PIN(INLC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(VCC_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLC_pad.PIN_TYPE = 6'b011001;
    defparam INLC_pad.PULLUP = 1'b0;
    defparam INLC_pad.NEG_TRIGGER = 1'b0;
    defparam INLC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_27 (.CI(n40528), 
            .I0(GND_net), .I1(n8_adj_4997), .CO(n40529));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_26_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n9_adj_4998), .I3(n40527), .O(n9_adj_4933)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_26 (.CI(n40527), 
            .I0(GND_net), .I1(n9_adj_4998), .CO(n40528));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_25_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n10_adj_4999), .I3(n40526), .O(n10_adj_4932)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_25 (.CI(n40526), 
            .I0(GND_net), .I1(n10_adj_4999), .CO(n40527));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_24_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n11_adj_5000), .I3(n40525), .O(n11_adj_4931)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n5722), 
            .D(n688), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_24 (.CI(n40525), 
            .I0(GND_net), .I1(n11_adj_5000), .CO(n40526));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_23_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n12_adj_5001), .I3(n40524), .O(n12_adj_4930)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15563_3_lut (.I0(\data_out_frame[10] [1]), .I1(encoder1_position_scaled[9]), 
            .I2(n23935), .I3(GND_net), .O(n28626));   // verilog/coms.v(127[12] 300[6])
    defparam i15563_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15564_3_lut (.I0(\data_out_frame[10] [0]), .I1(encoder1_position_scaled[8]), 
            .I2(n23935), .I3(GND_net), .O(n28627));   // verilog/coms.v(127[12] 300[6])
    defparam i15564_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_23 (.CI(n40524), 
            .I0(GND_net), .I1(n12_adj_5001), .CO(n40525));
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n5722), 
            .D(n689), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_22_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n13_adj_5002), .I3(n40523), .O(n13_adj_4929)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15565_3_lut (.I0(\data_out_frame[9] [7]), .I1(encoder1_position_scaled[23]), 
            .I2(n23935), .I3(GND_net), .O(n28628));   // verilog/coms.v(127[12] 300[6])
    defparam i15565_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15566_3_lut (.I0(\data_out_frame[9] [6]), .I1(encoder1_position_scaled[22]), 
            .I2(n23935), .I3(GND_net), .O(n28629));   // verilog/coms.v(127[12] 300[6])
    defparam i15566_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15567_3_lut (.I0(\data_out_frame[9] [5]), .I1(encoder1_position_scaled[21]), 
            .I2(n23935), .I3(GND_net), .O(n28630));   // verilog/coms.v(127[12] 300[6])
    defparam i15567_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15568_3_lut (.I0(\data_out_frame[9] [4]), .I1(encoder1_position_scaled[20]), 
            .I2(n23935), .I3(GND_net), .O(n28631));   // verilog/coms.v(127[12] 300[6])
    defparam i15568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15569_3_lut (.I0(\data_out_frame[9] [3]), .I1(encoder1_position_scaled[19]), 
            .I2(n23935), .I3(GND_net), .O(n28632));   // verilog/coms.v(127[12] 300[6])
    defparam i15569_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_22 (.CI(n40523), 
            .I0(GND_net), .I1(n13_adj_5002), .CO(n40524));
    SB_LUT4 i15570_3_lut (.I0(\data_out_frame[9] [2]), .I1(encoder1_position_scaled[18]), 
            .I2(n23935), .I3(GND_net), .O(n28633));   // verilog/coms.v(127[12] 300[6])
    defparam i15570_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_21_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n14_adj_5003), .I3(n40522), .O(n14_adj_4928)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_21 (.CI(n40522), 
            .I0(GND_net), .I1(n14_adj_5003), .CO(n40523));
    SB_LUT4 i15571_3_lut (.I0(\data_out_frame[9] [1]), .I1(encoder1_position_scaled[17]), 
            .I2(n23935), .I3(GND_net), .O(n28634));   // verilog/coms.v(127[12] 300[6])
    defparam i15571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15572_3_lut (.I0(\data_out_frame[9] [0]), .I1(encoder1_position_scaled[16]), 
            .I2(n23935), .I3(GND_net), .O(n28635));   // verilog/coms.v(127[12] 300[6])
    defparam i15572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_20_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n15_adj_5004), .I3(n40521), .O(n15_adj_4927)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_20 (.CI(n40521), 
            .I0(GND_net), .I1(n15_adj_5004), .CO(n40522));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_19_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n16_adj_5005), .I3(n40520), .O(n16_adj_4926)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15573_3_lut (.I0(\data_out_frame[8] [7]), .I1(encoder0_position_scaled[7]), 
            .I2(n23935), .I3(GND_net), .O(n28636));   // verilog/coms.v(127[12] 300[6])
    defparam i15573_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_19 (.CI(n40520), 
            .I0(GND_net), .I1(n16_adj_5005), .CO(n40521));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_18_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n17_adj_5006), .I3(n40519), .O(n17_adj_4925)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15574_3_lut (.I0(\data_out_frame[8] [6]), .I1(encoder0_position_scaled[6]), 
            .I2(n23935), .I3(GND_net), .O(n28637));   // verilog/coms.v(127[12] 300[6])
    defparam i15574_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15575_3_lut (.I0(\data_out_frame[8] [5]), .I1(encoder0_position_scaled[5]), 
            .I2(n23935), .I3(GND_net), .O(n28638));   // verilog/coms.v(127[12] 300[6])
    defparam i15575_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_18 (.CI(n40519), 
            .I0(GND_net), .I1(n17_adj_5006), .CO(n40520));
    SB_LUT4 i15576_3_lut (.I0(\data_out_frame[8] [4]), .I1(encoder0_position_scaled[4]), 
            .I2(n23935), .I3(GND_net), .O(n28639));   // verilog/coms.v(127[12] 300[6])
    defparam i15576_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15577_3_lut (.I0(\data_out_frame[8] [3]), .I1(encoder0_position_scaled[3]), 
            .I2(n23935), .I3(GND_net), .O(n28640));   // verilog/coms.v(127[12] 300[6])
    defparam i15577_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15578_3_lut (.I0(\data_out_frame[8] [2]), .I1(encoder0_position_scaled[2]), 
            .I2(n23935), .I3(GND_net), .O(n28641));   // verilog/coms.v(127[12] 300[6])
    defparam i15578_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15579_3_lut (.I0(\data_out_frame[8] [1]), .I1(encoder0_position_scaled[1]), 
            .I2(n23935), .I3(GND_net), .O(n28642));   // verilog/coms.v(127[12] 300[6])
    defparam i15579_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_17_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n18_adj_5007), .I3(n40518), .O(n18_adj_4924)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_17 (.CI(n40518), 
            .I0(GND_net), .I1(n18_adj_5007), .CO(n40519));
    SB_LUT4 encoder0_position_31__I_0_add_1235_16_lut (.I0(GND_net), .I1(n1820), 
            .I2(VCC_net), .I3(n39763), .O(n1887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_16_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n19_adj_5008), .I3(n40517), .O(n19_adj_4923)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_16 (.CI(n40517), 
            .I0(GND_net), .I1(n19_adj_5008), .CO(n40518));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_15_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n20_adj_5009), .I3(n40516), .O(n20_adj_4922)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15580_3_lut (.I0(\data_out_frame[8] [0]), .I1(encoder0_position_scaled[0]), 
            .I2(n23935), .I3(GND_net), .O(n28643));   // verilog/coms.v(127[12] 300[6])
    defparam i15580_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_15 (.CI(n40516), 
            .I0(GND_net), .I1(n20_adj_5009), .CO(n40517));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_14_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n21_adj_5010), .I3(n40515), .O(n21_adj_4921)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_14 (.CI(n40515), 
            .I0(GND_net), .I1(n21_adj_5010), .CO(n40516));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_13_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n22_adj_5011), .I3(n40514), .O(n22_adj_4920)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_13 (.CI(n40514), 
            .I0(GND_net), .I1(n22_adj_5011), .CO(n40515));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_12_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n23_adj_5012), .I3(n40513), .O(n23_adj_4919)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_12 (.CI(n40513), 
            .I0(GND_net), .I1(n23_adj_5012), .CO(n40514));
    SB_DFFESR delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n5722), 
            .D(n682), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_11_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n24_adj_5013), .I3(n40512), .O(n24_adj_4918)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_11 (.CI(n40512), 
            .I0(GND_net), .I1(n24_adj_5013), .CO(n40513));
    SB_LUT4 i15581_3_lut (.I0(\data_out_frame[7] [7]), .I1(encoder0_position_scaled[15]), 
            .I2(n23935), .I3(GND_net), .O(n28644));   // verilog/coms.v(127[12] 300[6])
    defparam i15581_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_10_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n25_adj_5014), .I3(n40511), .O(n25_adj_4917)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_10 (.CI(n40511), 
            .I0(GND_net), .I1(n25_adj_5014), .CO(n40512));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_9_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n26_adj_5015), .I3(n40510), .O(n26)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_9 (.CI(n40510), 
            .I0(GND_net), .I1(n26_adj_5015), .CO(n40511));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_8_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n27_adj_5016), .I3(n40509), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_16 (.CI(n39763), .I0(n1820), 
            .I1(VCC_net), .CO(n39764));
    SB_LUT4 encoder0_position_31__I_0_add_1235_15_lut (.I0(GND_net), .I1(n1821), 
            .I2(VCC_net), .I3(n39762), .O(n1888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15582_3_lut (.I0(\data_out_frame[7] [6]), .I1(encoder0_position_scaled[14]), 
            .I2(n23935), .I3(GND_net), .O(n28645));   // verilog/coms.v(127[12] 300[6])
    defparam i15582_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15583_3_lut (.I0(\data_out_frame[7] [5]), .I1(encoder0_position_scaled[13]), 
            .I2(n23935), .I3(GND_net), .O(n28646));   // verilog/coms.v(127[12] 300[6])
    defparam i15583_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15584_3_lut (.I0(\data_out_frame[7] [4]), .I1(encoder0_position_scaled[12]), 
            .I2(n23935), .I3(GND_net), .O(n28647));   // verilog/coms.v(127[12] 300[6])
    defparam i15584_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15585_3_lut (.I0(\data_out_frame[7] [3]), .I1(encoder0_position_scaled[11]), 
            .I2(n23935), .I3(GND_net), .O(n28648));   // verilog/coms.v(127[12] 300[6])
    defparam i15585_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15586_3_lut (.I0(\data_out_frame[7] [2]), .I1(encoder0_position_scaled[10]), 
            .I2(n23935), .I3(GND_net), .O(n28649));   // verilog/coms.v(127[12] 300[6])
    defparam i15586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15587_3_lut (.I0(\data_out_frame[7] [1]), .I1(encoder0_position_scaled[9]), 
            .I2(n23935), .I3(GND_net), .O(n28650));   // verilog/coms.v(127[12] 300[6])
    defparam i15587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15588_3_lut (.I0(\data_out_frame[7] [0]), .I1(encoder0_position_scaled[8]), 
            .I2(n23935), .I3(GND_net), .O(n28651));   // verilog/coms.v(127[12] 300[6])
    defparam i15588_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15589_3_lut (.I0(\data_out_frame[6] [7]), .I1(encoder0_position_scaled[23]), 
            .I2(n23935), .I3(GND_net), .O(n28652));   // verilog/coms.v(127[12] 300[6])
    defparam i15589_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15590_3_lut (.I0(\data_out_frame[6] [6]), .I1(encoder0_position_scaled[22]), 
            .I2(n23935), .I3(GND_net), .O(n28653));   // verilog/coms.v(127[12] 300[6])
    defparam i15590_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15591_3_lut (.I0(\data_out_frame[6] [5]), .I1(encoder0_position_scaled[21]), 
            .I2(n23935), .I3(GND_net), .O(n28654));   // verilog/coms.v(127[12] 300[6])
    defparam i15591_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15592_3_lut (.I0(\data_out_frame[6] [4]), .I1(encoder0_position_scaled[20]), 
            .I2(n23935), .I3(GND_net), .O(n28655));   // verilog/coms.v(127[12] 300[6])
    defparam i15592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15593_3_lut (.I0(\data_out_frame[6] [3]), .I1(encoder0_position_scaled[19]), 
            .I2(n23935), .I3(GND_net), .O(n28656));   // verilog/coms.v(127[12] 300[6])
    defparam i15593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15594_3_lut (.I0(\data_out_frame[6] [2]), .I1(encoder0_position_scaled[18]), 
            .I2(n23935), .I3(GND_net), .O(n28657));   // verilog/coms.v(127[12] 300[6])
    defparam i15594_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15595_3_lut (.I0(\data_out_frame[6] [1]), .I1(encoder0_position_scaled[17]), 
            .I2(n23935), .I3(GND_net), .O(n28658));   // verilog/coms.v(127[12] 300[6])
    defparam i15595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15596_3_lut (.I0(\data_out_frame[6] [0]), .I1(encoder0_position_scaled[16]), 
            .I2(n23935), .I3(GND_net), .O(n28659));   // verilog/coms.v(127[12] 300[6])
    defparam i15596_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15597_3_lut (.I0(\data_out_frame[5] [7]), .I1(control_mode[7]), 
            .I2(n23935), .I3(GND_net), .O(n28660));   // verilog/coms.v(127[12] 300[6])
    defparam i15597_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15598_3_lut (.I0(\data_out_frame[5] [6]), .I1(control_mode[6]), 
            .I2(n23935), .I3(GND_net), .O(n28661));   // verilog/coms.v(127[12] 300[6])
    defparam i15598_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15599_3_lut (.I0(\data_out_frame[5] [5]), .I1(control_mode[5]), 
            .I2(n23935), .I3(GND_net), .O(n28662));   // verilog/coms.v(127[12] 300[6])
    defparam i15599_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15600_3_lut (.I0(\data_out_frame[5] [4]), .I1(control_mode[4]), 
            .I2(n23935), .I3(GND_net), .O(n28663));   // verilog/coms.v(127[12] 300[6])
    defparam i15600_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15601_3_lut (.I0(\data_out_frame[5] [3]), .I1(control_mode[3]), 
            .I2(n23935), .I3(GND_net), .O(n28664));   // verilog/coms.v(127[12] 300[6])
    defparam i15601_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15602_3_lut (.I0(\data_out_frame[5] [2]), .I1(control_mode[2]), 
            .I2(n23935), .I3(GND_net), .O(n28665));   // verilog/coms.v(127[12] 300[6])
    defparam i15602_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15603_3_lut (.I0(\data_out_frame[5] [1]), .I1(control_mode[1]), 
            .I2(n23935), .I3(GND_net), .O(n28666));   // verilog/coms.v(127[12] 300[6])
    defparam i15603_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15604_3_lut (.I0(\data_out_frame[5] [0]), .I1(control_mode[0]), 
            .I2(n23935), .I3(GND_net), .O(n28667));   // verilog/coms.v(127[12] 300[6])
    defparam i15604_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15605_3_lut (.I0(\data_out_frame[4] [7]), .I1(ID[7]), .I2(n23935), 
            .I3(GND_net), .O(n28668));   // verilog/coms.v(127[12] 300[6])
    defparam i15605_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i970_3_lut (.I0(n1423), .I1(n1490), 
            .I2(n1455), .I3(GND_net), .O(n1522));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i970_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15606_3_lut (.I0(\data_out_frame[4] [6]), .I1(ID[6]), .I2(n23935), 
            .I3(GND_net), .O(n28669));   // verilog/coms.v(127[12] 300[6])
    defparam i15606_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15607_3_lut (.I0(\data_out_frame[4] [5]), .I1(ID[5]), .I2(n23935), 
            .I3(GND_net), .O(n28670));   // verilog/coms.v(127[12] 300[6])
    defparam i15607_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15608_3_lut (.I0(\data_out_frame[4] [4]), .I1(ID[4]), .I2(n23935), 
            .I3(GND_net), .O(n28671));   // verilog/coms.v(127[12] 300[6])
    defparam i15608_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15609_3_lut (.I0(\data_out_frame[4] [3]), .I1(ID[3]), .I2(n23935), 
            .I3(GND_net), .O(n28672));   // verilog/coms.v(127[12] 300[6])
    defparam i15609_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15610_3_lut (.I0(\data_out_frame[4] [2]), .I1(ID[2]), .I2(n23935), 
            .I3(GND_net), .O(n28673));   // verilog/coms.v(127[12] 300[6])
    defparam i15610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15611_3_lut (.I0(\data_out_frame[4] [1]), .I1(ID[1]), .I2(n23935), 
            .I3(GND_net), .O(n28674));   // verilog/coms.v(127[12] 300[6])
    defparam i15611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15612_3_lut (.I0(\data_out_frame[4] [0]), .I1(ID[0]), .I2(n23935), 
            .I3(GND_net), .O(n28675));   // verilog/coms.v(127[12] 300[6])
    defparam i15612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15613_3_lut (.I0(Ki[15]), .I1(\data_in_frame[4] [7]), .I2(n27771), 
            .I3(GND_net), .O(n28676));   // verilog/coms.v(127[12] 300[6])
    defparam i15613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15614_3_lut (.I0(Ki[14]), .I1(\data_in_frame[4] [6]), .I2(n27771), 
            .I3(GND_net), .O(n28677));   // verilog/coms.v(127[12] 300[6])
    defparam i15614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15615_3_lut (.I0(Ki[13]), .I1(\data_in_frame[4] [5]), .I2(n27771), 
            .I3(GND_net), .O(n28678));   // verilog/coms.v(127[12] 300[6])
    defparam i15615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15616_3_lut (.I0(Ki[12]), .I1(\data_in_frame[4] [4]), .I2(n27771), 
            .I3(GND_net), .O(n28679));   // verilog/coms.v(127[12] 300[6])
    defparam i15616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15617_3_lut (.I0(Ki[11]), .I1(\data_in_frame[4] [3]), .I2(n27771), 
            .I3(GND_net), .O(n28680));   // verilog/coms.v(127[12] 300[6])
    defparam i15617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15618_3_lut (.I0(Ki[10]), .I1(\data_in_frame[4] [2]), .I2(n27771), 
            .I3(GND_net), .O(n28681));   // verilog/coms.v(127[12] 300[6])
    defparam i15618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15619_3_lut (.I0(Ki[9]), .I1(\data_in_frame[4] [1]), .I2(n27771), 
            .I3(GND_net), .O(n28682));   // verilog/coms.v(127[12] 300[6])
    defparam i15619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15620_3_lut (.I0(Ki[8]), .I1(\data_in_frame[4] [0]), .I2(n27771), 
            .I3(GND_net), .O(n28683));   // verilog/coms.v(127[12] 300[6])
    defparam i15620_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15621_3_lut (.I0(Ki[7]), .I1(\data_in_frame[5] [7]), .I2(n27771), 
            .I3(GND_net), .O(n28684));   // verilog/coms.v(127[12] 300[6])
    defparam i15621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15622_3_lut (.I0(Ki[6]), .I1(\data_in_frame[5] [6]), .I2(n27771), 
            .I3(GND_net), .O(n28685));   // verilog/coms.v(127[12] 300[6])
    defparam i15622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15623_3_lut (.I0(Ki[5]), .I1(\data_in_frame[5] [5]), .I2(n27771), 
            .I3(GND_net), .O(n28686));   // verilog/coms.v(127[12] 300[6])
    defparam i15623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15624_3_lut (.I0(Ki[4]), .I1(\data_in_frame[5] [4]), .I2(n27771), 
            .I3(GND_net), .O(n28687));   // verilog/coms.v(127[12] 300[6])
    defparam i15624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15625_3_lut (.I0(Ki[3]), .I1(\data_in_frame[5] [3]), .I2(n27771), 
            .I3(GND_net), .O(n28688));   // verilog/coms.v(127[12] 300[6])
    defparam i15625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15626_3_lut (.I0(Ki[2]), .I1(\data_in_frame[5] [2]), .I2(n27771), 
            .I3(GND_net), .O(n28689));   // verilog/coms.v(127[12] 300[6])
    defparam i15626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15627_3_lut (.I0(Ki[1]), .I1(\data_in_frame[5] [1]), .I2(n27771), 
            .I3(GND_net), .O(n28690));   // verilog/coms.v(127[12] 300[6])
    defparam i15627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15628_3_lut (.I0(Kp[15]), .I1(\data_in_frame[2] [7]), .I2(n27771), 
            .I3(GND_net), .O(n28691));   // verilog/coms.v(127[12] 300[6])
    defparam i15628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15629_3_lut (.I0(Kp[14]), .I1(\data_in_frame[2] [6]), .I2(n27771), 
            .I3(GND_net), .O(n28692));   // verilog/coms.v(127[12] 300[6])
    defparam i15629_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15630_3_lut (.I0(Kp[13]), .I1(\data_in_frame[2] [5]), .I2(n27771), 
            .I3(GND_net), .O(n28693));   // verilog/coms.v(127[12] 300[6])
    defparam i15630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15631_3_lut (.I0(Kp[12]), .I1(\data_in_frame[2] [4]), .I2(n27771), 
            .I3(GND_net), .O(n28694));   // verilog/coms.v(127[12] 300[6])
    defparam i15631_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15632_3_lut (.I0(Kp[11]), .I1(\data_in_frame[2] [3]), .I2(n27771), 
            .I3(GND_net), .O(n28695));   // verilog/coms.v(127[12] 300[6])
    defparam i15632_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15633_3_lut (.I0(Kp[10]), .I1(\data_in_frame[2] [2]), .I2(n27771), 
            .I3(GND_net), .O(n28696));   // verilog/coms.v(127[12] 300[6])
    defparam i15633_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15634_3_lut (.I0(Kp[9]), .I1(\data_in_frame[2] [1]), .I2(n27771), 
            .I3(GND_net), .O(n28697));   // verilog/coms.v(127[12] 300[6])
    defparam i15634_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15635_3_lut (.I0(Kp[8]), .I1(\data_in_frame[2] [0]), .I2(n27771), 
            .I3(GND_net), .O(n28698));   // verilog/coms.v(127[12] 300[6])
    defparam i15635_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15636_3_lut (.I0(Kp[7]), .I1(\data_in_frame[3] [7]), .I2(n27771), 
            .I3(GND_net), .O(n28699));   // verilog/coms.v(127[12] 300[6])
    defparam i15636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15637_3_lut (.I0(Kp[6]), .I1(\data_in_frame[3] [6]), .I2(n27771), 
            .I3(GND_net), .O(n28700));   // verilog/coms.v(127[12] 300[6])
    defparam i15637_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15638_3_lut (.I0(Kp[5]), .I1(\data_in_frame[3] [5]), .I2(n27771), 
            .I3(GND_net), .O(n28701));   // verilog/coms.v(127[12] 300[6])
    defparam i15638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15639_3_lut (.I0(Kp[4]), .I1(\data_in_frame[3] [4]), .I2(n27771), 
            .I3(GND_net), .O(n28702));   // verilog/coms.v(127[12] 300[6])
    defparam i15639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15640_3_lut (.I0(Kp[3]), .I1(\data_in_frame[3] [3]), .I2(n27771), 
            .I3(GND_net), .O(n28703));   // verilog/coms.v(127[12] 300[6])
    defparam i15640_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15641_3_lut (.I0(Kp[2]), .I1(\data_in_frame[3] [2]), .I2(n27771), 
            .I3(GND_net), .O(n28704));   // verilog/coms.v(127[12] 300[6])
    defparam i15641_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15642_3_lut (.I0(Kp[1]), .I1(\data_in_frame[3] [1]), .I2(n27771), 
            .I3(GND_net), .O(n28705));   // verilog/coms.v(127[12] 300[6])
    defparam i15642_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15643_3_lut (.I0(\data_in[3] [7]), .I1(rx_data[7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28706));   // verilog/coms.v(127[12] 300[6])
    defparam i15643_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15644_3_lut (.I0(\data_in[3] [6]), .I1(rx_data[6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28707));   // verilog/coms.v(127[12] 300[6])
    defparam i15644_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15645_3_lut (.I0(\data_in[3] [5]), .I1(rx_data[5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28708));   // verilog/coms.v(127[12] 300[6])
    defparam i15645_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15646_3_lut (.I0(\data_in[3] [4]), .I1(rx_data[4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28709));   // verilog/coms.v(127[12] 300[6])
    defparam i15646_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_8 (.CI(n40509), 
            .I0(GND_net), .I1(n27_adj_5016), .CO(n40510));
    SB_LUT4 encoder0_position_31__I_0_i978_3_lut (.I0(n1431), .I1(n1498), 
            .I2(n1455), .I3(GND_net), .O(n1530));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_7_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n28_adj_5017), .I3(n40508), .O(n28)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n5722), 
            .D(n683), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_7 (.CI(n40508), 
            .I0(GND_net), .I1(n28_adj_5017), .CO(n40509));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_6_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n29_adj_5018), .I3(n40507), .O(n29)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_6 (.CI(n40507), 
            .I0(GND_net), .I1(n29_adj_5018), .CO(n40508));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_5_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n30_adj_5019), .I3(n40506), .O(n30)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_5 (.CI(n40506), 
            .I0(GND_net), .I1(n30_adj_5019), .CO(n40507));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_4_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n31_adj_5020), .I3(n40505), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15647_3_lut (.I0(\data_in[3] [3]), .I1(rx_data[3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28710));   // verilog/coms.v(127[12] 300[6])
    defparam i15647_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_4 (.CI(n40505), 
            .I0(GND_net), .I1(n31_adj_5020), .CO(n40506));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_3_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n32_adj_5021), .I3(n40504), .O(n32)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_3 (.CI(n40504), 
            .I0(GND_net), .I1(n32_adj_5021), .CO(n40505));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_add_3_2_lut (.I0(GND_net), 
            .I1(GND_net), .I2(n33_adj_5022), .I3(VCC_net), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_unary_minus_2_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_unary_minus_2_add_3_2 (.CI(VCC_net), 
            .I0(GND_net), .I1(n33_adj_5022), .CO(n40504));
    SB_CARRY encoder0_position_31__I_0_add_1235_15 (.CI(n39762), .I0(n1821), 
            .I1(VCC_net), .CO(n39763));
    SB_LUT4 i15648_3_lut (.I0(\data_in[3] [2]), .I1(rx_data[2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28711));   // verilog/coms.v(127[12] 300[6])
    defparam i15648_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1235_14_lut (.I0(GND_net), .I1(n1822), 
            .I2(VCC_net), .I3(n39761), .O(n1889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_77_8 (.CI(n39026), .I0(encoder1_position[9]), .I1(GND_net), 
            .CO(n39027));
    SB_LUT4 i15649_3_lut (.I0(\data_in[3] [1]), .I1(rx_data[1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28712));   // verilog/coms.v(127[12] 300[6])
    defparam i15649_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1235_14 (.CI(n39761), .I0(n1822), 
            .I1(VCC_net), .CO(n39762));
    SB_LUT4 i15650_3_lut (.I0(\data_in[3] [0]), .I1(rx_data[0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28713));   // verilog/coms.v(127[12] 300[6])
    defparam i15650_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15651_3_lut (.I0(\data_in[2] [7]), .I1(\data_in[3] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28714));   // verilog/coms.v(127[12] 300[6])
    defparam i15651_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15652_3_lut (.I0(\data_in[2] [6]), .I1(\data_in[3] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28715));   // verilog/coms.v(127[12] 300[6])
    defparam i15652_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15653_3_lut (.I0(\data_in[2] [5]), .I1(\data_in[3] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28716));   // verilog/coms.v(127[12] 300[6])
    defparam i15653_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36149_1_lut (.I0(n2742), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51102));
    defparam i36149_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15654_3_lut (.I0(\data_in[2] [4]), .I1(\data_in[3] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28717));   // verilog/coms.v(127[12] 300[6])
    defparam i15654_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15655_3_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28718));   // verilog/coms.v(127[12] 300[6])
    defparam i15655_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15656_3_lut (.I0(\data_in[2] [2]), .I1(\data_in[3] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28719));   // verilog/coms.v(127[12] 300[6])
    defparam i15656_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15657_3_lut (.I0(\data_in[2] [1]), .I1(\data_in[3] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28720));   // verilog/coms.v(127[12] 300[6])
    defparam i15657_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15658_3_lut (.I0(\data_in[2] [0]), .I1(\data_in[3] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28721));   // verilog/coms.v(127[12] 300[6])
    defparam i15658_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15659_3_lut (.I0(\data_in[1] [7]), .I1(\data_in[2] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28722));   // verilog/coms.v(127[12] 300[6])
    defparam i15659_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15660_3_lut (.I0(\data_in[1] [6]), .I1(\data_in[2] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28723));   // verilog/coms.v(127[12] 300[6])
    defparam i15660_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15661_3_lut (.I0(\data_in[1] [5]), .I1(\data_in[2] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28724));   // verilog/coms.v(127[12] 300[6])
    defparam i15661_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15662_3_lut (.I0(\data_in[1] [4]), .I1(\data_in[2] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28725));   // verilog/coms.v(127[12] 300[6])
    defparam i15662_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15663_3_lut (.I0(\data_in[1] [3]), .I1(\data_in[2] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28726));   // verilog/coms.v(127[12] 300[6])
    defparam i15663_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15664_3_lut (.I0(\data_in[1] [2]), .I1(\data_in[2] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28727));   // verilog/coms.v(127[12] 300[6])
    defparam i15664_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15665_3_lut (.I0(\data_in[1] [1]), .I1(\data_in[2] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28728));   // verilog/coms.v(127[12] 300[6])
    defparam i15665_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15666_3_lut (.I0(\data_in[1] [0]), .I1(\data_in[2] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28729));   // verilog/coms.v(127[12] 300[6])
    defparam i15666_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15667_3_lut (.I0(\data_in[0] [7]), .I1(\data_in[1] [7]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28730));   // verilog/coms.v(127[12] 300[6])
    defparam i15667_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15668_3_lut (.I0(\data_in[0] [6]), .I1(\data_in[1] [6]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28731));   // verilog/coms.v(127[12] 300[6])
    defparam i15668_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15669_3_lut (.I0(\data_in[0] [5]), .I1(\data_in[1] [5]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28732));   // verilog/coms.v(127[12] 300[6])
    defparam i15669_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15670_3_lut (.I0(\data_in[0] [4]), .I1(\data_in[1] [4]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28733));   // verilog/coms.v(127[12] 300[6])
    defparam i15670_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15671_3_lut (.I0(\data_in[0] [3]), .I1(\data_in[1] [3]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28734));   // verilog/coms.v(127[12] 300[6])
    defparam i15671_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15672_3_lut (.I0(\data_in[0] [2]), .I1(\data_in[1] [2]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28735));   // verilog/coms.v(127[12] 300[6])
    defparam i15672_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15673_3_lut (.I0(\data_in[0] [1]), .I1(\data_in[1] [1]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28736));   // verilog/coms.v(127[12] 300[6])
    defparam i15673_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15674_3_lut (.I0(IntegralLimit[23]), .I1(\data_in_frame[11] [7]), 
            .I2(n27771), .I3(GND_net), .O(n28737));   // verilog/coms.v(127[12] 300[6])
    defparam i15674_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1235_13_lut (.I0(GND_net), .I1(n1823), 
            .I2(VCC_net), .I3(n39760), .O(n1890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_13_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i26 (.Q(delay_counter[26]), .C(CLK_c), .E(n5722), 
            .D(n664), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 i15675_3_lut (.I0(IntegralLimit[22]), .I1(\data_in_frame[11] [6]), 
            .I2(n27771), .I3(GND_net), .O(n28738));   // verilog/coms.v(127[12] 300[6])
    defparam i15675_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15676_3_lut (.I0(IntegralLimit[21]), .I1(\data_in_frame[11] [5]), 
            .I2(n27771), .I3(GND_net), .O(n28739));   // verilog/coms.v(127[12] 300[6])
    defparam i15676_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i25 (.Q(delay_counter[25]), .C(CLK_c), .E(n5722), 
            .D(n665), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 i15677_3_lut (.I0(IntegralLimit[20]), .I1(\data_in_frame[11] [4]), 
            .I2(n27771), .I3(GND_net), .O(n28740));   // verilog/coms.v(127[12] 300[6])
    defparam i15677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15678_3_lut (.I0(IntegralLimit[19]), .I1(\data_in_frame[11] [3]), 
            .I2(n27771), .I3(GND_net), .O(n28741));   // verilog/coms.v(127[12] 300[6])
    defparam i15678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15679_3_lut (.I0(IntegralLimit[18]), .I1(\data_in_frame[11] [2]), 
            .I2(n27771), .I3(GND_net), .O(n28742));   // verilog/coms.v(127[12] 300[6])
    defparam i15679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15680_3_lut (.I0(IntegralLimit[17]), .I1(\data_in_frame[11] [1]), 
            .I2(n27771), .I3(GND_net), .O(n28743));   // verilog/coms.v(127[12] 300[6])
    defparam i15680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15681_3_lut (.I0(IntegralLimit[16]), .I1(\data_in_frame[11] [0]), 
            .I2(n27771), .I3(GND_net), .O(n28744));   // verilog/coms.v(127[12] 300[6])
    defparam i15681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15682_3_lut (.I0(IntegralLimit[15]), .I1(\data_in_frame[12] [7]), 
            .I2(n27771), .I3(GND_net), .O(n28745));   // verilog/coms.v(127[12] 300[6])
    defparam i15682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15683_3_lut (.I0(IntegralLimit[14]), .I1(\data_in_frame[12] [6]), 
            .I2(n27771), .I3(GND_net), .O(n28746));   // verilog/coms.v(127[12] 300[6])
    defparam i15683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15684_3_lut (.I0(IntegralLimit[13]), .I1(\data_in_frame[12] [5]), 
            .I2(n27771), .I3(GND_net), .O(n28747));   // verilog/coms.v(127[12] 300[6])
    defparam i15684_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n5722), 
            .D(n684), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 i15685_3_lut (.I0(IntegralLimit[12]), .I1(\data_in_frame[12] [4]), 
            .I2(n27771), .I3(GND_net), .O(n28748));   // verilog/coms.v(127[12] 300[6])
    defparam i15685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15686_3_lut (.I0(IntegralLimit[11]), .I1(\data_in_frame[12] [3]), 
            .I2(n27771), .I3(GND_net), .O(n28749));   // verilog/coms.v(127[12] 300[6])
    defparam i15686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15687_3_lut (.I0(IntegralLimit[10]), .I1(\data_in_frame[12] [2]), 
            .I2(n27771), .I3(GND_net), .O(n28750));   // verilog/coms.v(127[12] 300[6])
    defparam i15687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15688_3_lut (.I0(IntegralLimit[9]), .I1(\data_in_frame[12] [1]), 
            .I2(n27771), .I3(GND_net), .O(n28751));   // verilog/coms.v(127[12] 300[6])
    defparam i15688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15689_3_lut (.I0(IntegralLimit[8]), .I1(\data_in_frame[12] [0]), 
            .I2(n27771), .I3(GND_net), .O(n28752));   // verilog/coms.v(127[12] 300[6])
    defparam i15689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15690_3_lut (.I0(IntegralLimit[7]), .I1(\data_in_frame[13] [7]), 
            .I2(n27771), .I3(GND_net), .O(n28753));   // verilog/coms.v(127[12] 300[6])
    defparam i15690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15691_3_lut (.I0(IntegralLimit[6]), .I1(\data_in_frame[13] [6]), 
            .I2(n27771), .I3(GND_net), .O(n28754));   // verilog/coms.v(127[12] 300[6])
    defparam i15691_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1235_13 (.CI(n39760), .I0(n1823), 
            .I1(VCC_net), .CO(n39761));
    SB_LUT4 i15692_3_lut (.I0(IntegralLimit[5]), .I1(\data_in_frame[13] [5]), 
            .I2(n27771), .I3(GND_net), .O(n28755));   // verilog/coms.v(127[12] 300[6])
    defparam i15692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15693_3_lut (.I0(IntegralLimit[4]), .I1(\data_in_frame[13] [4]), 
            .I2(n27771), .I3(GND_net), .O(n28756));   // verilog/coms.v(127[12] 300[6])
    defparam i15693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1235_12_lut (.I0(GND_net), .I1(n1824), 
            .I2(VCC_net), .I3(n39759), .O(n1891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15694_3_lut (.I0(IntegralLimit[3]), .I1(\data_in_frame[13] [3]), 
            .I2(n27771), .I3(GND_net), .O(n28757));   // verilog/coms.v(127[12] 300[6])
    defparam i15694_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1235_12 (.CI(n39759), .I0(n1824), 
            .I1(VCC_net), .CO(n39760));
    SB_LUT4 i15695_3_lut (.I0(IntegralLimit[2]), .I1(\data_in_frame[13] [2]), 
            .I2(n27771), .I3(GND_net), .O(n28758));   // verilog/coms.v(127[12] 300[6])
    defparam i15695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15696_3_lut (.I0(IntegralLimit[1]), .I1(\data_in_frame[13] [1]), 
            .I2(n27771), .I3(GND_net), .O(n28759));   // verilog/coms.v(127[12] 300[6])
    defparam i15696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_77_7_lut (.I0(GND_net), .I1(encoder1_position[8]), .I2(GND_net), 
            .I3(n39025), .O(encoder1_position_scaled_23__N_58[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1235_11_lut (.I0(GND_net), .I1(n1825), 
            .I2(VCC_net), .I3(n39758), .O(n1892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35098_4_lut (.I0(state[0]), .I1(start), .I2(n34525), .I3(\neo_pixel_transmitter.done ), 
            .O(n49724));   // verilog/neopixel.v(35[12] 117[6])
    defparam i35098_4_lut.LUT_INIT = 16'hccdc;
    SB_LUT4 encoder0_position_31__I_0_add_766_11_lut (.I0(n50798), .I1(n1125), 
            .I2(VCC_net), .I3(n39654), .O(n1224)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i34946_2_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n49726));   // verilog/neopixel.v(35[12] 117[6])
    defparam i34946_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i15208_3_lut (.I0(PWMLimit[7]), .I1(\data_in_frame[10] [7]), 
            .I2(n27771), .I3(GND_net), .O(n28271));   // verilog/coms.v(127[12] 300[6])
    defparam i15208_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18_4_lut (.I0(n49726), .I1(n49724), .I2(state[1]), .I3(n34629), 
            .O(n42985));   // verilog/neopixel.v(35[12] 117[6])
    defparam i18_4_lut.LUT_INIT = 16'hcac0;
    SB_LUT4 i15702_3_lut (.I0(ID[1]), .I1(data[1]), .I2(n46808), .I3(GND_net), 
            .O(n28765));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i15702_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15209_3_lut (.I0(PWMLimit[6]), .I1(\data_in_frame[10] [6]), 
            .I2(n27771), .I3(GND_net), .O(n28272));   // verilog/coms.v(127[12] 300[6])
    defparam i15209_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15703_3_lut (.I0(ID[2]), .I1(data[2]), .I2(n46808), .I3(GND_net), 
            .O(n28766));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i15703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15704_3_lut (.I0(ID[3]), .I1(data[3]), .I2(n46808), .I3(GND_net), 
            .O(n28767));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i15704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15705_3_lut (.I0(ID[4]), .I1(data[4]), .I2(n46808), .I3(GND_net), 
            .O(n28768));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i15705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_766_10_lut (.I0(GND_net), .I1(n1126), 
            .I2(VCC_net), .I3(n39653), .O(n1193_adj_4956)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15706_3_lut (.I0(ID[5]), .I1(data[5]), .I2(n46808), .I3(GND_net), 
            .O(n28769));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i15706_3_lut.LUT_INIT = 16'hacac;
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n5722), 
            .D(n685), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 i15707_3_lut (.I0(ID[6]), .I1(data[6]), .I2(n46808), .I3(GND_net), 
            .O(n28770));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i15707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15708_3_lut (.I0(ID[7]), .I1(data[7]), .I2(n46808), .I3(GND_net), 
            .O(n28771));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i15708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35005_4_lut (.I0(n5_adj_4947), .I1(n6_adj_5041), .I2(n5855), 
            .I3(n1419), .O(n49758));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i35005_4_lut.LUT_INIT = 16'h080c;
    SB_LUT4 i49_4_lut (.I0(n49758), .I1(n5855), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(data_ready), .O(n43285));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i49_4_lut.LUT_INIT = 16'hcafa;
    SB_LUT4 i273_2_lut (.I0(n777), .I1(n26483), .I2(GND_net), .I3(GND_net), 
            .O(n1419));   // verilog/TinyFPGA_B.v(278[9] 284[12])
    defparam i273_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1680 (.I0(n5_adj_4947), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(n1419), .I3(read_N_321), .O(n25_adj_4889));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i1_4_lut_adj_1680.LUT_INIT = 16'h7350;
    SB_LUT4 i33899_2_lut (.I0(data_ready), .I1(\ID_READOUT_FSM.state [0]), 
            .I2(GND_net), .I3(GND_net), .O(n48793));
    defparam i33899_2_lut.LUT_INIT = 16'h8888;
    SB_DFFESR delay_counter_i0_i24 (.Q(delay_counter[24]), .C(CLK_c), .E(n5722), 
            .D(n666), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 i35936_4_lut (.I0(\ID_READOUT_FSM.state [1]), .I1(n5855), .I2(n48793), 
            .I3(n25_adj_4889), .O(n17_adj_4890));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i35936_4_lut.LUT_INIT = 16'h88ba;
    SB_LUT4 add_29_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(GND_net), 
            .I3(n39000), .O(n679)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_11 (.CI(n39758), .I0(n1825), 
            .I1(VCC_net), .CO(n39759));
    SB_CARRY encoder0_position_31__I_0_add_766_10 (.CI(n39653), .I0(n1126), 
            .I1(VCC_net), .CO(n39654));
    SB_LUT4 encoder0_position_31__I_0_add_766_9_lut (.I0(GND_net), .I1(n1127), 
            .I2(VCC_net), .I3(n39652), .O(n1194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_77_25_lut (.I0(GND_net), .I1(encoder1_position[26]), .I2(GND_net), 
            .I3(n39043), .O(encoder1_position_scaled_23__N_58[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_77_24_lut (.I0(GND_net), .I1(encoder1_position[25]), .I2(GND_net), 
            .I3(n39042), .O(encoder1_position_scaled_23__N_58[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_77_7 (.CI(n39025), .I0(encoder1_position[8]), .I1(GND_net), 
            .CO(n39026));
    SB_LUT4 add_29_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(GND_net), 
            .I3(n38992), .O(n687)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29974_4_lut (.I0(n7_adj_4961), .I1(state_adj_5100[0]), .I2(n6_adj_4984), 
            .I3(state_adj_5116[0]), .O(n44859));
    defparam i29974_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 i1_3_lut_adj_1681 (.I0(state_adj_5100[1]), .I1(read), .I2(n44120), 
            .I3(GND_net), .O(n12_adj_4957));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_3_lut_adj_1681.LUT_INIT = 16'ha2a2;
    SB_LUT4 i1_4_lut_adj_1682 (.I0(n34334), .I1(n12_adj_4957), .I2(state_adj_5100[0]), 
            .I3(n44120), .O(n43693));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1682.LUT_INIT = 16'h88a8;
    SB_LUT4 i15143_4_lut (.I0(state_7__N_4003[3]), .I1(data[2]), .I2(n4_adj_4914), 
            .I3(n26645), .O(n28206));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15143_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_29_13 (.CI(n39000), .I0(delay_counter[11]), .I1(GND_net), 
            .CO(n39001));
    SB_LUT4 encoder0_position_31__I_0_add_1235_10_lut (.I0(GND_net), .I1(n1826), 
            .I2(VCC_net), .I3(n39757), .O(n1893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_10 (.CI(n39757), .I0(n1826), 
            .I1(VCC_net), .CO(n39758));
    SB_CARRY encoder0_position_31__I_0_add_766_9 (.CI(n39652), .I0(n1127), 
            .I1(VCC_net), .CO(n39653));
    SB_CARRY add_77_24 (.CI(n39042), .I0(encoder1_position[25]), .I1(GND_net), 
            .CO(n39043));
    SB_LUT4 add_77_23_lut (.I0(GND_net), .I1(encoder1_position[24]), .I2(GND_net), 
            .I3(n39041), .O(encoder1_position_scaled_23__N_58[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15144_4_lut (.I0(state_7__N_4003[3]), .I1(data[1]), .I2(n10_adj_5039), 
            .I3(n26650), .O(n28207));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15144_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 unary_minus_4_inv_0_i8_1_lut (.I0(duty[7]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n18));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_77_23 (.CI(n39041), .I0(encoder1_position[24]), .I1(GND_net), 
            .CO(n39042));
    SB_LUT4 add_77_6_lut (.I0(GND_net), .I1(encoder1_position[7]), .I2(GND_net), 
            .I3(n39024), .O(encoder1_position_scaled_23__N_58[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_77_6 (.CI(n39024), .I0(encoder1_position[7]), .I1(GND_net), 
            .CO(n39025));
    SB_LUT4 add_77_5_lut (.I0(GND_net), .I1(encoder1_position[6]), .I2(GND_net), 
            .I3(n39023), .O(encoder1_position_scaled_23__N_58[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_77_5 (.CI(n39023), .I0(encoder1_position[6]), .I1(GND_net), 
            .CO(n39024));
    SB_LUT4 encoder0_position_31__I_0_add_766_8_lut (.I0(GND_net), .I1(n1128), 
            .I2(VCC_net), .I3(n39651), .O(n1195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_8 (.CI(n39651), .I0(n1128), 
            .I1(VCC_net), .CO(n39652));
    SB_LUT4 unary_minus_4_inv_0_i9_1_lut (.I0(duty[8]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n17));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36184_1_lut (.I0(n2841), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51137));
    defparam i36184_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_77_22_lut (.I0(GND_net), .I1(encoder1_position[23]), .I2(GND_net), 
            .I3(n39040), .O(encoder1_position_scaled_23__N_58[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_77_4_lut (.I0(GND_net), .I1(encoder1_position[5]), .I2(GND_net), 
            .I3(n39022), .O(encoder1_position_scaled_23__N_58[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n5722), 
            .D(n690), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY add_29_5 (.CI(n38992), .I0(delay_counter[3]), .I1(GND_net), 
            .CO(n38993));
    SB_LUT4 encoder0_position_31__I_0_add_1235_9_lut (.I0(GND_net), .I1(n1827), 
            .I2(VCC_net), .I3(n39756), .O(n1894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_77_22 (.CI(n39040), .I0(encoder1_position[23]), .I1(GND_net), 
            .CO(n39041));
    SB_LUT4 add_29_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(GND_net), 
            .I3(n38999), .O(n680)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_12_lut.LUT_INIT = 16'hC33C;
    SB_IO RX_pad (.PACKAGE_PIN(RX), .OUTPUT_ENABLE(VCC_net), .D_IN_0(RX_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam RX_pad.PIN_TYPE = 6'b000001;
    defparam RX_pad.PULLUP = 1'b0;
    defparam RX_pad.NEG_TRIGGER = 1'b0;
    defparam RX_pad.IO_STANDARD = "SB_LVCMOS";
    SB_CARRY add_29_12 (.CI(n38999), .I0(delay_counter[10]), .I1(GND_net), 
            .CO(n39000));
    SB_LUT4 encoder0_position_31__I_0_add_766_7_lut (.I0(GND_net), .I1(n1129), 
            .I2(GND_net), .I3(n39650), .O(n1196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_9 (.CI(n39756), .I0(n1827), 
            .I1(VCC_net), .CO(n39757));
    SB_LUT4 encoder0_position_31__I_0_i1039_3_lut (.I0(n1524), .I1(n1591), 
            .I2(n1554), .I3(GND_net), .O(n1623));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1039_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_766_7 (.CI(n39650), .I0(n1129), 
            .I1(GND_net), .CO(n39651));
    SB_CARRY add_77_4 (.CI(n39022), .I0(encoder1_position[5]), .I1(GND_net), 
            .CO(n39023));
    SB_LUT4 add_29_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(GND_net), 
            .I3(n38991), .O(n688)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_77_21_lut (.I0(GND_net), .I1(encoder1_position[22]), .I2(GND_net), 
            .I3(n39039), .O(encoder1_position_scaled_23__N_58[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_21_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i23 (.Q(delay_counter[23]), .C(CLK_c), .E(n5722), 
            .D(n667), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY add_77_21 (.CI(n39039), .I0(encoder1_position[22]), .I1(GND_net), 
            .CO(n39040));
    SB_LUT4 add_29_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(GND_net), 
            .I3(n38998), .O(n681)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1235_8_lut (.I0(GND_net), .I1(n1828), 
            .I2(VCC_net), .I3(n39755), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_77_3_lut (.I0(GND_net), .I1(encoder1_position[4]), .I2(GND_net), 
            .I3(n39021), .O(encoder1_position_scaled_23__N_58[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_77_3 (.CI(n39021), .I0(encoder1_position[4]), .I1(GND_net), 
            .CO(n39022));
    SB_CARRY encoder0_position_31__I_0_add_1235_8 (.CI(n39755), .I0(n1828), 
            .I1(VCC_net), .CO(n39756));
    SB_LUT4 encoder0_position_31__I_0_add_766_6_lut (.I0(GND_net), .I1(n1130), 
            .I2(GND_net), .I3(n39649), .O(n1197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_77_20_lut (.I0(GND_net), .I1(encoder1_position[21]), .I2(GND_net), 
            .I3(n39038), .O(encoder1_position_scaled_23__N_58[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1235_7_lut (.I0(GND_net), .I1(n1829), 
            .I2(GND_net), .I3(n39754), .O(n1896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_7 (.CI(n39754), .I0(n1829), 
            .I1(GND_net), .CO(n39755));
    SB_CARRY add_77_20 (.CI(n39038), .I0(encoder1_position[21]), .I1(GND_net), 
            .CO(n39039));
    SB_LUT4 add_77_2_lut (.I0(GND_net), .I1(encoder1_position[3]), .I2(encoder1_position_scaled_23__N_231), 
            .I3(GND_net), .O(encoder1_position_scaled_23__N_58[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_77_19_lut (.I0(GND_net), .I1(encoder1_position[20]), .I2(GND_net), 
            .I3(n39037), .O(encoder1_position_scaled_23__N_58[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1235_6_lut (.I0(GND_net), .I1(n1830), 
            .I2(GND_net), .I3(n39753), .O(n1897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_6 (.CI(n39753), .I0(n1830), 
            .I1(GND_net), .CO(n39754));
    SB_CARRY add_77_19 (.CI(n39037), .I0(encoder1_position[20]), .I1(GND_net), 
            .CO(n39038));
    SB_LUT4 add_77_9_lut (.I0(GND_net), .I1(encoder1_position[10]), .I2(GND_net), 
            .I3(n39027), .O(encoder1_position_scaled_23__N_58[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_77_2 (.CI(GND_net), .I0(encoder1_position[3]), .I1(encoder1_position_scaled_23__N_231), 
            .CO(n39021));
    SB_LUT4 add_77_18_lut (.I0(GND_net), .I1(encoder1_position[19]), .I2(GND_net), 
            .I3(n39036), .O(encoder1_position_scaled_23__N_58[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_4_inv_0_i10_1_lut (.I0(duty[9]), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n16));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_766_6 (.CI(n39649), .I0(n1130), 
            .I1(GND_net), .CO(n39650));
    SB_LUT4 i36103_1_lut (.I0(n2148), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51056));
    defparam i36103_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i11_1_lut (.I0(duty[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4887));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1235_5_lut (.I0(GND_net), .I1(n1831), 
            .I2(VCC_net), .I3(n39752), .O(n1898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_766_5_lut (.I0(GND_net), .I1(n1131), 
            .I2(VCC_net), .I3(n39648), .O(n1198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_766_5 (.CI(n39648), .I0(n1131), 
            .I1(VCC_net), .CO(n39649));
    SB_LUT4 encoder0_position_31__I_0_add_766_4_lut (.I0(GND_net), .I1(n1132), 
            .I2(GND_net), .I3(n39647), .O(n1199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_5 (.CI(n39752), .I0(n1831), 
            .I1(VCC_net), .CO(n39753));
    SB_LUT4 encoder1_position_scaled_23__I_2_4_lut (.I0(encoder1_position[0]), 
            .I1(encoder1_position[31]), .I2(encoder1_position[1]), .I3(encoder1_position[2]), 
            .O(encoder1_position_scaled_23__N_231));   // verilog/TinyFPGA_B.v(223[33:52])
    defparam encoder1_position_scaled_23__I_2_4_lut.LUT_INIT = 16'hccc8;
    SB_CARRY add_77_18 (.CI(n39036), .I0(encoder1_position[19]), .I1(GND_net), 
            .CO(n39037));
    SB_LUT4 encoder0_position_31__I_0_add_1235_4_lut (.I0(GND_net), .I1(n1832), 
            .I2(GND_net), .I3(n39751), .O(n1899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35980_1_lut (.I0(n1554), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50933));
    defparam i35980_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15145_3_lut (.I0(\data_in[0] [0]), .I1(\data_in[1] [0]), .I2(rx_data_ready), 
            .I3(GND_net), .O(n28208));   // verilog/coms.v(127[12] 300[6])
    defparam i15145_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_766_4 (.CI(n39647), .I0(n1132), 
            .I1(GND_net), .CO(n39648));
    SB_LUT4 add_77_17_lut (.I0(GND_net), .I1(encoder1_position[18]), .I2(GND_net), 
            .I3(n39035), .O(encoder1_position_scaled_23__N_58[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_766_3_lut (.I0(GND_net), .I1(n1133), 
            .I2(VCC_net), .I3(n39646), .O(n1200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1235_4 (.CI(n39751), .I0(n1832), 
            .I1(GND_net), .CO(n39752));
    SB_CARRY add_77_17 (.CI(n39035), .I0(encoder1_position[18]), .I1(GND_net), 
            .CO(n39036));
    SB_LUT4 add_77_16_lut (.I0(GND_net), .I1(encoder1_position[17]), .I2(GND_net), 
            .I3(n39034), .O(encoder1_position_scaled_23__N_58[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i977_3_lut (.I0(n1430), .I1(n1497), 
            .I2(n1455), .I3(GND_net), .O(n1529));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1235_3_lut (.I0(GND_net), .I1(n1833), 
            .I2(VCC_net), .I3(n39750), .O(n1900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_77_16 (.CI(n39034), .I0(encoder1_position[17]), .I1(GND_net), 
            .CO(n39035));
    SB_CARRY encoder0_position_31__I_0_add_766_3 (.CI(n39646), .I0(n1133), 
            .I1(VCC_net), .CO(n39647));
    SB_LUT4 encoder0_position_31__I_0_i1047_3_lut (.I0(n1532), .I1(n1599), 
            .I2(n1554), .I3(GND_net), .O(n1631));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_766_2_lut (.I0(GND_net), .I1(n936), 
            .I2(GND_net), .I3(VCC_net), .O(n1201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_766_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15146_3_lut (.I0(Kp[0]), .I1(\data_in_frame[3] [0]), .I2(n27771), 
            .I3(GND_net), .O(n28209));   // verilog/coms.v(127[12] 300[6])
    defparam i15146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15147_3_lut (.I0(Ki[0]), .I1(\data_in_frame[5] [0]), .I2(n27771), 
            .I3(GND_net), .O(n28210));   // verilog/coms.v(127[12] 300[6])
    defparam i15147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15148_3_lut (.I0(neopxl_color[0]), .I1(\data_in_frame[6] [0]), 
            .I2(n46360), .I3(GND_net), .O(n28211));   // verilog/coms.v(127[12] 300[6])
    defparam i15148_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_77_11 (.CI(n39029), .I0(encoder1_position[12]), .I1(GND_net), 
            .CO(n39030));
    SB_LUT4 unary_minus_4_inv_0_i12_1_lut (.I0(duty[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n14));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i13_1_lut (.I0(duty[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n13));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1235_3 (.CI(n39750), .I0(n1833), 
            .I1(VCC_net), .CO(n39751));
    SB_LUT4 i15249_3_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(timer[4]), 
            .I2(n43085), .I3(GND_net), .O(n28312));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15249_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_77_15_lut (.I0(GND_net), .I1(encoder1_position[16]), .I2(GND_net), 
            .I3(n39033), .O(encoder1_position_scaled_23__N_58[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_77_15 (.CI(n39033), .I0(encoder1_position[16]), .I1(GND_net), 
            .CO(n39034));
    SB_LUT4 i36216_1_lut (.I0(n2940), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51169));
    defparam i36216_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1235_2_lut (.I0(GND_net), .I1(n943), 
            .I2(GND_net), .I3(VCC_net), .O(n1901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1235_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_77_14_lut (.I0(GND_net), .I1(encoder1_position[15]), .I2(GND_net), 
            .I3(n39032), .O(encoder1_position_scaled_23__N_58[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35330_4_lut (.I0(n9_adj_4966), .I1(n7_adj_4964), .I2(pwm_counter[2]), 
            .I3(pwm_setpoint[2]), .O(n50283));
    defparam i35330_4_lut.LUT_INIT = 16'heffe;
    SB_CARRY add_77_14 (.CI(n39032), .I0(encoder1_position[15]), .I1(GND_net), 
            .CO(n39033));
    SB_LUT4 i15150_3_lut (.I0(control_mode[0]), .I1(\data_in_frame[1] [0]), 
            .I2(n27771), .I3(GND_net), .O(n28213));   // verilog/coms.v(127[12] 300[6])
    defparam i15150_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_766_2 (.CI(VCC_net), .I0(n936), 
            .I1(GND_net), .CO(n39646));
    SB_CARRY encoder0_position_31__I_0_add_1235_2 (.CI(VCC_net), .I0(n943), 
            .I1(GND_net), .CO(n39750));
    SB_LUT4 add_29_33_lut (.I0(GND_net), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(n39020), .O(n659)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_77_13_lut (.I0(GND_net), .I1(encoder1_position[14]), .I2(GND_net), 
            .I3(n39031), .O(encoder1_position_scaled_23__N_58[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_699_10_lut (.I0(GND_net), .I1(n1026), 
            .I2(VCC_net), .I3(n39645), .O(n1093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1168_17_lut (.I0(n50974), .I1(n1719), 
            .I2(VCC_net), .I3(n39749), .O(n1818)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1168_16_lut (.I0(GND_net), .I1(n1720), 
            .I2(VCC_net), .I3(n39748), .O(n1787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_699_9_lut (.I0(GND_net), .I1(n1027), 
            .I2(VCC_net), .I3(n39644), .O(n1094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_9 (.CI(n39644), .I0(n1027), 
            .I1(VCC_net), .CO(n39645));
    SB_LUT4 encoder0_position_31__I_0_add_565_8_lut (.I0(n861), .I1(n828), 
            .I2(VCC_net), .I3(n39539), .O(n927)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_8_lut.LUT_INIT = 16'h8228;
    SB_LUT4 unary_minus_4_inv_0_i14_1_lut (.I0(duty[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n12));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_699_8_lut (.I0(GND_net), .I1(n1028), 
            .I2(VCC_net), .I3(n39643), .O(n1095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_565_7_lut (.I0(GND_net), .I1(n829), 
            .I2(GND_net), .I3(n39538), .O(n896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_7 (.CI(n39538), .I0(n829), 
            .I1(GND_net), .CO(n39539));
    SB_LUT4 encoder0_position_31__I_0_add_565_6_lut (.I0(GND_net), .I1(n830), 
            .I2(GND_net), .I3(n39537), .O(n897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_6 (.CI(n39537), .I0(n830), 
            .I1(GND_net), .CO(n39538));
    SB_LUT4 add_29_32_lut (.I0(GND_net), .I1(delay_counter[30]), .I2(GND_net), 
            .I3(n39019), .O(n660)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_8 (.CI(n39643), .I0(n1028), 
            .I1(VCC_net), .CO(n39644));
    SB_LUT4 encoder0_position_31__I_0_add_565_5_lut (.I0(GND_net), .I1(n831), 
            .I2(VCC_net), .I3(n39536), .O(n898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_5 (.CI(n39536), .I0(n831), 
            .I1(VCC_net), .CO(n39537));
    SB_LUT4 encoder0_position_31__I_0_add_699_7_lut (.I0(GND_net), .I1(n1029), 
            .I2(GND_net), .I3(n39642), .O(n1096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_565_4_lut (.I0(GND_net), .I1(n832), 
            .I2(GND_net), .I3(n39535), .O(n899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_4_inv_0_i15_1_lut (.I0(duty[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n11));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_699_7 (.CI(n39642), .I0(n1029), 
            .I1(GND_net), .CO(n39643));
    SB_IO ENCODER1_B_pad (.PACKAGE_PIN(ENCODER1_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_B_pad.PULLUP = 1'b0;
    defparam ENCODER1_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER1_A_pad (.PACKAGE_PIN(ENCODER1_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER1_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER1_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER1_A_pad.PULLUP = 1'b0;
    defparam ENCODER1_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER1_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_B_pad (.PACKAGE_PIN(ENCODER0_B), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_B_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_B_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_B_pad.PULLUP = 1'b0;
    defparam ENCODER0_B_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_B_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ENCODER0_A_pad (.PACKAGE_PIN(ENCODER0_A), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(ENCODER0_A_N));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ENCODER0_A_pad.PIN_TYPE = 6'b000001;
    defparam ENCODER0_A_pad.PULLUP = 1'b0;
    defparam ENCODER0_A_pad.NEG_TRIGGER = 1'b0;
    defparam ENCODER0_A_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO CLK_pad (.PACKAGE_PIN(CLK), .OUTPUT_ENABLE(VCC_net), .GLOBAL_BUFFER_OUTPUT(CLK_c));   // verilog/TinyFPGA_B.v(3[9:12])
    defparam CLK_pad.PIN_TYPE = 6'b000001;
    defparam CLK_pad.PULLUP = 1'b0;
    defparam CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHA_pad (.PACKAGE_PIN(INHA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHA_pad.PIN_TYPE = 6'b011001;
    defparam INHA_pad.PULLUP = 1'b0;
    defparam INHA_pad.NEG_TRIGGER = 1'b0;
    defparam INHA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLA_pad (.PACKAGE_PIN(INLA), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLA_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLA_pad.PIN_TYPE = 6'b011001;
    defparam INLA_pad.PULLUP = 1'b0;
    defparam INLA_pad.NEG_TRIGGER = 1'b0;
    defparam INLA_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHB_pad (.PACKAGE_PIN(INHB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHB_pad.PIN_TYPE = 6'b011001;
    defparam INHB_pad.PULLUP = 1'b0;
    defparam INHB_pad.NEG_TRIGGER = 1'b0;
    defparam INHB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INLB_pad (.PACKAGE_PIN(INLB), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INLB_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INLB_pad.PIN_TYPE = 6'b011001;
    defparam INLB_pad.PULLUP = 1'b0;
    defparam INLB_pad.NEG_TRIGGER = 1'b0;
    defparam INLB_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO INHC_pad (.PACKAGE_PIN(INHC), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(INHC_c)) /* synthesis IO_FF_OUT=TRUE */ ;   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam INHC_pad.PIN_TYPE = 6'b011001;
    defparam INHC_pad.PULLUP = 1'b0;
    defparam INHC_pad.NEG_TRIGGER = 1'b0;
    defparam INHC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO CS_CLK_pad (.PACKAGE_PIN(CS_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam CS_CLK_pad.PIN_TYPE = 6'b011001;
    defparam CS_CLK_pad.PULLUP = 1'b0;
    defparam CS_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam CS_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 unary_minus_4_inv_0_i16_1_lut (.I0(duty[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n10));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_IO DE_pad (.PACKAGE_PIN(DE), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(DE_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DE_pad.PIN_TYPE = 6'b011001;
    defparam DE_pad.PULLUP = 1'b0;
    defparam DE_pad.NEG_TRIGGER = 1'b0;
    defparam DE_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_31__I_0_i974_3_lut (.I0(n1427), .I1(n1494), 
            .I2(n1455), .I3(GND_net), .O(n1526));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i974_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i973_3_lut (.I0(n1426), .I1(n1493), 
            .I2(n1455), .I3(GND_net), .O(n1525));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i973_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i972_3_lut (.I0(n1425), .I1(n1492), 
            .I2(n1455), .I3(GND_net), .O(n1524));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i972_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i981_3_lut (.I0(n939), .I1(n1501), 
            .I2(n1455), .I3(GND_net), .O(n1533));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i980_3_lut (.I0(n1433), .I1(n1500), 
            .I2(n1455), .I3(GND_net), .O(n1532));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i979_3_lut (.I0(n1432), .I1(n1499), 
            .I2(n1455), .I3(GND_net), .O(n1531));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i903_3_lut (.I0(n1324), .I1(n1391), 
            .I2(n1356), .I3(GND_net), .O(n1423));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i903_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i906_3_lut (.I0(n1327), .I1(n1394), 
            .I2(n1356), .I3(GND_net), .O(n1426));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i906_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i905_3_lut (.I0(n1326), .I1(n1393), 
            .I2(n1356), .I3(GND_net), .O(n1425));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i905_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i904_3_lut (.I0(n1325), .I1(n1392), 
            .I2(n1356), .I3(GND_net), .O(n1424));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i904_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i911_3_lut (.I0(n1332), .I1(n1399), 
            .I2(n1356), .I3(GND_net), .O(n1431));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i910_3_lut (.I0(n1331), .I1(n1398), 
            .I2(n1356), .I3(GND_net), .O(n1430));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i909_3_lut (.I0(n1330), .I1(n1397), 
            .I2(n1356), .I3(GND_net), .O(n1429));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i907_3_lut (.I0(n1328), .I1(n1395), 
            .I2(n1356), .I3(GND_net), .O(n1427));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i907_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i836_3_lut (.I0(n1225), .I1(n1292), 
            .I2(n1257), .I3(GND_net), .O(n1324));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i836_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i843_3_lut (.I0(n1232), .I1(n1299), 
            .I2(n1257), .I3(GND_net), .O(n1331));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i842_3_lut (.I0(n1231), .I1(n1298), 
            .I2(n1257), .I3(GND_net), .O(n1330));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i841_3_lut (.I0(n1230), .I1(n1297), 
            .I2(n1257), .I3(GND_net), .O(n1329));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i840_3_lut (.I0(n1229), .I1(n1296), 
            .I2(n1257), .I3(GND_net), .O(n1328));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i840_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i839_3_lut (.I0(n1228), .I1(n1295), 
            .I2(n1257), .I3(GND_net), .O(n1327));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i839_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i838_3_lut (.I0(n1227), .I1(n1294), 
            .I2(n1257), .I3(GND_net), .O(n1326));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i838_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i837_3_lut (.I0(n1226), .I1(n1293), 
            .I2(n1257), .I3(GND_net), .O(n1325));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i837_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i775_3_lut (.I0(n1132), .I1(n1199), 
            .I2(n1158), .I3(GND_net), .O(n1231));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i775_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i774_3_lut (.I0(n1131), .I1(n1198), 
            .I2(n1158), .I3(GND_net), .O(n1230));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15210_3_lut (.I0(PWMLimit[5]), .I1(\data_in_frame[10] [5]), 
            .I2(n27771), .I3(GND_net), .O(n28273));   // verilog/coms.v(127[12] 300[6])
    defparam i15210_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15211_3_lut (.I0(PWMLimit[4]), .I1(\data_in_frame[10] [4]), 
            .I2(n27771), .I3(GND_net), .O(n28274));   // verilog/coms.v(127[12] 300[6])
    defparam i15211_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15212_3_lut (.I0(PWMLimit[3]), .I1(\data_in_frame[10] [3]), 
            .I2(n27771), .I3(GND_net), .O(n28275));   // verilog/coms.v(127[12] 300[6])
    defparam i15212_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_77_13 (.CI(n39031), .I0(encoder1_position[14]), .I1(GND_net), 
            .CO(n39032));
    SB_CARRY encoder0_position_31__I_0_add_565_4 (.CI(n39535), .I0(n832), 
            .I1(GND_net), .CO(n39536));
    SB_CARRY encoder0_position_31__I_0_add_1168_16 (.CI(n39748), .I0(n1720), 
            .I1(VCC_net), .CO(n39749));
    SB_LUT4 i15213_3_lut (.I0(PWMLimit[2]), .I1(\data_in_frame[10] [2]), 
            .I2(n27771), .I3(GND_net), .O(n28276));   // verilog/coms.v(127[12] 300[6])
    defparam i15213_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_29_32 (.CI(n39019), .I0(delay_counter[30]), .I1(GND_net), 
            .CO(n39020));
    SB_LUT4 i15214_3_lut (.I0(PWMLimit[1]), .I1(\data_in_frame[10] [1]), 
            .I2(n27771), .I3(GND_net), .O(n28277));   // verilog/coms.v(127[12] 300[6])
    defparam i15214_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1168_15_lut (.I0(GND_net), .I1(n1721), 
            .I2(VCC_net), .I3(n39747), .O(n1788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_77_12_lut (.I0(GND_net), .I1(encoder1_position[13]), .I2(GND_net), 
            .I3(n39030), .O(encoder1_position_scaled_23__N_58[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15215_3_lut (.I0(control_mode[7]), .I1(\data_in_frame[1] [7]), 
            .I2(n27771), .I3(GND_net), .O(n28278));   // verilog/coms.v(127[12] 300[6])
    defparam i15215_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1168_15 (.CI(n39747), .I0(n1721), 
            .I1(VCC_net), .CO(n39748));
    SB_LUT4 encoder0_position_31__I_0_i773_3_lut (.I0(n1130), .I1(n1197), 
            .I2(n1158), .I3(GND_net), .O(n1229));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i773_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_699_6_lut (.I0(GND_net), .I1(n1030), 
            .I2(GND_net), .I3(n39641), .O(n1097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i772_3_lut (.I0(n1129), .I1(n1196), 
            .I2(n1158), .I3(GND_net), .O(n1228));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i772_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15216_3_lut (.I0(control_mode[6]), .I1(\data_in_frame[1] [6]), 
            .I2(n27771), .I3(GND_net), .O(n28279));   // verilog/coms.v(127[12] 300[6])
    defparam i15216_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15217_3_lut (.I0(control_mode[5]), .I1(\data_in_frame[1] [5]), 
            .I2(n27771), .I3(GND_net), .O(n28280));   // verilog/coms.v(127[12] 300[6])
    defparam i15217_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1168_14_lut (.I0(GND_net), .I1(n1722), 
            .I2(VCC_net), .I3(n39746), .O(n1789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15218_3_lut (.I0(control_mode[4]), .I1(\data_in_frame[1] [4]), 
            .I2(n27771), .I3(GND_net), .O(n28281));   // verilog/coms.v(127[12] 300[6])
    defparam i15218_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_699_6 (.CI(n39641), .I0(n1030), 
            .I1(GND_net), .CO(n39642));
    SB_CARRY encoder0_position_31__I_0_add_1168_14 (.CI(n39746), .I0(n1722), 
            .I1(VCC_net), .CO(n39747));
    SB_LUT4 encoder0_position_31__I_0_add_1168_13_lut (.I0(GND_net), .I1(n1723), 
            .I2(VCC_net), .I3(n39745), .O(n1790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15219_3_lut (.I0(control_mode[3]), .I1(\data_in_frame[1] [3]), 
            .I2(n27771), .I3(GND_net), .O(n28282));   // verilog/coms.v(127[12] 300[6])
    defparam i15219_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_565_3_lut (.I0(GND_net), .I1(n833), 
            .I2(VCC_net), .I3(n39534), .O(n900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_3 (.CI(n39534), .I0(n833), 
            .I1(VCC_net), .CO(n39535));
    SB_CARRY encoder0_position_31__I_0_add_1168_13 (.CI(n39745), .I0(n1723), 
            .I1(VCC_net), .CO(n39746));
    SB_LUT4 unary_minus_4_inv_0_i17_1_lut (.I0(duty[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i18_1_lut (.I0(duty[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n8));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15220_3_lut (.I0(control_mode[2]), .I1(\data_in_frame[1] [2]), 
            .I2(n27771), .I3(GND_net), .O(n28283));   // verilog/coms.v(127[12] 300[6])
    defparam i15220_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_77_12 (.CI(n39030), .I0(encoder1_position[13]), .I1(GND_net), 
            .CO(n39031));
    SB_LUT4 i15221_3_lut (.I0(control_mode[1]), .I1(\data_in_frame[1] [1]), 
            .I2(n27771), .I3(GND_net), .O(n28284));   // verilog/coms.v(127[12] 300[6])
    defparam i15221_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15222_3_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(timer[31]), 
            .I2(n43085), .I3(GND_net), .O(n28285));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15222_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1168_12_lut (.I0(GND_net), .I1(n1724), 
            .I2(VCC_net), .I3(n39744), .O(n1791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_699_5_lut (.I0(GND_net), .I1(n1031), 
            .I2(VCC_net), .I3(n39640), .O(n1098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_12 (.CI(n39744), .I0(n1724), 
            .I1(VCC_net), .CO(n39745));
    SB_LUT4 i15223_3_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(timer[30]), 
            .I2(n43085), .I3(GND_net), .O(n28286));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15223_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15224_3_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(timer[29]), 
            .I2(n43085), .I3(GND_net), .O(n28287));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15224_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_699_5 (.CI(n39640), .I0(n1031), 
            .I1(VCC_net), .CO(n39641));
    SB_LUT4 encoder0_position_31__I_0_add_565_2_lut (.I0(GND_net), .I1(n834), 
            .I2(GND_net), .I3(VCC_net), .O(n901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_565_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_77_11_lut (.I0(GND_net), .I1(encoder1_position[12]), .I2(GND_net), 
            .I3(n39029), .O(encoder1_position_scaled_23__N_58[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1168_11_lut (.I0(GND_net), .I1(n1725), 
            .I2(VCC_net), .I3(n39743), .O(n1792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_77_9 (.CI(n39027), .I0(encoder1_position[10]), .I1(GND_net), 
            .CO(n39028));
    SB_CARRY encoder0_position_31__I_0_add_1168_11 (.CI(n39743), .I0(n1725), 
            .I1(VCC_net), .CO(n39744));
    SB_LUT4 encoder0_position_31__I_0_add_699_4_lut (.I0(GND_net), .I1(n1032), 
            .I2(GND_net), .I3(n39639), .O(n1099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_4 (.CI(n39639), .I0(n1032), 
            .I1(GND_net), .CO(n39640));
    SB_LUT4 encoder0_position_31__I_0_i771_3_lut (.I0(n1128), .I1(n1195), 
            .I2(n1158), .I3(GND_net), .O(n1227));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i771_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_699_3_lut (.I0(GND_net), .I1(n1033), 
            .I2(VCC_net), .I3(n39638), .O(n1100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_565_2 (.CI(VCC_net), .I0(n834), 
            .I1(GND_net), .CO(n39534));
    SB_LUT4 encoder0_position_31__I_0_add_1168_10_lut (.I0(GND_net), .I1(n1726), 
            .I2(VCC_net), .I3(n39742), .O(n1793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_10 (.CI(n39742), .I0(n1726), 
            .I1(VCC_net), .CO(n39743));
    SB_CARRY encoder0_position_31__I_0_add_699_3 (.CI(n39638), .I0(n1033), 
            .I1(VCC_net), .CO(n39639));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_25_lut (.I0(GND_net), .I1(encoder0_position_scaled[23]), 
            .I2(n2), .I3(n39323), .O(displacement_23__N_82[23])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_699_2_lut (.I0(GND_net), .I1(n935), 
            .I2(GND_net), .I3(VCC_net), .O(n1101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_699_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_77_10_lut (.I0(GND_net), .I1(encoder1_position[11]), .I2(GND_net), 
            .I3(n39028), .O(encoder1_position_scaled_23__N_58[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1168_9_lut (.I0(GND_net), .I1(n1727), 
            .I2(VCC_net), .I3(n39741), .O(n1794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_29_31_lut (.I0(GND_net), .I1(delay_counter[29]), .I2(GND_net), 
            .I3(n39018), .O(n661)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_699_2 (.CI(VCC_net), .I0(n935), 
            .I1(GND_net), .CO(n39638));
    SB_CARRY add_77_10 (.CI(n39028), .I0(encoder1_position[11]), .I1(GND_net), 
            .CO(n39029));
    SB_CARRY encoder0_position_31__I_0_add_1168_9 (.CI(n39741), .I0(n1727), 
            .I1(VCC_net), .CO(n39742));
    SB_LUT4 encoder0_position_31__I_0_add_632_9_lut (.I0(n960), .I1(n927), 
            .I2(VCC_net), .I3(n39637), .O(n1026)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1168_8_lut (.I0(GND_net), .I1(n1728), 
            .I2(VCC_net), .I3(n39740), .O(n1795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_8 (.CI(n39740), .I0(n1728), 
            .I1(VCC_net), .CO(n39741));
    SB_LUT4 encoder0_position_31__I_0_add_632_8_lut (.I0(GND_net), .I1(n928), 
            .I2(VCC_net), .I3(n39636), .O(n995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i22 (.Q(delay_counter[22]), .C(CLK_c), .E(n5722), 
            .D(n668), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY encoder0_position_31__I_0_add_632_8 (.CI(n39636), .I0(n928), 
            .I1(VCC_net), .CO(n39637));
    SB_LUT4 encoder0_position_31__I_0_add_1168_7_lut (.I0(GND_net), .I1(n1729), 
            .I2(GND_net), .I3(n39739), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_24_lut (.I0(GND_net), .I1(encoder0_position_scaled[22]), 
            .I2(n3_adj_4936), .I3(n39322), .O(displacement_23__N_82[22])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_31 (.CI(n39018), .I0(delay_counter[29]), .I1(GND_net), 
            .CO(n39019));
    SB_LUT4 encoder0_position_31__I_0_add_632_7_lut (.I0(GND_net), .I1(n929), 
            .I2(GND_net), .I3(n39635), .O(n996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_7 (.CI(n39635), .I0(n929), 
            .I1(GND_net), .CO(n39636));
    SB_LUT4 i15225_3_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(timer[28]), 
            .I2(n43085), .I3(GND_net), .O(n28288));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15225_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i770_3_lut (.I0(n1127), .I1(n1194), 
            .I2(n1158), .I3(GND_net), .O(n1226));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i770_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i777_3_lut (.I0(n936), .I1(n1201), 
            .I2(n1158), .I3(GND_net), .O(n1233));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i777_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i776_3_lut (.I0(n1133), .I1(n1200), 
            .I2(n1158), .I3(GND_net), .O(n1232));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21468_3_lut (.I0(n937), .I1(n1232), .I2(n1233), .I3(GND_net), 
            .O(n34531));
    defparam i21468_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_adj_1683 (.I0(n1226), .I1(n1227), .I2(n1228), .I3(GND_net), 
            .O(n47239));
    defparam i1_3_lut_adj_1683.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1684 (.I0(n1229), .I1(n34531), .I2(n1230), .I3(n1231), 
            .O(n45026));
    defparam i1_4_lut_adj_1684.LUT_INIT = 16'ha080;
    SB_LUT4 i35867_4_lut (.I0(n1225), .I1(n1224), .I2(n45026), .I3(n47239), 
            .O(n1257));
    defparam i35867_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i22_3_lut (.I0(encoder0_position[21]), 
            .I1(n12_adj_4930), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n937));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i845_3_lut (.I0(n937), .I1(n1301), 
            .I2(n1257), .I3(GND_net), .O(n1333));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i844_3_lut (.I0(n1233), .I1(n1300), 
            .I2(n1257), .I3(GND_net), .O(n1332));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21412_3_lut (.I0(n938), .I1(n1332), .I2(n1333), .I3(GND_net), 
            .O(n34475));
    defparam i21412_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1685 (.I0(n1325), .I1(n1326), .I2(n1327), .I3(n1328), 
            .O(n46953));
    defparam i1_4_lut_adj_1685.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1686 (.I0(n1329), .I1(n34475), .I2(n1330), .I3(n1331), 
            .O(n45023));
    defparam i1_4_lut_adj_1686.LUT_INIT = 16'ha080;
    SB_LUT4 i35883_4_lut (.I0(n45023), .I1(n1323), .I2(n1324), .I3(n46953), 
            .O(n1356));
    defparam i35883_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i21_3_lut (.I0(encoder0_position[20]), 
            .I1(n13_adj_4929), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n938));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i913_3_lut (.I0(n938), .I1(n1401), 
            .I2(n1356), .I3(GND_net), .O(n1433));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i912_3_lut (.I0(n1333), .I1(n1400), 
            .I2(n1356), .I3(GND_net), .O(n1432));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i20_3_lut (.I0(encoder0_position[19]), 
            .I1(n14_adj_4928), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n939));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21408_3_lut (.I0(n939), .I1(n1432), .I2(n1433), .I3(GND_net), 
            .O(n34471));
    defparam i21408_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1687 (.I0(n1427), .I1(n1428), .I2(GND_net), .I3(GND_net), 
            .O(n47247));
    defparam i1_2_lut_adj_1687.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1688 (.I0(n1429), .I1(n34471), .I2(n1430), .I3(n1431), 
            .O(n45042));
    defparam i1_4_lut_adj_1688.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1689 (.I0(n1424), .I1(n1425), .I2(n1426), .I3(n47247), 
            .O(n47253));
    defparam i1_4_lut_adj_1689.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_632_6_lut (.I0(GND_net), .I1(n930), 
            .I2(GND_net), .I3(n39634), .O(n997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35845_1_lut (.I0(n1158), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50798));
    defparam i35845_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_1168_7 (.CI(n39739), .I0(n1729), 
            .I1(GND_net), .CO(n39740));
    SB_CARRY encoder0_position_31__I_0_add_632_6 (.CI(n39634), .I0(n930), 
            .I1(GND_net), .CO(n39635));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_24 (.CI(n39322), .I0(encoder0_position_scaled[22]), 
            .I1(n3_adj_4936), .CO(n39323));
    SB_LUT4 i35955_4_lut (.I0(n1423), .I1(n1422), .I2(n47253), .I3(n45042), 
            .O(n1455));
    defparam i35955_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_632_5_lut (.I0(GND_net), .I1(n931), 
            .I2(VCC_net), .I3(n39633), .O(n998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_23_lut (.I0(GND_net), .I1(encoder0_position_scaled[21]), 
            .I2(n4_adj_4937), .I3(n39321), .O(displacement_23__N_82[21])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i908_3_lut (.I0(n1329), .I1(n1396), 
            .I2(n1356), .I3(GND_net), .O(n1428));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i908_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_29_11 (.CI(n38998), .I0(delay_counter[9]), .I1(GND_net), 
            .CO(n38999));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_23 (.CI(n39321), .I0(encoder0_position_scaled[21]), 
            .I1(n4_adj_4937), .CO(n39322));
    SB_LUT4 add_29_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(GND_net), 
            .I3(n38997), .O(n682)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_10_lut.LUT_INIT = 16'hC33C;
    SB_DFF displacement_i23 (.Q(displacement[23]), .C(CLK_c), .D(displacement_23__N_82[23]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_LUT4 i36002_1_lut (.I0(n1653), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50955));
    defparam i36002_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i19_1_lut (.I0(duty[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4886));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36250_1_lut (.I0(n3039), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51203));
    defparam i36250_1_lut.LUT_INIT = 16'h5555;
    SB_DFF displacement_i22 (.Q(displacement[22]), .C(CLK_c), .D(displacement_23__N_82[22]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i21 (.Q(displacement[21]), .C(CLK_c), .D(displacement_23__N_82[21]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i20 (.Q(displacement[20]), .C(CLK_c), .D(displacement_23__N_82[20]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i19 (.Q(displacement[19]), .C(CLK_c), .D(displacement_23__N_82[19]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i18 (.Q(displacement[18]), .C(CLK_c), .D(displacement_23__N_82[18]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i17 (.Q(displacement[17]), .C(CLK_c), .D(displacement_23__N_82[17]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i16 (.Q(displacement[16]), .C(CLK_c), .D(displacement_23__N_82[16]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i15 (.Q(displacement[15]), .C(CLK_c), .D(displacement_23__N_82[15]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i14 (.Q(displacement[14]), .C(CLK_c), .D(displacement_23__N_82[14]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i13 (.Q(displacement[13]), .C(CLK_c), .D(displacement_23__N_82[13]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i12 (.Q(displacement[12]), .C(CLK_c), .D(displacement_23__N_82[12]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i11 (.Q(displacement[11]), .C(CLK_c), .D(displacement_23__N_82[11]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i10 (.Q(displacement[10]), .C(CLK_c), .D(displacement_23__N_82[10]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i9 (.Q(displacement[9]), .C(CLK_c), .D(displacement_23__N_82[9]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i8 (.Q(displacement[8]), .C(CLK_c), .D(displacement_23__N_82[8]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i7 (.Q(displacement[7]), .C(CLK_c), .D(displacement_23__N_82[7]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i6 (.Q(displacement[6]), .C(CLK_c), .D(displacement_23__N_82[6]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i5 (.Q(displacement[5]), .C(CLK_c), .D(displacement_23__N_82[5]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i4 (.Q(displacement[4]), .C(CLK_c), .D(displacement_23__N_82[4]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i3 (.Q(displacement[3]), .C(CLK_c), .D(displacement_23__N_82[3]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i2 (.Q(displacement[2]), .C(CLK_c), .D(displacement_23__N_82[2]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF displacement_i1 (.Q(displacement[1]), .C(CLK_c), .D(displacement_23__N_82[1]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i23 (.Q(encoder1_position_scaled[23]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[23]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i22 (.Q(encoder1_position_scaled[22]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[22]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i21 (.Q(encoder1_position_scaled[21]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[21]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i20 (.Q(encoder1_position_scaled[20]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[20]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i19 (.Q(encoder1_position_scaled[19]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[19]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i18 (.Q(encoder1_position_scaled[18]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[18]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i17 (.Q(encoder1_position_scaled[17]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[17]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i16 (.Q(encoder1_position_scaled[16]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[16]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i15 (.Q(encoder1_position_scaled[15]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[15]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i14 (.Q(encoder1_position_scaled[14]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[14]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i13 (.Q(encoder1_position_scaled[13]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[13]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i12 (.Q(encoder1_position_scaled[12]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[12]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i11 (.Q(encoder1_position_scaled[11]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[11]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i10 (.Q(encoder1_position_scaled[10]), 
           .C(CLK_c), .D(encoder1_position_scaled_23__N_58[10]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i9 (.Q(encoder1_position_scaled[9]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[9]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i8 (.Q(encoder1_position_scaled[8]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[8]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i7 (.Q(encoder1_position_scaled[7]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[7]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i6 (.Q(encoder1_position_scaled[6]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[6]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i5 (.Q(encoder1_position_scaled[5]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[5]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i4 (.Q(encoder1_position_scaled[4]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[4]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i3 (.Q(encoder1_position_scaled[3]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[3]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i2 (.Q(encoder1_position_scaled[2]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[2]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder1_position_scaled_i1 (.Q(encoder1_position_scaled[1]), .C(CLK_c), 
           .D(encoder1_position_scaled_23__N_58[1]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_LUT4 add_29_30_lut (.I0(GND_net), .I1(delay_counter[28]), .I2(GND_net), 
            .I3(n39017), .O(n662)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1168_6_lut (.I0(GND_net), .I1(n1730), 
            .I2(GND_net), .I3(n39738), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_6 (.CI(n39738), .I0(n1730), 
            .I1(GND_net), .CO(n39739));
    SB_LUT4 encoder0_position_31__I_0_i975_3_lut (.I0(n1428), .I1(n1495), 
            .I2(n1455), .I3(GND_net), .O(n1527));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 unary_minus_4_inv_0_i20_1_lut (.I0(duty[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n6));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i976_3_lut (.I0(n1429), .I1(n1496), 
            .I2(n1455), .I3(GND_net), .O(n1528));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1690 (.I0(n1528), .I1(n1527), .I2(GND_net), .I3(GND_net), 
            .O(n47151));
    defparam i1_2_lut_adj_1690.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_31__I_0_add_1168_5_lut (.I0(GND_net), .I1(n1731), 
            .I2(VCC_net), .I3(n39737), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_5 (.CI(n39633), .I0(n931), 
            .I1(VCC_net), .CO(n39634));
    SB_CARRY encoder0_position_31__I_0_add_1168_5 (.CI(n39737), .I0(n1731), 
            .I1(VCC_net), .CO(n39738));
    SB_LUT4 i15151_3_lut (.I0(PWMLimit[0]), .I1(\data_in_frame[10] [0]), 
            .I2(n27771), .I3(GND_net), .O(n28214));   // verilog/coms.v(127[12] 300[6])
    defparam i15151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21590_4_lut (.I0(n940), .I1(n1531), .I2(n1532), .I3(n1533), 
            .O(n34657));
    defparam i21590_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1691 (.I0(n1524), .I1(n1525), .I2(n1526), .I3(n47151), 
            .O(n47157));
    defparam i1_4_lut_adj_1691.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1692 (.I0(n1529), .I1(n47157), .I2(n34657), .I3(n1530), 
            .O(n47159));
    defparam i1_4_lut_adj_1692.LUT_INIT = 16'heccc;
    SB_LUT4 unary_minus_4_inv_0_i21_1_lut (.I0(duty[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n5));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_4_inv_0_i22_1_lut (.I0(duty[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35984_4_lut (.I0(n1522), .I1(n1521), .I2(n47159), .I3(n1523), 
            .O(n1554));
    defparam i35984_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 unary_minus_4_inv_0_i23_1_lut (.I0(duty[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n3));   // verilog/TinyFPGA_B.v(106[23:28])
    defparam unary_minus_4_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i19_3_lut (.I0(encoder0_position[18]), 
            .I1(n15_adj_4927), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n940));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1049_3_lut (.I0(n940), .I1(n1601), 
            .I2(n1554), .I3(GND_net), .O(n1633));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15226_3_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(timer[27]), 
            .I2(n43085), .I3(GND_net), .O(n28289));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15226_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1048_3_lut (.I0(n1533), .I1(n1600), 
            .I2(n1554), .I3(GND_net), .O(n1632));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15227_3_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(timer[26]), 
            .I2(n43085), .I3(GND_net), .O(n28290));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15227_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15228_3_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(timer[25]), 
            .I2(n43085), .I3(GND_net), .O(n28291));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15228_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21398_3_lut (.I0(n941), .I1(n1632), .I2(n1633), .I3(GND_net), 
            .O(n34461));
    defparam i21398_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1693 (.I0(n1625), .I1(n1627), .I2(n1626), .I3(n1628), 
            .O(n47263));
    defparam i1_4_lut_adj_1693.LUT_INIT = 16'hfffe;
    SB_LUT4 i15229_3_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(timer[24]), 
            .I2(n43085), .I3(GND_net), .O(n28292));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15229_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15230_3_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(timer[23]), 
            .I2(n43085), .I3(GND_net), .O(n28293));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15230_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_83_i1_4_lut (.I0(encoder1_position_scaled[0]), .I1(displacement[0]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[0]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i1_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_4_lut_adj_1694 (.I0(n1629), .I1(n34461), .I2(n1630), .I3(n1631), 
            .O(n45051));
    defparam i1_4_lut_adj_1694.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_31__I_0_add_1168_4_lut (.I0(GND_net), .I1(n1732), 
            .I2(GND_net), .I3(n39736), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_22_lut (.I0(GND_net), .I1(encoder0_position_scaled[20]), 
            .I2(n5_adj_4891), .I3(n39320), .O(displacement_23__N_82[20])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_22 (.CI(n39320), .I0(encoder0_position_scaled[20]), 
            .I1(n5_adj_4891), .CO(n39321));
    SB_DFF read_66 (.Q(read), .C(CLK_c), .D(n46845));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 i1_4_lut_adj_1695 (.I0(n1623), .I1(n45051), .I2(n1624), .I3(n47263), 
            .O(n47269));
    defparam i1_4_lut_adj_1695.LUT_INIT = 16'hfffe;
    SB_LUT4 i36006_4_lut (.I0(n1621), .I1(n1620), .I2(n1622), .I3(n47269), 
            .O(n1653));
    defparam i36006_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_83_i2_4_lut (.I0(encoder1_position_scaled[1]), .I1(displacement[1]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[1]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i2_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i1_1_lut (.I0(encoder1_position_scaled[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_4911));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_632_4_lut (.I0(GND_net), .I1(n932), 
            .I2(GND_net), .I3(n39632), .O(n999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_30 (.CI(n39017), .I0(delay_counter[28]), .I1(GND_net), 
            .CO(n39018));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_21_lut (.I0(GND_net), .I1(encoder0_position_scaled[19]), 
            .I2(n6_adj_4892), .I3(n39319), .O(displacement_23__N_82[19])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_83_i3_4_lut (.I0(encoder1_position_scaled[2]), .I1(displacement[2]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[2]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i3_4_lut.LUT_INIT = 16'h0aca;
    SB_CARRY add_29_4 (.CI(n38991), .I0(delay_counter[2]), .I1(GND_net), 
            .CO(n38992));
    SB_DFF encoder0_position_scaled_i23 (.Q(encoder0_position_scaled[23]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[23]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_LUT4 encoder0_position_31__I_0_mux_3_i18_3_lut (.I0(encoder0_position[17]), 
            .I1(n16_adj_4926), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n941));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_29_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(GND_net), 
            .I3(n38990), .O(n689)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_10 (.CI(n38997), .I0(delay_counter[8]), .I1(GND_net), 
            .CO(n38998));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_21 (.CI(n39319), .I0(encoder0_position_scaled[19]), 
            .I1(n6_adj_4892), .CO(n39320));
    SB_LUT4 add_29_29_lut (.I0(GND_net), .I1(delay_counter[27]), .I2(GND_net), 
            .I3(n39016), .O(n663)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_29 (.CI(n39016), .I0(delay_counter[27]), .I1(GND_net), 
            .CO(n39017));
    SB_LUT4 i15231_3_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(timer[22]), 
            .I2(n43085), .I3(GND_net), .O(n28294));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15231_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1117_3_lut (.I0(n941), .I1(n1701), 
            .I2(n1653), .I3(GND_net), .O(n1733));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1117_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1116_3_lut (.I0(n1633), .I1(n1700), 
            .I2(n1653), .I3(GND_net), .O(n1732));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i17_3_lut (.I0(encoder0_position[16]), 
            .I1(n17_adj_4925), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n942));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21396_3_lut (.I0(n942), .I1(n1732), .I2(n1733), .I3(GND_net), 
            .O(n34459));
    defparam i21396_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1696 (.I0(n1723), .I1(n1724), .I2(n1728), .I3(n1726), 
            .O(n47229));
    defparam i1_4_lut_adj_1696.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut (.I0(encoder0_position[0]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n33_adj_5022));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut (.I0(encoder0_position[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n32_adj_5021));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i2_1_lut (.I0(encoder1_position_scaled[1]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_4910));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_DFF encoder0_position_scaled_i22 (.Q(encoder0_position_scaled[22]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[22]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_LUT4 mux_83_i4_4_lut (.I0(encoder1_position_scaled[3]), .I1(displacement[3]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[3]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i4_4_lut.LUT_INIT = 16'h0aca;
    SB_DFF encoder0_position_scaled_i21 (.Q(encoder0_position_scaled[21]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[21]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i20 (.Q(encoder0_position_scaled[20]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[20]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i19 (.Q(encoder0_position_scaled[19]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[19]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i18 (.Q(encoder0_position_scaled[18]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[18]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i17 (.Q(encoder0_position_scaled[17]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[17]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i16 (.Q(encoder0_position_scaled[16]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[16]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i15 (.Q(encoder0_position_scaled[15]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[15]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_CARRY encoder0_position_31__I_0_add_1168_4 (.CI(n39736), .I0(n1732), 
            .I1(GND_net), .CO(n39737));
    SB_LUT4 i1_4_lut_adj_1697 (.I0(n1729), .I1(n34459), .I2(n1730), .I3(n1731), 
            .O(n45047));
    defparam i1_4_lut_adj_1697.LUT_INIT = 16'ha080;
    SB_DFF ID_i0_i0 (.Q(ID[0]), .C(CLK_c), .D(n28225));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFF encoder0_position_scaled_i14 (.Q(encoder0_position_scaled[14]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[14]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i13 (.Q(encoder0_position_scaled[13]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[13]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i12 (.Q(encoder0_position_scaled[12]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[12]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i11 (.Q(encoder0_position_scaled[11]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[11]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i10 (.Q(encoder0_position_scaled[10]), 
           .C(CLK_c), .D(encoder0_position_scaled_23__N_34[10]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i9 (.Q(encoder0_position_scaled[9]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[9]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i8 (.Q(encoder0_position_scaled[8]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[8]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i7 (.Q(encoder0_position_scaled[7]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[7]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i6 (.Q(encoder0_position_scaled[6]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[6]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i5 (.Q(encoder0_position_scaled[5]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[5]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i4 (.Q(encoder0_position_scaled[4]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[4]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i3 (.Q(encoder0_position_scaled[3]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[3]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i2 (.Q(encoder0_position_scaled[2]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[2]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF encoder0_position_scaled_i1 (.Q(encoder0_position_scaled[1]), .C(CLK_c), 
           .D(encoder0_position_scaled_23__N_34[1]));   // verilog/TinyFPGA_B.v(221[10] 225[6])
    SB_DFF pwm_setpoint_i22 (.Q(pwm_setpoint[22]), .C(CLK_c), .D(pwm_setpoint_22__N_11[22]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i21 (.Q(pwm_setpoint[21]), .C(CLK_c), .D(pwm_setpoint_22__N_11[21]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i20 (.Q(pwm_setpoint[20]), .C(CLK_c), .D(pwm_setpoint_22__N_11[20]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i19 (.Q(pwm_setpoint[19]), .C(CLK_c), .D(pwm_setpoint_22__N_11[19]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i18 (.Q(pwm_setpoint[18]), .C(CLK_c), .D(pwm_setpoint_22__N_11[18]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i17 (.Q(pwm_setpoint[17]), .C(CLK_c), .D(pwm_setpoint_22__N_11[17]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i16 (.Q(pwm_setpoint[16]), .C(CLK_c), .D(pwm_setpoint_22__N_11[16]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i15 (.Q(pwm_setpoint[15]), .C(CLK_c), .D(pwm_setpoint_22__N_11[15]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i14 (.Q(pwm_setpoint[14]), .C(CLK_c), .D(pwm_setpoint_22__N_11[14]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i13 (.Q(pwm_setpoint[13]), .C(CLK_c), .D(pwm_setpoint_22__N_11[13]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i12 (.Q(pwm_setpoint[12]), .C(CLK_c), .D(pwm_setpoint_22__N_11[12]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i11 (.Q(pwm_setpoint[11]), .C(CLK_c), .D(pwm_setpoint_22__N_11[11]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i10 (.Q(pwm_setpoint[10]), .C(CLK_c), .D(pwm_setpoint_22__N_11[10]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i9 (.Q(pwm_setpoint[9]), .C(CLK_c), .D(pwm_setpoint_22__N_11[9]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i8 (.Q(pwm_setpoint[8]), .C(CLK_c), .D(pwm_setpoint_22__N_11[8]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i7 (.Q(pwm_setpoint[7]), .C(CLK_c), .D(pwm_setpoint_22__N_11[7]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i6 (.Q(pwm_setpoint[6]), .C(CLK_c), .D(pwm_setpoint_22__N_11[6]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i5 (.Q(pwm_setpoint[5]), .C(CLK_c), .D(pwm_setpoint_22__N_11[5]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i4 (.Q(pwm_setpoint[4]), .C(CLK_c), .D(pwm_setpoint_22__N_11[4]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i3 (.Q(pwm_setpoint[3]), .C(CLK_c), .D(pwm_setpoint_22__N_11[3]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i2 (.Q(pwm_setpoint[2]), .C(CLK_c), .D(pwm_setpoint_22__N_11[2]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_DFF pwm_setpoint_i1 (.Q(pwm_setpoint[1]), .C(CLK_c), .D(pwm_setpoint_22__N_11[1]));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 i1_2_lut_adj_1698 (.I0(n1725), .I1(n1727), .I2(GND_net), .I3(GND_net), 
            .O(n47145));
    defparam i1_2_lut_adj_1698.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1699 (.I0(n45047), .I1(n1721), .I2(n1722), .I3(n47229), 
            .O(n46363));
    defparam i1_4_lut_adj_1699.LUT_INIT = 16'hfffe;
    SB_LUT4 i36026_4_lut (.I0(n1720), .I1(n1719), .I2(n46363), .I3(n47145), 
            .O(n1752));
    defparam i36026_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1111_3_lut (.I0(n1628), .I1(n1695), 
            .I2(n1653), .I3(GND_net), .O(n1727));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1111_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1178_3_lut (.I0(n1727), .I1(n1794), 
            .I2(n1752), .I3(GND_net), .O(n1826));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1178_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1179_3_lut (.I0(n1728), .I1(n1795), 
            .I2(n1752), .I3(GND_net), .O(n1827));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1179_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1177_3_lut (.I0(n1726), .I1(n1793), 
            .I2(n1752), .I3(GND_net), .O(n1825));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1177_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1700 (.I0(n1825), .I1(n1827), .I2(n1828), .I3(n1826), 
            .O(n47287));
    defparam i1_4_lut_adj_1700.LUT_INIT = 16'hfffe;
    SB_LUT4 i21394_3_lut (.I0(n943), .I1(n1832), .I2(n1833), .I3(GND_net), 
            .O(n34457));
    defparam i21394_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_adj_1701 (.I0(n1823), .I1(n1824), .I2(n47287), .I3(GND_net), 
            .O(n47291));
    defparam i1_3_lut_adj_1701.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1702 (.I0(n1829), .I1(n34457), .I2(n1830), .I3(n1831), 
            .O(n45088));
    defparam i1_4_lut_adj_1702.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1703 (.I0(n1821), .I1(n1822), .I2(n45088), .I3(n47291), 
            .O(n47297));
    defparam i1_4_lut_adj_1703.LUT_INIT = 16'hfffe;
    SB_LUT4 i36049_4_lut (.I0(n1819), .I1(n1818), .I2(n1820), .I3(n47297), 
            .O(n1851));
    defparam i36049_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1180_rep_50_3_lut (.I0(n1729), .I1(n1796), 
            .I2(n1752), .I3(GND_net), .O(n1828));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1180_rep_50_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1247_3_lut (.I0(n1828), .I1(n1895), 
            .I2(n1851), .I3(GND_net), .O(n1927));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1247_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15232_3_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(timer[21]), 
            .I2(n43085), .I3(GND_net), .O(n28295));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15232_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_632_4 (.CI(n39632), .I0(n932), 
            .I1(GND_net), .CO(n39633));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut (.I0(encoder0_position[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n31_adj_5020));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut (.I0(encoder0_position[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n30_adj_5019));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut (.I0(encoder0_position[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n29_adj_5018));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_29_28_lut (.I0(GND_net), .I1(delay_counter[26]), .I2(GND_net), 
            .I3(n39015), .O(n664)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_20_lut (.I0(GND_net), .I1(encoder0_position_scaled[18]), 
            .I2(n7_adj_4893), .I3(n39318), .O(displacement_23__N_82[18])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1168_3_lut (.I0(GND_net), .I1(n1733), 
            .I2(VCC_net), .I3(n39735), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i3_1_lut (.I0(encoder1_position_scaled[2]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_4909));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36284_1_lut (.I0(n3138), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51237));
    defparam i36284_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15233_3_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(timer[20]), 
            .I2(n43085), .I3(GND_net), .O(n28296));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15233_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_632_3_lut (.I0(GND_net), .I1(n933), 
            .I2(VCC_net), .I3(n39631), .O(n1000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_20 (.CI(n39318), .I0(encoder0_position_scaled[18]), 
            .I1(n7_adj_4893), .CO(n39319));
    SB_CARRY encoder0_position_31__I_0_add_632_3 (.CI(n39631), .I0(n933), 
            .I1(VCC_net), .CO(n39632));
    SB_CARRY encoder0_position_31__I_0_add_1168_3 (.CI(n39735), .I0(n1733), 
            .I1(VCC_net), .CO(n39736));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_19_lut (.I0(GND_net), .I1(encoder0_position_scaled[17]), 
            .I2(n8_adj_4894), .I3(n39317), .O(displacement_23__N_82[17])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_632_2_lut (.I0(GND_net), .I1(n934), 
            .I2(GND_net), .I3(VCC_net), .O(n1001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_632_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_632_2 (.CI(VCC_net), .I0(n934), 
            .I1(GND_net), .CO(n39631));
    SB_LUT4 encoder0_position_31__I_0_add_1168_2_lut (.I0(GND_net), .I1(n942), 
            .I2(GND_net), .I3(VCC_net), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1168_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1168_2 (.CI(VCC_net), .I0(n942), 
            .I1(GND_net), .CO(n39735));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_19 (.CI(n39317), .I0(encoder0_position_scaled[17]), 
            .I1(n8_adj_4894), .CO(n39318));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_18_lut (.I0(GND_net), .I1(encoder0_position_scaled[16]), 
            .I2(n9_adj_4895), .I3(n39316), .O(displacement_23__N_82[16])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_18 (.CI(n39316), .I0(encoder0_position_scaled[16]), 
            .I1(n9_adj_4895), .CO(n39317));
    SB_CARRY add_29_28 (.CI(n39015), .I0(delay_counter[26]), .I1(GND_net), 
            .CO(n39016));
    SB_LUT4 add_29_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(GND_net), 
            .I3(n38996), .O(n683)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_29_27_lut (.I0(GND_net), .I1(delay_counter[25]), .I2(GND_net), 
            .I3(n39014), .O(n665)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_27 (.CI(n39014), .I0(delay_counter[25]), .I1(GND_net), 
            .CO(n39015));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_17_lut (.I0(GND_net), .I1(encoder0_position_scaled[15]), 
            .I2(n10_adj_4896), .I3(n39315), .O(displacement_23__N_82[15])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_17 (.CI(n39315), .I0(encoder0_position_scaled[15]), 
            .I1(n10_adj_4896), .CO(n39316));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_16_lut (.I0(GND_net), .I1(encoder0_position_scaled[14]), 
            .I2(n11_adj_4897), .I3(n39314), .O(displacement_23__N_82[14])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_16 (.CI(n39314), .I0(encoder0_position_scaled[14]), 
            .I1(n11_adj_4897), .CO(n39315));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_15_lut (.I0(GND_net), .I1(encoder0_position_scaled[13]), 
            .I2(n12_adj_4898), .I3(n39313), .O(displacement_23__N_82[13])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_83_i5_4_lut (.I0(encoder1_position_scaled[4]), .I1(displacement[4]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[4]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i5_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i4_1_lut (.I0(encoder1_position_scaled[3]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_4908));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut (.I0(encoder0_position[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n28_adj_5017));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i5_1_lut (.I0(encoder1_position_scaled[4]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_4907));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15246_3_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(timer[7]), 
            .I2(n43085), .I3(GND_net), .O(n28309));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15246_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut (.I0(encoder0_position[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n27_adj_5016));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15247_3_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(timer[6]), 
            .I2(n43085), .I3(GND_net), .O(n28310));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15247_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut (.I0(encoder0_position[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n26_adj_5015));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut (.I0(encoder0_position[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n25_adj_5014));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut (.I0(encoder0_position[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n24_adj_5013));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_83_i6_4_lut (.I0(encoder1_position_scaled[5]), .I1(displacement[5]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[5]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i6_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut (.I0(encoder0_position[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n23_adj_5012));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut (.I0(encoder0_position[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n22_adj_5011));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut (.I0(encoder0_position[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n21_adj_5010));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15250_3_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(timer[3]), 
            .I2(n43085), .I3(GND_net), .O(n28313));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut (.I0(encoder0_position[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_5009));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut (.I0(encoder0_position[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_5008));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut (.I0(encoder0_position[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_5007));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut (.I0(encoder0_position[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_5006));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_IO NEOPXL_pad (.PACKAGE_PIN(NEOPXL), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(NEOPXL_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam NEOPXL_pad.PIN_TYPE = 6'b011001;
    defparam NEOPXL_pad.PULLUP = 1'b0;
    defparam NEOPXL_pad.NEG_TRIGGER = 1'b0;
    defparam NEOPXL_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO USBPU_pad (.PACKAGE_PIN(USBPU), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(GND_net));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam USBPU_pad.PIN_TYPE = 6'b011001;
    defparam USBPU_pad.PULLUP = 1'b0;
    defparam USBPU_pad.NEG_TRIGGER = 1'b0;
    defparam USBPU_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // /home/letrend/lscc/iCEcube2.2017.08/LSE/userware/unix/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i6_1_lut (.I0(encoder1_position_scaled[5]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n20_adj_4906));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_15 (.CI(n39313), .I0(encoder0_position_scaled[13]), 
            .I1(n12_adj_4898), .CO(n39314));
    SB_LUT4 add_29_26_lut (.I0(GND_net), .I1(delay_counter[24]), .I2(GND_net), 
            .I3(n39013), .O(n666)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_14_lut (.I0(GND_net), .I1(encoder0_position_scaled[12]), 
            .I2(n13_adj_4899), .I3(n39312), .O(displacement_23__N_82[12])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35466_4_lut (.I0(n15_adj_4971), .I1(n13_adj_4970), .I2(n11_adj_4968), 
            .I3(n50283), .O(n50419));
    defparam i35466_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35464_4_lut (.I0(n21_adj_4974), .I1(n19_adj_4973), .I2(n17_adj_4972), 
            .I3(n50419), .O(n50417));
    defparam i35464_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35066_4_lut (.I0(n27_adj_4977), .I1(n25_adj_4976), .I2(n23_adj_4975), 
            .I3(n50417), .O(n50018));
    defparam i35066_4_lut.LUT_INIT = 16'haaab;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_14 (.CI(n39312), .I0(encoder0_position_scaled[12]), 
            .I1(n13_adj_4899), .CO(n39313));
    SB_DFFESR delay_counter_i0_i21 (.Q(delay_counter[21]), .C(CLK_c), .E(n5722), 
            .D(n669), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut (.I0(encoder0_position[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_5005));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut (.I0(encoder0_position[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_5004));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut (.I0(encoder0_position[19]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_5003));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 LessThan_699_i4_4_lut (.I0(pwm_setpoint[0]), .I1(pwm_setpoint[1]), 
            .I2(pwm_counter[1]), .I3(pwm_counter[0]), .O(n4_adj_4962));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i35552_3_lut (.I0(n4_adj_4962), .I1(pwm_setpoint[13]), .I2(n27_adj_4977), 
            .I3(GND_net), .O(n50505));   // verilog/pwm.v(21[8:24])
    defparam i35552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_1940_25_lut (.I0(n50783), .I1(n2_adj_4991), .I2(n1059), 
            .I3(n40325), .O(encoder0_position_scaled_23__N_34[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_25_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_1940_24_lut (.I0(n50798), .I1(n2_adj_4991), .I2(n1158), 
            .I3(n40324), .O(encoder0_position_scaled_23__N_34[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_24_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1940_24 (.CI(n40324), .I0(n2_adj_4991), .I1(n1158), .CO(n40325));
    SB_LUT4 add_1940_23_lut (.I0(n50817), .I1(n2_adj_4991), .I2(n1257), 
            .I3(n40323), .O(encoder0_position_scaled_23__N_34[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1940_23 (.CI(n40323), .I0(n2_adj_4991), .I1(n1257), .CO(n40324));
    SB_LUT4 add_1940_22_lut (.I0(n50832), .I1(n2_adj_4991), .I2(n1356), 
            .I3(n40322), .O(encoder0_position_scaled_23__N_34[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_22_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1940_22 (.CI(n40322), .I0(n2_adj_4991), .I1(n1356), .CO(n40323));
    SB_LUT4 add_1940_21_lut (.I0(n50904), .I1(n2_adj_4991), .I2(n1455), 
            .I3(n40321), .O(encoder0_position_scaled_23__N_34[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_21_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1940_21 (.CI(n40321), .I0(n2_adj_4991), .I1(n1455), .CO(n40322));
    SB_LUT4 add_1940_20_lut (.I0(n50933), .I1(n2_adj_4991), .I2(n1554), 
            .I3(n40320), .O(encoder0_position_scaled_23__N_34[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_20_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1940_20 (.CI(n40320), .I0(n2_adj_4991), .I1(n1554), .CO(n40321));
    SB_LUT4 add_1940_19_lut (.I0(n50955), .I1(n2_adj_4991), .I2(n1653), 
            .I3(n40319), .O(encoder0_position_scaled_23__N_34[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1940_19 (.CI(n40319), .I0(n2_adj_4991), .I1(n1653), .CO(n40320));
    SB_LUT4 add_1940_18_lut (.I0(n50974), .I1(n2_adj_4991), .I2(n1752), 
            .I3(n40318), .O(encoder0_position_scaled_23__N_34[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1940_18 (.CI(n40318), .I0(n2_adj_4991), .I1(n1752), .CO(n40319));
    SB_LUT4 add_1940_17_lut (.I0(n50998), .I1(n2_adj_4991), .I2(n1851), 
            .I3(n40317), .O(encoder0_position_scaled_23__N_34[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_17_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1940_17 (.CI(n40317), .I0(n2_adj_4991), .I1(n1851), .CO(n40318));
    SB_LUT4 mux_83_i7_4_lut (.I0(encoder1_position_scaled[6]), .I1(displacement[6]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[6]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i7_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 add_1940_16_lut (.I0(n51019), .I1(n2_adj_4991), .I2(n1950), 
            .I3(n40316), .O(encoder0_position_scaled_23__N_34[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 LessThan_699_i30_3_lut (.I0(n12_adj_4969), .I1(pwm_setpoint[17]), 
            .I2(n35), .I3(GND_net), .O(n30_adj_4979));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_1940_16 (.CI(n40316), .I0(n2_adj_4991), .I1(n1950), .CO(n40317));
    SB_LUT4 add_1940_15_lut (.I0(n51045), .I1(n2_adj_4991), .I2(n2049), 
            .I3(n40315), .O(encoder0_position_scaled_23__N_34[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i15251_3_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(timer[2]), 
            .I2(n43085), .I3(GND_net), .O(n28314));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15251_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1940_15 (.CI(n40315), .I0(n2_adj_4991), .I1(n2049), .CO(n40316));
    SB_LUT4 add_1940_14_lut (.I0(n51056), .I1(n2_adj_4991), .I2(n2148), 
            .I3(n40314), .O(encoder0_position_scaled_23__N_34[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_14_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1940_14 (.CI(n40314), .I0(n2_adj_4991), .I1(n2148), .CO(n40315));
    SB_LUT4 add_1940_13_lut (.I0(n51302), .I1(n2_adj_4991), .I2(n2247), 
            .I3(n40313), .O(encoder0_position_scaled_23__N_34[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_13_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1940_13 (.CI(n40313), .I0(n2_adj_4991), .I1(n2247), .CO(n40314));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_13_lut (.I0(GND_net), .I1(encoder0_position_scaled[11]), 
            .I2(n14_adj_4900), .I3(n39311), .O(displacement_23__N_82[11])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut (.I0(encoder0_position[20]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_5002));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_1940_12_lut (.I0(n51327), .I1(n2_adj_4991), .I2(n2346), 
            .I3(n40312), .O(encoder0_position_scaled_23__N_34[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_12_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1940_12 (.CI(n40312), .I0(n2_adj_4991), .I1(n2346), .CO(n40313));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_13 (.CI(n39311), .I0(encoder0_position_scaled[11]), 
            .I1(n14_adj_4900), .CO(n39312));
    SB_LUT4 add_1940_11_lut (.I0(n51356), .I1(n2_adj_4991), .I2(n2445), 
            .I3(n40311), .O(encoder0_position_scaled_23__N_34[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1940_11 (.CI(n40311), .I0(n2_adj_4991), .I1(n2445), .CO(n40312));
    SB_LUT4 add_1940_10_lut (.I0(n51390), .I1(n2_adj_4991), .I2(n2544), 
            .I3(n40310), .O(encoder0_position_scaled_23__N_34[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_10_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1940_10 (.CI(n40310), .I0(n2_adj_4991), .I1(n2544), .CO(n40311));
    SB_LUT4 add_1940_9_lut (.I0(n50740), .I1(n2_adj_4991), .I2(n2643), 
            .I3(n40309), .O(encoder0_position_scaled_23__N_34[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_9_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1940_9 (.CI(n40309), .I0(n2_adj_4991), .I1(n2643), .CO(n40310));
    SB_LUT4 add_1940_8_lut (.I0(n51102), .I1(n2_adj_4991), .I2(n2742), 
            .I3(n40308), .O(encoder0_position_scaled_23__N_34[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_12_lut (.I0(GND_net), .I1(encoder0_position_scaled[10]), 
            .I2(n15_adj_4901), .I3(n39310), .O(displacement_23__N_82[10])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1940_8 (.CI(n40308), .I0(n2_adj_4991), .I1(n2742), .CO(n40309));
    SB_LUT4 add_1940_7_lut (.I0(n51137), .I1(n2_adj_4991), .I2(n2841), 
            .I3(n40307), .O(encoder0_position_scaled_23__N_34[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_7_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_12 (.CI(n39310), .I0(encoder0_position_scaled[10]), 
            .I1(n15_adj_4901), .CO(n39311));
    SB_CARRY add_1940_7 (.CI(n40307), .I0(n2_adj_4991), .I1(n2841), .CO(n40308));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i7_1_lut (.I0(encoder1_position_scaled[6]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n19_adj_4905));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_1940_6_lut (.I0(n51169), .I1(n2_adj_4991), .I2(n2940), 
            .I3(n40306), .O(encoder0_position_scaled_23__N_34[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_6_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_11_lut (.I0(GND_net), .I1(encoder0_position_scaled[9]), 
            .I2(n16_adj_4902), .I3(n39309), .O(displacement_23__N_82[9])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_1940_6 (.CI(n40306), .I0(n2_adj_4991), .I1(n2940), .CO(n40307));
    SB_LUT4 add_1940_5_lut (.I0(n51203), .I1(n2_adj_4991), .I2(n3039), 
            .I3(n40305), .O(encoder0_position_scaled_23__N_34[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1940_5 (.CI(n40305), .I0(n2_adj_4991), .I1(n3039), .CO(n40306));
    SB_LUT4 add_1940_4_lut (.I0(n51237), .I1(n2_adj_4991), .I2(n3138), 
            .I3(n40304), .O(encoder0_position_scaled_23__N_34[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_4_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1940_4 (.CI(n40304), .I0(n2_adj_4991), .I1(n3138), .CO(n40305));
    SB_LUT4 add_1940_3_lut (.I0(n51241), .I1(n2_adj_4991), .I2(n3237), 
            .I3(n40303), .O(encoder0_position_scaled_23__N_34[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1940_3 (.CI(n40303), .I0(n2_adj_4991), .I1(n3237), .CO(n40304));
    SB_LUT4 add_1940_2_lut (.I0(n51275), .I1(n2_adj_4991), .I2(n34801), 
            .I3(VCC_net), .O(encoder0_position_scaled_23__N_34[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_1940_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1940_2 (.CI(VCC_net), .I0(n2_adj_4991), .I1(n34801), 
            .CO(n40303));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i8_1_lut (.I0(encoder1_position_scaled[7]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n18_adj_4904));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_11 (.CI(n39309), .I0(encoder0_position_scaled[9]), 
            .I1(n16_adj_4902), .CO(n39310));
    SB_LUT4 encoder0_position_31__I_0_add_2173_33_lut (.I0(n51241), .I1(n3204), 
            .I2(VCC_net), .I3(n40302), .O(n48729)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_2173_32_lut (.I0(GND_net), .I1(n3205), 
            .I2(VCC_net), .I3(n40301), .O(n3272)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_32 (.CI(n40301), .I0(n3205), 
            .I1(VCC_net), .CO(n40302));
    SB_LUT4 encoder0_position_31__I_0_add_2173_31_lut (.I0(GND_net), .I1(n3206), 
            .I2(VCC_net), .I3(n40300), .O(n3273)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_31 (.CI(n40300), .I0(n3206), 
            .I1(VCC_net), .CO(n40301));
    SB_LUT4 encoder0_position_31__I_0_add_2173_30_lut (.I0(GND_net), .I1(n3207), 
            .I2(VCC_net), .I3(n40299), .O(n3274)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_30 (.CI(n40299), .I0(n3207), 
            .I1(VCC_net), .CO(n40300));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut (.I0(encoder0_position[21]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_5001));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_2173_29_lut (.I0(GND_net), .I1(n3208), 
            .I2(VCC_net), .I3(n40298), .O(n3275)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_29 (.CI(n40298), .I0(n3208), 
            .I1(VCC_net), .CO(n40299));
    SB_LUT4 encoder0_position_31__I_0_add_2173_28_lut (.I0(GND_net), .I1(n3209), 
            .I2(VCC_net), .I3(n40297), .O(n3276)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_28 (.CI(n40297), .I0(n3209), 
            .I1(VCC_net), .CO(n40298));
    SB_LUT4 encoder0_position_31__I_0_add_2173_27_lut (.I0(GND_net), .I1(n3210), 
            .I2(VCC_net), .I3(n40296), .O(n3277)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_27 (.CI(n40296), .I0(n3210), 
            .I1(VCC_net), .CO(n40297));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_10_lut (.I0(GND_net), .I1(encoder0_position_scaled[8]), 
            .I2(n17_adj_4903), .I3(n39308), .O(displacement_23__N_82[8])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_10 (.CI(n39308), .I0(encoder0_position_scaled[8]), 
            .I1(n17_adj_4903), .CO(n39309));
    SB_LUT4 encoder0_position_31__I_0_add_2173_26_lut (.I0(GND_net), .I1(n3211), 
            .I2(VCC_net), .I3(n40295), .O(n3278)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut (.I0(encoder0_position[22]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_5000));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_2173_26 (.CI(n40295), .I0(n3211), 
            .I1(VCC_net), .CO(n40296));
    SB_LUT4 encoder0_position_31__I_0_add_2173_25_lut (.I0(GND_net), .I1(n3212), 
            .I2(VCC_net), .I3(n40294), .O(n3279)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_25 (.CI(n40294), .I0(n3212), 
            .I1(VCC_net), .CO(n40295));
    SB_LUT4 encoder0_position_31__I_0_add_2173_24_lut (.I0(GND_net), .I1(n3213), 
            .I2(VCC_net), .I3(n40293), .O(n3280)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_26 (.CI(n39013), .I0(delay_counter[24]), .I1(GND_net), 
            .CO(n39014));
    SB_CARRY encoder0_position_31__I_0_add_2173_24 (.CI(n40293), .I0(n3213), 
            .I1(VCC_net), .CO(n40294));
    SB_LUT4 encoder0_position_31__I_0_add_2173_23_lut (.I0(GND_net), .I1(n3214), 
            .I2(VCC_net), .I3(n40292), .O(n3281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_9_lut (.I0(GND_net), .I1(encoder0_position_scaled[7]), 
            .I2(n18_adj_4904), .I3(n39307), .O(displacement_23__N_82[7])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut (.I0(encoder0_position[23]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4999));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_9 (.CI(n39307), .I0(encoder0_position_scaled[7]), 
            .I1(n18_adj_4904), .CO(n39308));
    SB_CARRY encoder0_position_31__I_0_add_2173_23 (.CI(n40292), .I0(n3214), 
            .I1(VCC_net), .CO(n40293));
    SB_LUT4 encoder0_position_31__I_0_add_2173_22_lut (.I0(GND_net), .I1(n3215), 
            .I2(VCC_net), .I3(n40291), .O(n3282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_22 (.CI(n40291), .I0(n3215), 
            .I1(VCC_net), .CO(n40292));
    SB_LUT4 encoder0_position_31__I_0_add_2173_21_lut (.I0(GND_net), .I1(n3216), 
            .I2(VCC_net), .I3(n40290), .O(n3283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut (.I0(encoder0_position[24]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4998));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_8_lut (.I0(GND_net), .I1(encoder0_position_scaled[6]), 
            .I2(n19_adj_4905), .I3(n39306), .O(displacement_23__N_82[6])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_8 (.CI(n39306), .I0(encoder0_position_scaled[6]), 
            .I1(n19_adj_4905), .CO(n39307));
    SB_CARRY encoder0_position_31__I_0_add_2173_21 (.CI(n40290), .I0(n3216), 
            .I1(VCC_net), .CO(n40291));
    SB_LUT4 encoder0_position_31__I_0_add_2173_20_lut (.I0(GND_net), .I1(n3217), 
            .I2(VCC_net), .I3(n40289), .O(n3284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_20 (.CI(n40289), .I0(n3217), 
            .I1(VCC_net), .CO(n40290));
    SB_LUT4 encoder0_position_31__I_0_add_2173_19_lut (.I0(GND_net), .I1(n3218), 
            .I2(VCC_net), .I3(n40288), .O(n3285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut (.I0(encoder0_position[25]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4997));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut (.I0(encoder0_position[26]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4996));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_2173_19 (.CI(n40288), .I0(n3218), 
            .I1(VCC_net), .CO(n40289));
    SB_LUT4 i15248_3_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(timer[5]), 
            .I2(n43085), .I3(GND_net), .O(n28311));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15248_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_18_lut (.I0(GND_net), .I1(n3219), 
            .I2(VCC_net), .I3(n40287), .O(n3286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_18 (.CI(n40287), .I0(n3219), 
            .I1(VCC_net), .CO(n40288));
    SB_LUT4 add_29_25_lut (.I0(GND_net), .I1(delay_counter[23]), .I2(GND_net), 
            .I3(n39012), .O(n667)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2173_17_lut (.I0(GND_net), .I1(n3220), 
            .I2(VCC_net), .I3(n40286), .O(n3287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_17 (.CI(n40286), .I0(n3220), 
            .I1(VCC_net), .CO(n40287));
    SB_LUT4 encoder0_position_31__I_0_add_2173_16_lut (.I0(GND_net), .I1(n3221), 
            .I2(VCC_net), .I3(n40285), .O(n3288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_16 (.CI(n40285), .I0(n3221), 
            .I1(VCC_net), .CO(n40286));
    SB_LUT4 encoder0_position_31__I_0_add_2173_15_lut (.I0(GND_net), .I1(n3222), 
            .I2(VCC_net), .I3(n40284), .O(n3289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_15 (.CI(n40284), .I0(n3222), 
            .I1(VCC_net), .CO(n40285));
    SB_LUT4 encoder0_position_31__I_0_add_2173_14_lut (.I0(GND_net), .I1(n3223), 
            .I2(VCC_net), .I3(n40283), .O(n3290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_14 (.CI(n40283), .I0(n3223), 
            .I1(VCC_net), .CO(n40284));
    SB_LUT4 encoder0_position_31__I_0_add_2173_13_lut (.I0(GND_net), .I1(n3224), 
            .I2(VCC_net), .I3(n40282), .O(n3291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut (.I0(encoder0_position[27]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n6_adj_4995));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_2173_13 (.CI(n40282), .I0(n3224), 
            .I1(VCC_net), .CO(n40283));
    SB_LUT4 encoder0_position_31__I_0_add_2173_12_lut (.I0(GND_net), .I1(n3225), 
            .I2(VCC_net), .I3(n40281), .O(n3292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_9 (.CI(n38996), .I0(delay_counter[7]), .I1(GND_net), 
            .CO(n38997));
    SB_LUT4 i15252_3_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(timer[1]), 
            .I2(n43085), .I3(GND_net), .O(n28315));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15252_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2173_12 (.CI(n40281), .I0(n3225), 
            .I1(VCC_net), .CO(n40282));
    SB_LUT4 encoder0_position_31__I_0_add_2173_11_lut (.I0(GND_net), .I1(n3226), 
            .I2(VCC_net), .I3(n40280), .O(n3293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_11 (.CI(n40280), .I0(n3226), 
            .I1(VCC_net), .CO(n40281));
    SB_LUT4 encoder0_position_31__I_0_add_2173_10_lut (.I0(GND_net), .I1(n3227), 
            .I2(VCC_net), .I3(n40279), .O(n3294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_10 (.CI(n40279), .I0(n3227), 
            .I1(VCC_net), .CO(n40280));
    SB_LUT4 encoder0_position_31__I_0_add_2173_9_lut (.I0(GND_net), .I1(n3228), 
            .I2(VCC_net), .I3(n40278), .O(n3295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_7_lut (.I0(GND_net), .I1(encoder0_position_scaled[5]), 
            .I2(n20_adj_4906), .I3(n39305), .O(displacement_23__N_82[5])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_9 (.CI(n40278), .I0(n3228), 
            .I1(VCC_net), .CO(n40279));
    SB_LUT4 encoder0_position_31__I_0_add_2173_8_lut (.I0(GND_net), .I1(n3229), 
            .I2(GND_net), .I3(n40277), .O(n3296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_7 (.CI(n39305), .I0(encoder0_position_scaled[5]), 
            .I1(n20_adj_4906), .CO(n39306));
    SB_CARRY encoder0_position_31__I_0_add_2173_8 (.CI(n40277), .I0(n3229), 
            .I1(GND_net), .CO(n40278));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_6_lut (.I0(GND_net), .I1(encoder0_position_scaled[4]), 
            .I2(n21_adj_4907), .I3(n39304), .O(displacement_23__N_82[4])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15234_3_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(timer[19]), 
            .I2(n43085), .I3(GND_net), .O(n28297));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15234_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2173_7_lut (.I0(n3298), .I1(n3230), 
            .I2(GND_net), .I3(n40276), .O(n49734)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_6 (.CI(n39304), .I0(encoder0_position_scaled[4]), 
            .I1(n21_adj_4907), .CO(n39305));
    SB_CARRY encoder0_position_31__I_0_add_2173_7 (.CI(n40276), .I0(n3230), 
            .I1(GND_net), .CO(n40277));
    SB_LUT4 encoder0_position_31__I_0_add_2173_6_lut (.I0(GND_net), .I1(n3231), 
            .I2(VCC_net), .I3(n40275), .O(n3298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_6 (.CI(n40275), .I0(n3231), 
            .I1(VCC_net), .CO(n40276));
    SB_LUT4 encoder0_position_31__I_0_add_2173_5_lut (.I0(GND_net), .I1(n3232), 
            .I2(GND_net), .I3(n40274), .O(n3299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_5 (.CI(n40274), .I0(n3232), 
            .I1(GND_net), .CO(n40275));
    SB_LUT4 encoder0_position_31__I_0_add_2173_4_lut (.I0(GND_net), .I1(n3233), 
            .I2(VCC_net), .I3(n40273), .O(n3300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_4 (.CI(n40273), .I0(n3233), 
            .I1(VCC_net), .CO(n40274));
    SB_LUT4 encoder0_position_31__I_0_add_2173_3_lut (.I0(GND_net), .I1(n957), 
            .I2(GND_net), .I3(n40272), .O(n3301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2173_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut (.I0(encoder0_position[28]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n5_adj_4994));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_83_i8_4_lut (.I0(encoder1_position_scaled[7]), .I1(displacement[7]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[7]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i8_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_5_lut (.I0(GND_net), .I1(encoder0_position_scaled[3]), 
            .I2(n22_adj_4908), .I3(n39303), .O(displacement_23__N_82[3])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2173_3 (.CI(n40272), .I0(n957), 
            .I1(GND_net), .CO(n40273));
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_5 (.CI(n39303), .I0(encoder0_position_scaled[3]), 
            .I1(n22_adj_4908), .CO(n39304));
    SB_CARRY encoder0_position_31__I_0_add_2173_2 (.CI(VCC_net), .I0(n652), 
            .I1(VCC_net), .CO(n40272));
    SB_LUT4 encoder0_position_31__I_0_add_2106_31_lut (.I0(n51237), .I1(n3105), 
            .I2(VCC_net), .I3(n40271), .O(n3204)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_2106_30_lut (.I0(GND_net), .I1(n3106), 
            .I2(VCC_net), .I3(n40270), .O(n3173)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_4_lut (.I0(GND_net), .I1(encoder0_position_scaled[2]), 
            .I2(n23_adj_4909), .I3(n39302), .O(displacement_23__N_82[2])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_30 (.CI(n40270), .I0(n3106), 
            .I1(VCC_net), .CO(n40271));
    SB_LUT4 encoder0_position_31__I_0_add_2106_29_lut (.I0(GND_net), .I1(n3107), 
            .I2(VCC_net), .I3(n40269), .O(n3174)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_4 (.CI(n39302), .I0(encoder0_position_scaled[2]), 
            .I1(n23_adj_4909), .CO(n39303));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i9_1_lut (.I0(encoder1_position_scaled[8]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n17_adj_4903));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_31__I_0_add_2106_29 (.CI(n40269), .I0(n3107), 
            .I1(VCC_net), .CO(n40270));
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_3_lut (.I0(GND_net), .I1(encoder0_position_scaled[1]), 
            .I2(n24_adj_4910), .I3(n39301), .O(displacement_23__N_82[1])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_28_lut (.I0(GND_net), .I1(n3108), 
            .I2(VCC_net), .I3(n40268), .O(n3175)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_28_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i36288_1_lut (.I0(n3237), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51241));
    defparam i36288_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_3 (.CI(n39301), .I0(encoder0_position_scaled[1]), 
            .I1(n24_adj_4910), .CO(n39302));
    SB_CARRY encoder0_position_31__I_0_add_2106_28 (.CI(n40268), .I0(n3108), 
            .I1(VCC_net), .CO(n40269));
    SB_LUT4 encoder0_position_31__I_0_add_2106_27_lut (.I0(GND_net), .I1(n3109), 
            .I2(VCC_net), .I3(n40267), .O(n3176)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_27 (.CI(n40267), .I0(n3109), 
            .I1(VCC_net), .CO(n40268));
    SB_LUT4 encoder0_position_31__I_0_add_2106_26_lut (.I0(GND_net), .I1(n3110), 
            .I2(VCC_net), .I3(n40266), .O(n3177)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_26 (.CI(n40266), .I0(n3110), 
            .I1(VCC_net), .CO(n40267));
    SB_LUT4 encoder0_position_31__I_0_add_2106_25_lut (.I0(GND_net), .I1(n3111), 
            .I2(VCC_net), .I3(n40265), .O(n3178)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_25 (.CI(n40265), .I0(n3111), 
            .I1(VCC_net), .CO(n40266));
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut (.I0(encoder0_position[29]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n4_adj_4993));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i1_3_lut (.I0(encoder0_position[0]), 
            .I1(n33), .I2(encoder0_position[31]), .I3(GND_net), .O(n652));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36322_1_lut (.I0(n34801), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51275));
    defparam i36322_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_add_2_2_lut (.I0(GND_net), .I1(encoder0_position_scaled[0]), 
            .I2(n25_adj_4911), .I3(VCC_net), .O(displacement_23__N_82[0])) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_scaled_23__I_0_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_24_lut (.I0(GND_net), .I1(n3112), 
            .I2(VCC_net), .I3(n40264), .O(n3179)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_24 (.CI(n40264), .I0(n3112), 
            .I1(VCC_net), .CO(n40265));
    SB_LUT4 encoder0_position_31__I_0_add_2106_23_lut (.I0(GND_net), .I1(n3113), 
            .I2(VCC_net), .I3(n40263), .O(n3180)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_scaled_23__I_0_add_2_2 (.CI(VCC_net), .I0(encoder0_position_scaled[0]), 
            .I1(n25_adj_4911), .CO(n39301));
    SB_LUT4 encoder0_position_31__I_0_i2198_3_lut (.I0(n3227), .I1(n3294), 
            .I2(n3237), .I3(GND_net), .O(n17_adj_5028));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2198_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut (.I0(encoder0_position[30]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n3_adj_4992));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2197_3_lut (.I0(n3226), .I1(n3293), 
            .I2(n3237), .I3(GND_net), .O(n19_adj_5029));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2197_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut (.I0(encoder0_position[31]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n2_adj_4991));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_unary_minus_2_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i2192_3_lut (.I0(n3221), .I1(n3288), 
            .I2(n3237), .I3(GND_net), .O(n29_adj_5031));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2192_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2199_3_lut (.I0(n3228), .I1(n3295), 
            .I2(n3237), .I3(GND_net), .O(n15_adj_5027));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2199_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2193_3_lut (.I0(n3222), .I1(n3289), 
            .I2(n3237), .I3(GND_net), .O(n27_adj_5030));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2193_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1704 (.I0(n3220), .I1(n17_adj_5028), .I2(n3287), 
            .I3(n3237), .O(n46959));
    defparam i1_4_lut_adj_1704.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_31__I_0_add_2106_23 (.CI(n40263), .I0(n3113), 
            .I1(VCC_net), .CO(n40264));
    SB_LUT4 i1_4_lut_adj_1705 (.I0(n3225), .I1(n19_adj_5029), .I2(n3292), 
            .I3(n3237), .O(n46961));
    defparam i1_4_lut_adj_1705.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_add_2106_22_lut (.I0(GND_net), .I1(n3114), 
            .I2(VCC_net), .I3(n40262), .O(n3181)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1706 (.I0(n3224), .I1(n27_adj_5030), .I2(n3291), 
            .I3(n3237), .O(n46963));
    defparam i1_4_lut_adj_1706.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_31__I_0_add_2106_22 (.CI(n40262), .I0(n3114), 
            .I1(VCC_net), .CO(n40263));
    SB_LUT4 encoder0_position_31__I_0_add_2106_21_lut (.I0(GND_net), .I1(n3115), 
            .I2(VCC_net), .I3(n40261), .O(n3182)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_25 (.CI(n39012), .I0(delay_counter[23]), .I1(GND_net), 
            .CO(n39013));
    SB_CARRY encoder0_position_31__I_0_add_2106_21 (.CI(n40261), .I0(n3115), 
            .I1(VCC_net), .CO(n40262));
    SB_LUT4 add_673_24_lut (.I0(duty[22]), .I1(n51409), .I2(n3), .I3(n39300), 
            .O(pwm_setpoint_22__N_11[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_24_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_2106_20_lut (.I0(GND_net), .I1(n3116), 
            .I2(VCC_net), .I3(n40260), .O(n3183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_673_23_lut (.I0(duty[21]), .I1(n51409), .I2(n4), .I3(n39299), 
            .O(pwm_setpoint_22__N_11[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_23_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_2106_20 (.CI(n40260), .I0(n3116), 
            .I1(VCC_net), .CO(n40261));
    SB_LUT4 i1_4_lut_adj_1707 (.I0(n3223), .I1(n15_adj_5027), .I2(n3290), 
            .I3(n3237), .O(n46967));
    defparam i1_4_lut_adj_1707.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_add_2106_19_lut (.I0(GND_net), .I1(n3117), 
            .I2(VCC_net), .I3(n40259), .O(n3184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2190_3_lut (.I0(n3219), .I1(n3286), 
            .I2(n3237), .I3(GND_net), .O(n33_adj_5032));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2190_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1708 (.I0(n3229), .I1(n29_adj_5031), .I2(n3296), 
            .I3(n3237), .O(n46965));
    defparam i1_4_lut_adj_1708.LUT_INIT = 16'heefc;
    SB_CARRY encoder0_position_31__I_0_add_2106_19 (.CI(n40259), .I0(n3117), 
            .I1(VCC_net), .CO(n40260));
    SB_LUT4 i1_4_lut_adj_1709 (.I0(n3218), .I1(n33_adj_5032), .I2(n3285), 
            .I3(n3237), .O(n46969));
    defparam i1_4_lut_adj_1709.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_add_2106_18_lut (.I0(GND_net), .I1(n3118), 
            .I2(VCC_net), .I3(n40258), .O(n3185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_18 (.CI(n40258), .I0(n3118), 
            .I1(VCC_net), .CO(n40259));
    SB_LUT4 encoder0_position_31__I_0_add_2106_17_lut (.I0(GND_net), .I1(n3119), 
            .I2(VCC_net), .I3(n40257), .O(n3186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_17 (.CI(n40257), .I0(n3119), 
            .I1(VCC_net), .CO(n40258));
    SB_LUT4 encoder0_position_31__I_0_add_2106_16_lut (.I0(GND_net), .I1(n3120), 
            .I2(VCC_net), .I3(n40256), .O(n3187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_16 (.CI(n40256), .I0(n3120), 
            .I1(VCC_net), .CO(n40257));
    SB_LUT4 encoder0_position_31__I_0_i2188_3_lut (.I0(n3217), .I1(n3284), 
            .I2(n3237), .I3(GND_net), .O(n37));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2188_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1710 (.I0(n46967), .I1(n46963), .I2(n46961), 
            .I3(n46959), .O(n46977));
    defparam i1_4_lut_adj_1710.LUT_INIT = 16'hfffe;
    SB_CARRY add_673_23 (.CI(n39299), .I0(n51409), .I1(n4), .CO(n39300));
    SB_LUT4 i21333_4_lut (.I0(n652), .I1(n957), .I2(n3301), .I3(n3237), 
            .O(n34393));
    defparam i21333_4_lut.LUT_INIT = 16'heefa;
    SB_LUT4 i21518_4_lut (.I0(n34393), .I1(n3233), .I2(n3300), .I3(n3237), 
            .O(n34583));
    defparam i21518_4_lut.LUT_INIT = 16'h88a0;
    SB_LUT4 add_29_24_lut (.I0(GND_net), .I1(delay_counter[22]), .I2(GND_net), 
            .I3(n39011), .O(n668)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_673_22_lut (.I0(duty[20]), .I1(n51409), .I2(n5), .I3(n39298), 
            .O(pwm_setpoint_22__N_11[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_22_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 i1_4_lut_adj_1711 (.I0(n46977), .I1(n37), .I2(n46969), .I3(n46965), 
            .O(n46981));
    defparam i1_4_lut_adj_1711.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n3231), .I1(n49734), .I2(n3237), .I3(n3230), 
            .O(n5_adj_5042));
    defparam i16_4_lut.LUT_INIT = 16'hac0c;
    SB_CARRY add_29_24 (.CI(n39011), .I0(delay_counter[22]), .I1(GND_net), 
            .CO(n39012));
    SB_LUT4 add_29_23_lut (.I0(GND_net), .I1(delay_counter[21]), .I2(GND_net), 
            .I3(n39010), .O(n669)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1712 (.I0(n3216), .I1(n46981), .I2(n3283), .I3(n3237), 
            .O(n46983));
    defparam i1_4_lut_adj_1712.LUT_INIT = 16'heefc;
    SB_CARRY add_29_23 (.CI(n39010), .I0(delay_counter[21]), .I1(GND_net), 
            .CO(n39011));
    SB_LUT4 encoder0_position_31__I_0_add_2106_15_lut (.I0(GND_net), .I1(n3121), 
            .I2(VCC_net), .I3(n40255), .O(n3188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_15 (.CI(n40255), .I0(n3121), 
            .I1(VCC_net), .CO(n40256));
    SB_LUT4 encoder0_position_31__I_0_add_2106_14_lut (.I0(GND_net), .I1(n3122), 
            .I2(VCC_net), .I3(n40254), .O(n3189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_14 (.CI(n40254), .I0(n3122), 
            .I1(VCC_net), .CO(n40255));
    SB_LUT4 i21625_4_lut (.I0(n34583), .I1(n3232), .I2(n3299), .I3(n3237), 
            .O(n34693));
    defparam i21625_4_lut.LUT_INIT = 16'heefa;
    SB_LUT4 encoder0_position_31__I_0_add_2106_13_lut (.I0(GND_net), .I1(n3123), 
            .I2(VCC_net), .I3(n40253), .O(n3190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_13 (.CI(n40253), .I0(n3123), 
            .I1(VCC_net), .CO(n40254));
    SB_LUT4 encoder0_position_31__I_0_i2186_3_lut (.I0(n3215), .I1(n3282), 
            .I2(n3237), .I3(GND_net), .O(n41));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2186_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1713 (.I0(n41), .I1(n34693), .I2(n46983), .I3(n5_adj_5042), 
            .O(n46987));
    defparam i1_4_lut_adj_1713.LUT_INIT = 16'hfefa;
    SB_LUT4 i1_4_lut_adj_1714 (.I0(n3214), .I1(n46987), .I2(n3281), .I3(n3237), 
            .O(n46989));
    defparam i1_4_lut_adj_1714.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1715 (.I0(n3213), .I1(n46989), .I2(n3280), .I3(n3237), 
            .O(n46991));
    defparam i1_4_lut_adj_1715.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1716 (.I0(n3212), .I1(n46991), .I2(n3279), .I3(n3237), 
            .O(n46993));
    defparam i1_4_lut_adj_1716.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1717 (.I0(n3211), .I1(n46993), .I2(n3278), .I3(n3237), 
            .O(n46995));
    defparam i1_4_lut_adj_1717.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1718 (.I0(n3210), .I1(n46995), .I2(n3277), .I3(n3237), 
            .O(n46997));
    defparam i1_4_lut_adj_1718.LUT_INIT = 16'heefc;
    SB_LUT4 i1_4_lut_adj_1719 (.I0(n3209), .I1(n46997), .I2(n3276), .I3(n3237), 
            .O(n46999));
    defparam i1_4_lut_adj_1719.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_add_2106_12_lut (.I0(GND_net), .I1(n3124), 
            .I2(VCC_net), .I3(n40252), .O(n3191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_12 (.CI(n40252), .I0(n3124), 
            .I1(VCC_net), .CO(n40253));
    SB_LUT4 encoder0_position_31__I_0_add_2106_11_lut (.I0(GND_net), .I1(n3125), 
            .I2(VCC_net), .I3(n40251), .O(n3192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_11 (.CI(n40251), .I0(n3125), 
            .I1(VCC_net), .CO(n40252));
    SB_LUT4 i1_4_lut_adj_1720 (.I0(n3208), .I1(n46999), .I2(n3275), .I3(n3237), 
            .O(n47001));
    defparam i1_4_lut_adj_1720.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_add_2106_10_lut (.I0(GND_net), .I1(n3126), 
            .I2(VCC_net), .I3(n40250), .O(n3193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1721 (.I0(n3207), .I1(n47001), .I2(n3274), .I3(n3237), 
            .O(n47003));
    defparam i1_4_lut_adj_1721.LUT_INIT = 16'heefc;
    SB_LUT4 encoder0_position_31__I_0_i2177_3_lut (.I0(n3206), .I1(n3273), 
            .I2(n3237), .I3(GND_net), .O(n59));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2177_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_10 (.CI(n40250), .I0(n3126), 
            .I1(VCC_net), .CO(n40251));
    SB_LUT4 encoder0_position_31__I_0_i2176_3_lut (.I0(n3205), .I1(n3272), 
            .I2(n3237), .I3(GND_net), .O(n61_adj_5033));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36325_4_lut (.I0(n61_adj_5033), .I1(n48729), .I2(n59), .I3(n47003), 
            .O(n34801));
    defparam i36325_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i2110_3_lut (.I0(n3107), .I1(n3174), 
            .I2(n3138), .I3(GND_net), .O(n3206));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2109_3_lut (.I0(n3106), .I1(n3173), 
            .I2(n3138), .I3(GND_net), .O(n3205));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_29_22_lut (.I0(GND_net), .I1(delay_counter[20]), .I2(GND_net), 
            .I3(n39009), .O(n670)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2118_3_lut (.I0(n3115), .I1(n3182), 
            .I2(n3138), .I3(GND_net), .O(n3214));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2118_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_9_lut (.I0(GND_net), .I1(n3127), 
            .I2(VCC_net), .I3(n40249), .O(n3194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_9 (.CI(n40249), .I0(n3127), 
            .I1(VCC_net), .CO(n40250));
    SB_LUT4 encoder0_position_31__I_0_add_2106_8_lut (.I0(GND_net), .I1(n3128), 
            .I2(VCC_net), .I3(n40248), .O(n3195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_8 (.CI(n40248), .I0(n3128), 
            .I1(VCC_net), .CO(n40249));
    SB_LUT4 encoder0_position_31__I_0_i2117_3_lut (.I0(n3114), .I1(n3181), 
            .I2(n3138), .I3(GND_net), .O(n3213));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2117_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_673_22 (.CI(n39298), .I0(n51409), .I1(n5), .CO(n39299));
    SB_LUT4 encoder0_position_31__I_0_i2113_3_lut (.I0(n3110), .I1(n3177), 
            .I2(n3138), .I3(GND_net), .O(n3209));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_7_lut (.I0(GND_net), .I1(n3129), 
            .I2(GND_net), .I3(n40247), .O(n3196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2112_3_lut (.I0(n3109), .I1(n3176), 
            .I2(n3138), .I3(GND_net), .O(n3208));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_673_21_lut (.I0(duty[19]), .I1(n51409), .I2(n6), .I3(n39297), 
            .O(pwm_setpoint_22__N_11[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_21_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i2111_3_lut (.I0(n3108), .I1(n3175), 
            .I2(n3138), .I3(GND_net), .O(n3207));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2111_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_2106_7 (.CI(n40247), .I0(n3129), 
            .I1(GND_net), .CO(n40248));
    SB_CARRY add_29_22 (.CI(n39009), .I0(delay_counter[20]), .I1(GND_net), 
            .CO(n39010));
    SB_LUT4 encoder0_position_31__I_0_add_2106_6_lut (.I0(GND_net), .I1(n3130), 
            .I2(GND_net), .I3(n40246), .O(n3197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_6 (.CI(n40246), .I0(n3130), 
            .I1(GND_net), .CO(n40247));
    SB_LUT4 encoder0_position_31__I_0_add_2106_5_lut (.I0(GND_net), .I1(n3131), 
            .I2(VCC_net), .I3(n40245), .O(n3198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15235_3_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(timer[18]), 
            .I2(n43085), .I3(GND_net), .O(n28298));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15235_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36045_1_lut (.I0(n1851), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50998));
    defparam i36045_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i15_3_lut (.I0(encoder0_position[14]), 
            .I1(n19_adj_4923), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n944));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_673_21 (.CI(n39297), .I0(n51409), .I1(n6), .CO(n39298));
    SB_CARRY encoder0_position_31__I_0_add_2106_5 (.CI(n40245), .I0(n3131), 
            .I1(VCC_net), .CO(n40246));
    SB_LUT4 encoder0_position_31__I_0_add_2106_4_lut (.I0(GND_net), .I1(n3132), 
            .I2(GND_net), .I3(n40244), .O(n3199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_4 (.CI(n40244), .I0(n3132), 
            .I1(GND_net), .CO(n40245));
    SB_LUT4 add_29_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(GND_net), 
            .I3(n38995), .O(n684)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2106_3_lut (.I0(GND_net), .I1(n3133), 
            .I2(VCC_net), .I3(n40243), .O(n3200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_3 (.CI(n40243), .I0(n3133), 
            .I1(VCC_net), .CO(n40244));
    SB_LUT4 encoder0_position_31__I_0_i2116_3_lut (.I0(n3113), .I1(n3180), 
            .I2(n3138), .I3(GND_net), .O(n3212));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2116_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2115_3_lut (.I0(n3112), .I1(n3179), 
            .I2(n3138), .I3(GND_net), .O(n3211));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2114_3_lut (.I0(n3111), .I1(n3178), 
            .I2(n3138), .I3(GND_net), .O(n3210));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2106_2_lut (.I0(GND_net), .I1(n956), 
            .I2(GND_net), .I3(VCC_net), .O(n3201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2106_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2106_2 (.CI(VCC_net), .I0(n956), 
            .I1(GND_net), .CO(n40243));
    SB_LUT4 encoder0_position_31__I_0_i2121_3_lut (.I0(n3118), .I1(n3185), 
            .I2(n3138), .I3(GND_net), .O(n3217));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2121_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2120_3_lut (.I0(n3117), .I1(n3184), 
            .I2(n3138), .I3(GND_net), .O(n3216));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2120_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_30_lut (.I0(n51203), .I1(n3006), 
            .I2(VCC_net), .I3(n40242), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_i1046_3_lut (.I0(n1531), .I1(n1598), 
            .I2(n1554), .I3(GND_net), .O(n1630));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2119_3_lut (.I0(n3116), .I1(n3183), 
            .I2(n3138), .I3(GND_net), .O(n3215));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2119_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2127_3_lut (.I0(n3124), .I1(n3191), 
            .I2(n3138), .I3(GND_net), .O(n3223));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2127_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15236_3_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(timer[17]), 
            .I2(n43085), .I3(GND_net), .O(n28299));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15236_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2132_3_lut (.I0(n3129), .I1(n3196), 
            .I2(n3138), .I3(GND_net), .O(n3228));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2132_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2124_3_lut (.I0(n3121), .I1(n3188), 
            .I2(n3138), .I3(GND_net), .O(n3220));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2124_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2130_3_lut (.I0(n3127), .I1(n3194), 
            .I2(n3138), .I3(GND_net), .O(n3226));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2130_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2123_3_lut (.I0(n3120), .I1(n3187), 
            .I2(n3138), .I3(GND_net), .O(n3219));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2123_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2128_3_lut (.I0(n3125), .I1(n3192), 
            .I2(n3138), .I3(GND_net), .O(n3224));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2128_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_29_lut (.I0(GND_net), .I1(n3007), 
            .I2(VCC_net), .I3(n40241), .O(n3074)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_29 (.CI(n40241), .I0(n3007), 
            .I1(VCC_net), .CO(n40242));
    SB_LUT4 encoder0_position_31__I_0_add_2039_28_lut (.I0(GND_net), .I1(n3008), 
            .I2(VCC_net), .I3(n40240), .O(n3075)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_28 (.CI(n40240), .I0(n3008), 
            .I1(VCC_net), .CO(n40241));
    SB_LUT4 add_673_20_lut (.I0(duty[18]), .I1(n51409), .I2(n7_adj_4886), 
            .I3(n39296), .O(pwm_setpoint_22__N_11[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_20_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_1101_16_lut (.I0(n50955), .I1(n1620), 
            .I2(VCC_net), .I3(n39724), .O(n1719)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_i2129_3_lut (.I0(n3126), .I1(n3193), 
            .I2(n3138), .I3(GND_net), .O(n3225));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2129_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_29_21_lut (.I0(GND_net), .I1(delay_counter[19]), .I2(GND_net), 
            .I3(n39008), .O(n671)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_2039_27_lut (.I0(GND_net), .I1(n3009), 
            .I2(VCC_net), .I3(n40239), .O(n3076)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2125_3_lut (.I0(n3122), .I1(n3189), 
            .I2(n3138), .I3(GND_net), .O(n3221));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2125_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_673_20 (.CI(n39296), .I0(n51409), .I1(n7_adj_4886), .CO(n39297));
    SB_CARRY encoder0_position_31__I_0_add_2039_27 (.CI(n40239), .I0(n3009), 
            .I1(VCC_net), .CO(n40240));
    SB_LUT4 encoder0_position_31__I_0_add_2039_26_lut (.I0(GND_net), .I1(n3010), 
            .I2(VCC_net), .I3(n40238), .O(n3077)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_26 (.CI(n40238), .I0(n3010), 
            .I1(VCC_net), .CO(n40239));
    SB_LUT4 encoder0_position_31__I_0_add_2039_25_lut (.I0(GND_net), .I1(n3011), 
            .I2(VCC_net), .I3(n40237), .O(n3078)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_673_19_lut (.I0(duty[17]), .I1(n51409), .I2(n8), .I3(n39295), 
            .O(pwm_setpoint_22__N_11[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_19_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_2039_25 (.CI(n40237), .I0(n3011), 
            .I1(VCC_net), .CO(n40238));
    SB_CARRY add_673_19 (.CI(n39295), .I0(n51409), .I1(n8), .CO(n39296));
    SB_LUT4 encoder0_position_31__I_0_add_1101_15_lut (.I0(GND_net), .I1(n1621), 
            .I2(VCC_net), .I3(n39723), .O(n1688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15237_3_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(timer[16]), 
            .I2(n43085), .I3(GND_net), .O(n28300));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15237_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_24_lut (.I0(GND_net), .I1(n3012), 
            .I2(VCC_net), .I3(n40236), .O(n3079)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_673_18_lut (.I0(duty[16]), .I1(n51409), .I2(n9), .I3(n39294), 
            .O(pwm_setpoint_22__N_11[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_18_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_2039_24 (.CI(n40236), .I0(n3012), 
            .I1(VCC_net), .CO(n40237));
    SB_LUT4 encoder0_position_31__I_0_add_2039_23_lut (.I0(GND_net), .I1(n3013), 
            .I2(VCC_net), .I3(n40235), .O(n3080)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_23 (.CI(n40235), .I0(n3013), 
            .I1(VCC_net), .CO(n40236));
    SB_DFFESR delay_counter_i0_i20 (.Q(delay_counter[20]), .C(CLK_c), .E(n5722), 
            .D(n670), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_add_2039_22_lut (.I0(GND_net), .I1(n3014), 
            .I2(VCC_net), .I3(n40234), .O(n3081)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_15 (.CI(n39723), .I0(n1621), 
            .I1(VCC_net), .CO(n39724));
    SB_LUT4 encoder0_position_31__I_0_i2137_3_lut (.I0(n956), .I1(n3201), 
            .I2(n3138), .I3(GND_net), .O(n3233));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2137_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1101_14_lut (.I0(GND_net), .I1(n1622), 
            .I2(VCC_net), .I3(n39722), .O(n1689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_22 (.CI(n40234), .I0(n3014), 
            .I1(VCC_net), .CO(n40235));
    SB_LUT4 encoder0_position_31__I_0_add_2039_21_lut (.I0(GND_net), .I1(n3015), 
            .I2(VCC_net), .I3(n40233), .O(n3082)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_21 (.CI(n40233), .I0(n3015), 
            .I1(VCC_net), .CO(n40234));
    SB_LUT4 encoder0_position_31__I_0_add_2039_20_lut (.I0(GND_net), .I1(n3016), 
            .I2(VCC_net), .I3(n40232), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_20 (.CI(n40232), .I0(n3016), 
            .I1(VCC_net), .CO(n40233));
    SB_LUT4 encoder0_position_31__I_0_add_2039_19_lut (.I0(GND_net), .I1(n3017), 
            .I2(VCC_net), .I3(n40231), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_19 (.CI(n40231), .I0(n3017), 
            .I1(VCC_net), .CO(n40232));
    SB_LUT4 encoder0_position_31__I_0_add_2039_18_lut (.I0(GND_net), .I1(n3018), 
            .I2(VCC_net), .I3(n40230), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_18 (.CI(n40230), .I0(n3018), 
            .I1(VCC_net), .CO(n40231));
    SB_LUT4 encoder0_position_31__I_0_add_2039_17_lut (.I0(GND_net), .I1(n3019), 
            .I2(VCC_net), .I3(n40229), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_14 (.CI(n39722), .I0(n1622), 
            .I1(VCC_net), .CO(n39723));
    SB_LUT4 encoder0_position_31__I_0_add_1101_13_lut (.I0(GND_net), .I1(n1623), 
            .I2(VCC_net), .I3(n39721), .O(n1690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2136_3_lut (.I0(n3133), .I1(n3200), 
            .I2(n3138), .I3(GND_net), .O(n3232));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2136_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1101_13 (.CI(n39721), .I0(n1623), 
            .I1(VCC_net), .CO(n39722));
    SB_LUT4 encoder0_position_31__I_0_add_1101_12_lut (.I0(GND_net), .I1(n1624), 
            .I2(VCC_net), .I3(n39720), .O(n1691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_673_18 (.CI(n39294), .I0(n51409), .I1(n9), .CO(n39295));
    SB_CARRY encoder0_position_31__I_0_add_1101_12 (.CI(n39720), .I0(n1624), 
            .I1(VCC_net), .CO(n39721));
    SB_LUT4 add_673_17_lut (.I0(duty[15]), .I1(n51409), .I2(n10), .I3(n39293), 
            .O(pwm_setpoint_22__N_11[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_17_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_1101_11_lut (.I0(GND_net), .I1(n1625), 
            .I2(VCC_net), .I3(n39719), .O(n1692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_673_17 (.CI(n39293), .I0(n51409), .I1(n10), .CO(n39294));
    SB_CARRY encoder0_position_31__I_0_add_1101_11 (.CI(n39719), .I0(n1625), 
            .I1(VCC_net), .CO(n39720));
    SB_CARRY encoder0_position_31__I_0_add_2039_17 (.CI(n40229), .I0(n3019), 
            .I1(VCC_net), .CO(n40230));
    SB_LUT4 encoder0_position_31__I_0_add_2039_16_lut (.I0(GND_net), .I1(n3020), 
            .I2(VCC_net), .I3(n40228), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_16 (.CI(n40228), .I0(n3020), 
            .I1(VCC_net), .CO(n40229));
    SB_LUT4 add_673_16_lut (.I0(duty[14]), .I1(n51409), .I2(n11), .I3(n39292), 
            .O(pwm_setpoint_22__N_11[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_16_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_2039_15_lut (.I0(GND_net), .I1(n3021), 
            .I2(VCC_net), .I3(n40227), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i2_3_lut (.I0(encoder0_position[1]), 
            .I1(n32), .I2(encoder0_position[31]), .I3(GND_net), .O(n957));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_2039_15 (.CI(n40227), .I0(n3021), 
            .I1(VCC_net), .CO(n40228));
    SB_LUT4 encoder0_position_31__I_0_add_2039_14_lut (.I0(GND_net), .I1(n3022), 
            .I2(VCC_net), .I3(n40226), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2135_3_lut (.I0(n3132), .I1(n3199), 
            .I2(n3138), .I3(GND_net), .O(n3231));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2135_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2134_3_lut (.I0(n3131), .I1(n3198), 
            .I2(n3138), .I3(GND_net), .O(n3230));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2134_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2133_3_lut (.I0(n3130), .I1(n3197), 
            .I2(n3138), .I3(GND_net), .O(n3229));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2133_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2122_3_lut (.I0(n3119), .I1(n3186), 
            .I2(n3138), .I3(GND_net), .O(n3218));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2122_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2126_3_lut (.I0(n3123), .I1(n3190), 
            .I2(n3138), .I3(GND_net), .O(n3222));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2126_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2131_3_lut (.I0(n3128), .I1(n3195), 
            .I2(n3138), .I3(GND_net), .O(n3227));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2131_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21526_3_lut (.I0(n957), .I1(n3232), .I2(n3233), .I3(GND_net), 
            .O(n34591));
    defparam i21526_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_31__I_0_i1253_3_lut (.I0(n943), .I1(n1901), 
            .I2(n1851), .I3(GND_net), .O(n1933));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1253_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1722 (.I0(n3221), .I1(n3225), .I2(n3224), .I3(n3219), 
            .O(n47547));
    defparam i1_4_lut_adj_1722.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1723 (.I0(n3227), .I1(n3222), .I2(GND_net), .I3(GND_net), 
            .O(n47537));
    defparam i1_2_lut_adj_1723.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1724 (.I0(n3226), .I1(n3220), .I2(n3228), .I3(n3223), 
            .O(n47549));
    defparam i1_4_lut_adj_1724.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_2039_14 (.CI(n40226), .I0(n3022), 
            .I1(VCC_net), .CO(n40227));
    SB_LUT4 encoder0_position_31__I_0_add_2039_13_lut (.I0(GND_net), .I1(n3023), 
            .I2(VCC_net), .I3(n40225), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_13 (.CI(n40225), .I0(n3023), 
            .I1(VCC_net), .CO(n40226));
    SB_LUT4 encoder0_position_31__I_0_add_2039_12_lut (.I0(GND_net), .I1(n3024), 
            .I2(VCC_net), .I3(n40224), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_673_16 (.CI(n39292), .I0(n51409), .I1(n11), .CO(n39293));
    SB_CARRY encoder0_position_31__I_0_add_2039_12 (.CI(n40224), .I0(n3024), 
            .I1(VCC_net), .CO(n40225));
    SB_LUT4 encoder0_position_31__I_0_add_2039_11_lut (.I0(GND_net), .I1(n3025), 
            .I2(VCC_net), .I3(n40223), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1101_10_lut (.I0(GND_net), .I1(n1626), 
            .I2(VCC_net), .I3(n39718), .O(n1693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_10 (.CI(n39718), .I0(n1626), 
            .I1(VCC_net), .CO(n39719));
    SB_LUT4 encoder0_position_31__I_0_add_1101_9_lut (.I0(GND_net), .I1(n1627), 
            .I2(VCC_net), .I3(n39717), .O(n1694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_11 (.CI(n40223), .I0(n3025), 
            .I1(VCC_net), .CO(n40224));
    SB_LUT4 encoder0_position_31__I_0_add_2039_10_lut (.I0(GND_net), .I1(n3026), 
            .I2(VCC_net), .I3(n40222), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_10 (.CI(n40222), .I0(n3026), 
            .I1(VCC_net), .CO(n40223));
    SB_LUT4 encoder0_position_31__I_0_add_2039_9_lut (.I0(GND_net), .I1(n3027), 
            .I2(VCC_net), .I3(n40221), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1725 (.I0(n47549), .I1(n47537), .I2(n47547), 
            .I3(n3218), .O(n47553));
    defparam i1_4_lut_adj_1725.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_2039_9 (.CI(n40221), .I0(n3027), 
            .I1(VCC_net), .CO(n40222));
    SB_LUT4 i1_4_lut_adj_1726 (.I0(n3229), .I1(n34591), .I2(n3230), .I3(n3231), 
            .O(n45178));
    defparam i1_4_lut_adj_1726.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1727 (.I0(n3215), .I1(n3216), .I2(n47553), .I3(n3217), 
            .O(n47559));
    defparam i1_4_lut_adj_1727.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1728 (.I0(n3213), .I1(n3214), .I2(n47559), .I3(n45178), 
            .O(n47565));
    defparam i1_4_lut_adj_1728.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1729 (.I0(n3210), .I1(n3211), .I2(n3212), .I3(n47565), 
            .O(n47571));
    defparam i1_4_lut_adj_1729.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1730 (.I0(n3207), .I1(n3208), .I2(n3209), .I3(n47571), 
            .O(n47577));
    defparam i1_4_lut_adj_1730.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1101_9 (.CI(n39717), .I0(n1627), 
            .I1(VCC_net), .CO(n39718));
    SB_LUT4 RX_I_0_1_lut (.I0(RX_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(RX_N_10));   // verilog/TinyFPGA_B.v(146[10:13])
    defparam RX_I_0_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36321_4_lut (.I0(n3205), .I1(n3204), .I2(n3206), .I3(n47577), 
            .O(n3237));
    defparam i36321_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_2039_8_lut (.I0(GND_net), .I1(n3028), 
            .I2(VCC_net), .I3(n40220), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_8 (.CI(n40220), .I0(n3028), 
            .I1(VCC_net), .CO(n40221));
    SB_LUT4 mux_83_i9_4_lut (.I0(encoder1_position_scaled[8]), .I1(displacement[8]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[8]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i9_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_add_2039_7_lut (.I0(GND_net), .I1(n3029), 
            .I2(GND_net), .I3(n40219), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_7 (.CI(n40219), .I0(n3029), 
            .I1(GND_net), .CO(n40220));
    SB_LUT4 encoder0_position_31__I_0_add_2039_6_lut (.I0(GND_net), .I1(n3030), 
            .I2(GND_net), .I3(n40218), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_6 (.CI(n40218), .I0(n3030), 
            .I1(GND_net), .CO(n40219));
    SB_LUT4 encoder0_position_31__I_0_add_1101_8_lut (.I0(GND_net), .I1(n1628), 
            .I2(VCC_net), .I3(n39716), .O(n1695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_21 (.CI(n39008), .I0(delay_counter[19]), .I1(GND_net), 
            .CO(n39009));
    SB_LUT4 encoder0_position_31__I_0_add_2039_5_lut (.I0(GND_net), .I1(n3031), 
            .I2(VCC_net), .I3(n40217), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_8 (.CI(n39716), .I0(n1628), 
            .I1(VCC_net), .CO(n39717));
    SB_LUT4 encoder0_position_31__I_0_i2043_3_lut (.I0(n3008), .I1(n3075), 
            .I2(n3039), .I3(GND_net), .O(n3107));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2043_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2042_3_lut (.I0(n3007), .I1(n3074), 
            .I2(n3039), .I3(GND_net), .O(n3106));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2046_3_lut (.I0(n3011), .I1(n3078), 
            .I2(n3039), .I3(GND_net), .O(n3110));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2046_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2045_3_lut (.I0(n3010), .I1(n3077), 
            .I2(n3039), .I3(GND_net), .O(n3109));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2044_3_lut (.I0(n3009), .I1(n3076), 
            .I2(n3039), .I3(GND_net), .O(n3108));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1101_7_lut (.I0(GND_net), .I1(n1629), 
            .I2(GND_net), .I3(n39715), .O(n1696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2049_3_lut (.I0(n3014), .I1(n3081), 
            .I2(n3039), .I3(GND_net), .O(n3113));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2049_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2048_3_lut (.I0(n3013), .I1(n3080), 
            .I2(n3039), .I3(GND_net), .O(n3112));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2048_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2047_3_lut (.I0(n3012), .I1(n3079), 
            .I2(n3039), .I3(GND_net), .O(n3111));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2047_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2051_3_lut (.I0(n3016), .I1(n3083), 
            .I2(n3039), .I3(GND_net), .O(n3115));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2051_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2050_3_lut (.I0(n3015), .I1(n3082), 
            .I2(n3039), .I3(GND_net), .O(n3114));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2050_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2067_3_lut (.I0(n3032), .I1(n3099), 
            .I2(n3039), .I3(GND_net), .O(n3131));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2067_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2066_3_lut (.I0(n3031), .I1(n3098), 
            .I2(n3039), .I3(GND_net), .O(n3130));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2066_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2065_3_lut (.I0(n3030), .I1(n3097), 
            .I2(n3039), .I3(GND_net), .O(n3129));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2065_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2053_3_lut (.I0(n3018), .I1(n3085), 
            .I2(n3039), .I3(GND_net), .O(n3117));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2053_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2052_3_lut (.I0(n3017), .I1(n3084), 
            .I2(n3039), .I3(GND_net), .O(n3116));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2052_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2069_3_lut (.I0(n955), .I1(n3101), 
            .I2(n3039), .I3(GND_net), .O(n3133));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2069_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2068_3_lut (.I0(n3033), .I1(n3100), 
            .I2(n3039), .I3(GND_net), .O(n3132));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2068_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i3_3_lut (.I0(encoder0_position[2]), 
            .I1(n31), .I2(encoder0_position[31]), .I3(GND_net), .O(n956));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i2057_3_lut (.I0(n3022), .I1(n3089), 
            .I2(n3039), .I3(GND_net), .O(n3121));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2057_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1101_7 (.CI(n39715), .I0(n1629), 
            .I1(GND_net), .CO(n39716));
    SB_LUT4 encoder0_position_31__I_0_add_1101_6_lut (.I0(GND_net), .I1(n1630), 
            .I2(GND_net), .I3(n39714), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_5 (.CI(n40217), .I0(n3031), 
            .I1(VCC_net), .CO(n40218));
    SB_CARRY encoder0_position_31__I_0_add_1101_6 (.CI(n39714), .I0(n1630), 
            .I1(GND_net), .CO(n39715));
    SB_LUT4 encoder0_position_31__I_0_i2054_3_lut (.I0(n3019), .I1(n3086), 
            .I2(n3039), .I3(GND_net), .O(n3118));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2054_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2060_3_lut (.I0(n3025), .I1(n3092), 
            .I2(n3039), .I3(GND_net), .O(n3124));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2060_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_673_15_lut (.I0(duty[13]), .I1(n51409), .I2(n12), .I3(n39291), 
            .O(pwm_setpoint_22__N_11[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_15_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i2062_3_lut (.I0(n3027), .I1(n3094), 
            .I2(n3039), .I3(GND_net), .O(n3126));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2062_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1101_5_lut (.I0(GND_net), .I1(n1631), 
            .I2(VCC_net), .I3(n39713), .O(n1698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i2063_3_lut (.I0(n3028), .I1(n3095), 
            .I2(n3039), .I3(GND_net), .O(n3127));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2063_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2058_3_lut (.I0(n3023), .I1(n3090), 
            .I2(n3039), .I3(GND_net), .O(n3122));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2058_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2055_3_lut (.I0(n3020), .I1(n3087), 
            .I2(n3039), .I3(GND_net), .O(n3119));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2055_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1101_5 (.CI(n39713), .I0(n1631), 
            .I1(VCC_net), .CO(n39714));
    SB_LUT4 encoder0_position_31__I_0_i2059_3_lut (.I0(n3024), .I1(n3091), 
            .I2(n3039), .I3(GND_net), .O(n3123));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2059_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2061_3_lut (.I0(n3026), .I1(n3093), 
            .I2(n3039), .I3(GND_net), .O(n3125));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2061_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2064_3_lut (.I0(n3029), .I1(n3096), 
            .I2(n3039), .I3(GND_net), .O(n3128));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2064_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2056_3_lut (.I0(n3021), .I1(n3088), 
            .I2(n3039), .I3(GND_net), .O(n3120));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2056_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_2039_4_lut (.I0(GND_net), .I1(n3032), 
            .I2(GND_net), .I3(n40216), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_4 (.CI(n40216), .I0(n3032), 
            .I1(GND_net), .CO(n40217));
    SB_LUT4 encoder0_position_31__I_0_add_2039_3_lut (.I0(GND_net), .I1(n3033), 
            .I2(VCC_net), .I3(n40215), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1731 (.I0(n3120), .I1(n3128), .I2(n3125), .I3(n3123), 
            .O(n47079));
    defparam i1_4_lut_adj_1731.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_2039_3 (.CI(n40215), .I0(n3033), 
            .I1(VCC_net), .CO(n40216));
    SB_LUT4 encoder0_position_31__I_0_add_2039_2_lut (.I0(GND_net), .I1(n955), 
            .I2(GND_net), .I3(VCC_net), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_2039_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_2039_2 (.CI(VCC_net), .I0(n955), 
            .I1(GND_net), .CO(n40215));
    SB_LUT4 i1_4_lut_adj_1732 (.I0(n3119), .I1(n3122), .I2(n3127), .I3(n3126), 
            .O(n47077));
    defparam i1_4_lut_adj_1732.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1733 (.I0(n47079), .I1(n3124), .I2(n3118), .I3(n3121), 
            .O(n47081));
    defparam i1_4_lut_adj_1733.LUT_INIT = 16'hfffe;
    SB_LUT4 i21528_3_lut (.I0(n956), .I1(n3132), .I2(n3133), .I3(GND_net), 
            .O(n34593));
    defparam i21528_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1734 (.I0(n3116), .I1(n47081), .I2(n3117), .I3(n47077), 
            .O(n47087));
    defparam i1_4_lut_adj_1734.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1735 (.I0(n3129), .I1(n34593), .I2(n3130), .I3(n3131), 
            .O(n45134));
    defparam i1_4_lut_adj_1735.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1736 (.I0(n3114), .I1(n3115), .I2(n45134), .I3(n47087), 
            .O(n47093));
    defparam i1_4_lut_adj_1736.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1737 (.I0(n3111), .I1(n3112), .I2(n3113), .I3(n47093), 
            .O(n47099));
    defparam i1_4_lut_adj_1737.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1738 (.I0(n3108), .I1(n3109), .I2(n3110), .I3(n47099), 
            .O(n47105));
    defparam i1_4_lut_adj_1738.LUT_INIT = 16'hfffe;
    SB_LUT4 i36287_4_lut (.I0(n3106), .I1(n3105), .I2(n3107), .I3(n47105), 
            .O(n3138));
    defparam i36287_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i36449_3_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n26483), .I3(GND_net), .O(n5722));
    defparam i36449_3_lut_3_lut.LUT_INIT = 16'h1515;
    SB_LUT4 i35036_2_lut (.I0(n51546), .I1(byte_transmit_counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n49817));
    defparam i35036_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i34997_2_lut_3_lut (.I0(n62), .I1(delay_counter[31]), .I2(\ID_READOUT_FSM.state [0]), 
            .I3(GND_net), .O(n49714));
    defparam i34997_2_lut_3_lut.LUT_INIT = 16'hf2f2;
    SB_LUT4 i1_2_lut_3_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n26483), .I3(GND_net), .O(n26484));   // verilog/TinyFPGA_B.v(277[7:11])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 encoder0_position_31__I_0_i1976_3_lut (.I0(n2909), .I1(n2976), 
            .I2(n2940), .I3(GND_net), .O(n3008));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1976_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1975_3_lut (.I0(n2908), .I1(n2975), 
            .I2(n2940), .I3(GND_net), .O(n3007));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1975_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1101_4_lut (.I0(GND_net), .I1(n1632), 
            .I2(GND_net), .I3(n39712), .O(n1699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1972_29_lut (.I0(n51169), .I1(n2907), 
            .I2(VCC_net), .I3(n40214), .O(n3006)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1972_28_lut (.I0(GND_net), .I1(n2908), 
            .I2(VCC_net), .I3(n40213), .O(n2975)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_28 (.CI(n40213), .I0(n2908), 
            .I1(VCC_net), .CO(n40214));
    SB_CARRY encoder0_position_31__I_0_add_1101_4 (.CI(n39712), .I0(n1632), 
            .I1(GND_net), .CO(n39713));
    SB_LUT4 encoder0_position_31__I_0_i1979_3_lut (.I0(n2912), .I1(n2979), 
            .I2(n2940), .I3(GND_net), .O(n3011));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1979_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1101_3_lut (.I0(GND_net), .I1(n1633), 
            .I2(VCC_net), .I3(n39711), .O(n1700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1978_3_lut (.I0(n2911), .I1(n2978), 
            .I2(n2940), .I3(GND_net), .O(n3010));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1978_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_27_lut (.I0(GND_net), .I1(n2909), 
            .I2(VCC_net), .I3(n40212), .O(n2976)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_27 (.CI(n40212), .I0(n2909), 
            .I1(VCC_net), .CO(n40213));
    SB_DFFESR delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n5722), 
            .D(n686), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_add_1972_26_lut (.I0(GND_net), .I1(n2910), 
            .I2(VCC_net), .I3(n40211), .O(n2977)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_26 (.CI(n40211), .I0(n2910), 
            .I1(VCC_net), .CO(n40212));
    SB_CARRY add_673_15 (.CI(n39291), .I0(n51409), .I1(n12), .CO(n39292));
    SB_LUT4 encoder0_position_31__I_0_add_1972_25_lut (.I0(GND_net), .I1(n2911), 
            .I2(VCC_net), .I3(n40210), .O(n2978)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_25 (.CI(n40210), .I0(n2911), 
            .I1(VCC_net), .CO(n40211));
    SB_LUT4 encoder0_position_31__I_0_add_1972_24_lut (.I0(GND_net), .I1(n2912), 
            .I2(VCC_net), .I3(n40209), .O(n2979)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_24 (.CI(n40209), .I0(n2912), 
            .I1(VCC_net), .CO(n40210));
    SB_LUT4 encoder0_position_31__I_0_i1977_3_lut (.I0(n2910), .I1(n2977), 
            .I2(n2940), .I3(GND_net), .O(n3009));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1977_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_23_lut (.I0(GND_net), .I1(n2913), 
            .I2(VCC_net), .I3(n40208), .O(n2980)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_23 (.CI(n40208), .I0(n2913), 
            .I1(VCC_net), .CO(n40209));
    SB_LUT4 encoder0_position_31__I_0_add_1972_22_lut (.I0(GND_net), .I1(n2914), 
            .I2(VCC_net), .I3(n40207), .O(n2981)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_22 (.CI(n40207), .I0(n2914), 
            .I1(VCC_net), .CO(n40208));
    SB_LUT4 encoder0_position_31__I_0_add_1972_21_lut (.I0(GND_net), .I1(n2915), 
            .I2(VCC_net), .I3(n40206), .O(n2982)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_21 (.CI(n40206), .I0(n2915), 
            .I1(VCC_net), .CO(n40207));
    SB_LUT4 encoder0_position_31__I_0_add_1972_20_lut (.I0(GND_net), .I1(n2916), 
            .I2(VCC_net), .I3(n40205), .O(n2983)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_20 (.CI(n40205), .I0(n2916), 
            .I1(VCC_net), .CO(n40206));
    SB_LUT4 encoder0_position_31__I_0_add_1972_19_lut (.I0(GND_net), .I1(n2917), 
            .I2(VCC_net), .I3(n40204), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_19 (.CI(n40204), .I0(n2917), 
            .I1(VCC_net), .CO(n40205));
    SB_LUT4 encoder0_position_31__I_0_add_1972_18_lut (.I0(GND_net), .I1(n2918), 
            .I2(VCC_net), .I3(n40203), .O(n2985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_673_14_lut (.I0(duty[12]), .I1(n51409), .I2(n13), .I3(n39290), 
            .O(pwm_setpoint_22__N_11[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_14_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_77_8_lut (.I0(GND_net), .I1(encoder1_position[9]), .I2(GND_net), 
            .I3(n39026), .O(encoder1_position_scaled_23__N_58[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_77_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_3 (.CI(n39711), .I0(n1633), 
            .I1(VCC_net), .CO(n39712));
    SB_LUT4 encoder0_position_31__I_0_add_1101_2_lut (.I0(GND_net), .I1(n941), 
            .I2(GND_net), .I3(VCC_net), .O(n1701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1101_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_673_14 (.CI(n39290), .I0(n51409), .I1(n13), .CO(n39291));
    SB_LUT4 add_673_13_lut (.I0(duty[11]), .I1(n51409), .I2(n14), .I3(n39289), 
            .O(pwm_setpoint_22__N_11[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_13_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i1984_3_lut (.I0(n2917), .I1(n2984), 
            .I2(n2940), .I3(GND_net), .O(n3016));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1984_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1983_3_lut (.I0(n2916), .I1(n2983), 
            .I2(n2940), .I3(GND_net), .O(n3015));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1983_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1972_18 (.CI(n40203), .I0(n2918), 
            .I1(VCC_net), .CO(n40204));
    SB_LUT4 encoder0_position_31__I_0_add_1972_17_lut (.I0(GND_net), .I1(n2919), 
            .I2(VCC_net), .I3(n40202), .O(n2986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_17_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i19 (.Q(delay_counter[19]), .C(CLK_c), .E(n5722), 
            .D(n671), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY encoder0_position_31__I_0_add_1972_17 (.CI(n40202), .I0(n2919), 
            .I1(VCC_net), .CO(n40203));
    SB_LUT4 encoder0_position_31__I_0_i1982_3_lut (.I0(n2915), .I1(n2982), 
            .I2(n2940), .I3(GND_net), .O(n3014));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1982_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1981_3_lut (.I0(n2914), .I1(n2981), 
            .I2(n2940), .I3(GND_net), .O(n3013));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1981_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1972_16_lut (.I0(GND_net), .I1(n2920), 
            .I2(VCC_net), .I3(n40201), .O(n2987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_16 (.CI(n40201), .I0(n2920), 
            .I1(VCC_net), .CO(n40202));
    SB_LUT4 encoder0_position_31__I_0_add_1972_15_lut (.I0(GND_net), .I1(n2921), 
            .I2(VCC_net), .I3(n40200), .O(n2988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_15 (.CI(n40200), .I0(n2921), 
            .I1(VCC_net), .CO(n40201));
    SB_LUT4 encoder0_position_31__I_0_add_1972_14_lut (.I0(GND_net), .I1(n2922), 
            .I2(VCC_net), .I3(n40199), .O(n2989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_14 (.CI(n40199), .I0(n2922), 
            .I1(VCC_net), .CO(n40200));
    SB_LUT4 encoder0_position_31__I_0_add_1972_13_lut (.I0(GND_net), .I1(n2923), 
            .I2(VCC_net), .I3(n40198), .O(n2990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_13 (.CI(n40198), .I0(n2923), 
            .I1(VCC_net), .CO(n40199));
    SB_LUT4 encoder0_position_31__I_0_add_1972_12_lut (.I0(GND_net), .I1(n2924), 
            .I2(VCC_net), .I3(n40197), .O(n2991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_12 (.CI(n40197), .I0(n2924), 
            .I1(VCC_net), .CO(n40198));
    SB_LUT4 encoder0_position_31__I_0_add_1972_11_lut (.I0(GND_net), .I1(n2925), 
            .I2(VCC_net), .I3(n40196), .O(n2992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_11 (.CI(n40196), .I0(n2925), 
            .I1(VCC_net), .CO(n40197));
    SB_LUT4 encoder0_position_31__I_0_add_1972_10_lut (.I0(GND_net), .I1(n2926), 
            .I2(VCC_net), .I3(n40195), .O(n2993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1980_3_lut (.I0(n2913), .I1(n2980), 
            .I2(n2940), .I3(GND_net), .O(n3012));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1980_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i2001_3_lut (.I0(n954), .I1(n3001), 
            .I2(n2940), .I3(GND_net), .O(n3033));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2001_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1972_10 (.CI(n40195), .I0(n2926), 
            .I1(VCC_net), .CO(n40196));
    SB_LUT4 encoder0_position_31__I_0_add_1972_9_lut (.I0(GND_net), .I1(n2927), 
            .I2(VCC_net), .I3(n40194), .O(n2994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1101_2 (.CI(VCC_net), .I0(n941), 
            .I1(GND_net), .CO(n39711));
    SB_LUT4 encoder0_position_31__I_0_add_1034_15_lut (.I0(n50933), .I1(n1521), 
            .I2(VCC_net), .I3(n39710), .O(n1620)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_673_13 (.CI(n39289), .I0(n51409), .I1(n14), .CO(n39290));
    SB_CARRY encoder0_position_31__I_0_add_1972_9 (.CI(n40194), .I0(n2927), 
            .I1(VCC_net), .CO(n40195));
    SB_LUT4 encoder0_position_31__I_0_add_1972_8_lut (.I0(GND_net), .I1(n2928), 
            .I2(VCC_net), .I3(n40193), .O(n2995)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1034_14_lut (.I0(GND_net), .I1(n1522), 
            .I2(VCC_net), .I3(n39709), .O(n1589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_8 (.CI(n40193), .I0(n2928), 
            .I1(VCC_net), .CO(n40194));
    SB_LUT4 encoder0_position_31__I_0_add_1972_7_lut (.I0(GND_net), .I1(n2929), 
            .I2(GND_net), .I3(n40192), .O(n2996)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_14 (.CI(n39709), .I0(n1522), 
            .I1(VCC_net), .CO(n39710));
    SB_LUT4 add_673_12_lut (.I0(duty[10]), .I1(n51409), .I2(n15_adj_4887), 
            .I3(n39288), .O(pwm_setpoint_22__N_11[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_12_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_1436_21_lut (.I0(n51056), .I1(n2115), 
            .I2(VCC_net), .I3(n39819), .O(n2214)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1436_20_lut (.I0(GND_net), .I1(n2116), 
            .I2(VCC_net), .I3(n39818), .O(n2183)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_20 (.CI(n39818), .I0(n2116), 
            .I1(VCC_net), .CO(n39819));
    SB_CARRY add_673_12 (.CI(n39288), .I0(n51409), .I1(n15_adj_4887), 
            .CO(n39289));
    SB_LUT4 encoder0_position_31__I_0_add_1436_19_lut (.I0(GND_net), .I1(n2117), 
            .I2(VCC_net), .I3(n39817), .O(n2184)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_7 (.CI(n40192), .I0(n2929), 
            .I1(GND_net), .CO(n40193));
    SB_CARRY encoder0_position_31__I_0_add_1436_19 (.CI(n39817), .I0(n2117), 
            .I1(VCC_net), .CO(n39818));
    SB_LUT4 encoder0_position_31__I_0_add_1972_6_lut (.I0(GND_net), .I1(n2930), 
            .I2(GND_net), .I3(n40191), .O(n2997)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1436_18_lut (.I0(GND_net), .I1(n2118), 
            .I2(VCC_net), .I3(n39816), .O(n2185)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_673_11_lut (.I0(duty[9]), .I1(n51409), .I2(n16), .I3(n39287), 
            .O(pwm_setpoint_22__N_11[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_11_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_1436_18 (.CI(n39816), .I0(n2118), 
            .I1(VCC_net), .CO(n39817));
    SB_CARRY encoder0_position_31__I_0_add_1972_6 (.CI(n40191), .I0(n2930), 
            .I1(GND_net), .CO(n40192));
    SB_LUT4 encoder0_position_31__I_0_add_1972_5_lut (.I0(GND_net), .I1(n2931), 
            .I2(VCC_net), .I3(n40190), .O(n2998)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_5 (.CI(n40190), .I0(n2931), 
            .I1(VCC_net), .CO(n40191));
    SB_LUT4 encoder0_position_31__I_0_add_1972_4_lut (.I0(GND_net), .I1(n2932), 
            .I2(GND_net), .I3(n40189), .O(n2999)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_4 (.CI(n40189), .I0(n2932), 
            .I1(GND_net), .CO(n40190));
    SB_LUT4 encoder0_position_31__I_0_add_1972_3_lut (.I0(GND_net), .I1(n2933), 
            .I2(VCC_net), .I3(n40188), .O(n3000)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_3 (.CI(n40188), .I0(n2933), 
            .I1(VCC_net), .CO(n40189));
    SB_LUT4 encoder0_position_31__I_0_add_1972_2_lut (.I0(GND_net), .I1(n954), 
            .I2(GND_net), .I3(VCC_net), .O(n3001)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1972_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1972_2 (.CI(VCC_net), .I0(n954), 
            .I1(GND_net), .CO(n40188));
    SB_LUT4 encoder0_position_31__I_0_add_1905_28_lut (.I0(n51137), .I1(n2808), 
            .I2(VCC_net), .I3(n40187), .O(n2907)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1905_27_lut (.I0(GND_net), .I1(n2809), 
            .I2(VCC_net), .I3(n40186), .O(n2876)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_27 (.CI(n40186), .I0(n2809), 
            .I1(VCC_net), .CO(n40187));
    SB_LUT4 encoder0_position_31__I_0_add_1905_26_lut (.I0(GND_net), .I1(n2810), 
            .I2(VCC_net), .I3(n40185), .O(n2877)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_26 (.CI(n40185), .I0(n2810), 
            .I1(VCC_net), .CO(n40186));
    SB_LUT4 encoder0_position_31__I_0_i2000_3_lut (.I0(n2933), .I1(n3000), 
            .I2(n2940), .I3(GND_net), .O(n3032));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i2000_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1905_25_lut (.I0(GND_net), .I1(n2811), 
            .I2(VCC_net), .I3(n40184), .O(n2878)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_25 (.CI(n40184), .I0(n2811), 
            .I1(VCC_net), .CO(n40185));
    SB_LUT4 encoder0_position_31__I_0_add_1034_13_lut (.I0(GND_net), .I1(n1523), 
            .I2(VCC_net), .I3(n39708), .O(n1590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_13 (.CI(n39708), .I0(n1523), 
            .I1(VCC_net), .CO(n39709));
    SB_LUT4 encoder0_position_31__I_0_add_1436_17_lut (.I0(GND_net), .I1(n2119), 
            .I2(VCC_net), .I3(n39815), .O(n2186)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_673_11 (.CI(n39287), .I0(n51409), .I1(n16), .CO(n39288));
    SB_CARRY encoder0_position_31__I_0_add_1436_17 (.CI(n39815), .I0(n2119), 
            .I1(VCC_net), .CO(n39816));
    SB_LUT4 encoder0_position_31__I_0_add_1905_24_lut (.I0(GND_net), .I1(n2812), 
            .I2(VCC_net), .I3(n40183), .O(n2879)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1436_16_lut (.I0(GND_net), .I1(n2120), 
            .I2(VCC_net), .I3(n39814), .O(n2187)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_24 (.CI(n40183), .I0(n2812), 
            .I1(VCC_net), .CO(n40184));
    SB_CARRY encoder0_position_31__I_0_add_1436_16 (.CI(n39814), .I0(n2120), 
            .I1(VCC_net), .CO(n39815));
    SB_LUT4 encoder0_position_31__I_0_add_1034_12_lut (.I0(GND_net), .I1(n1524), 
            .I2(VCC_net), .I3(n39707), .O(n1591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1905_23_lut (.I0(GND_net), .I1(n2813), 
            .I2(VCC_net), .I3(n40182), .O(n2880)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1436_15_lut (.I0(GND_net), .I1(n2121), 
            .I2(VCC_net), .I3(n39813), .O(n2188)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_12 (.CI(n39707), .I0(n1524), 
            .I1(VCC_net), .CO(n39708));
    SB_LUT4 encoder0_position_31__I_0_add_1034_11_lut (.I0(GND_net), .I1(n1525), 
            .I2(VCC_net), .I3(n39706), .O(n1592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_23 (.CI(n40182), .I0(n2813), 
            .I1(VCC_net), .CO(n40183));
    SB_LUT4 encoder0_position_31__I_0_add_1905_22_lut (.I0(GND_net), .I1(n2814), 
            .I2(VCC_net), .I3(n40181), .O(n2881)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_22 (.CI(n40181), .I0(n2814), 
            .I1(VCC_net), .CO(n40182));
    SB_LUT4 encoder0_position_31__I_0_add_1905_21_lut (.I0(GND_net), .I1(n2815), 
            .I2(VCC_net), .I3(n40180), .O(n2882)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_8 (.CI(n38995), .I0(delay_counter[6]), .I1(GND_net), 
            .CO(n38996));
    SB_CARRY encoder0_position_31__I_0_add_1905_21 (.CI(n40180), .I0(n2815), 
            .I1(VCC_net), .CO(n40181));
    SB_LUT4 encoder0_position_31__I_0_add_1905_20_lut (.I0(GND_net), .I1(n2816), 
            .I2(VCC_net), .I3(n40179), .O(n2883)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_20 (.CI(n40179), .I0(n2816), 
            .I1(VCC_net), .CO(n40180));
    SB_LUT4 encoder0_position_31__I_0_add_1905_19_lut (.I0(GND_net), .I1(n2817), 
            .I2(VCC_net), .I3(n40178), .O(n2884)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i4_3_lut (.I0(encoder0_position[3]), 
            .I1(n30), .I2(encoder0_position[31]), .I3(GND_net), .O(n955));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1905_19 (.CI(n40178), .I0(n2817), 
            .I1(VCC_net), .CO(n40179));
    SB_LUT4 encoder0_position_31__I_0_add_1905_18_lut (.I0(GND_net), .I1(n2818), 
            .I2(VCC_net), .I3(n40177), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_18 (.CI(n40177), .I0(n2818), 
            .I1(VCC_net), .CO(n40178));
    SB_CARRY encoder0_position_31__I_0_add_1034_11 (.CI(n39706), .I0(n1525), 
            .I1(VCC_net), .CO(n39707));
    SB_LUT4 add_673_10_lut (.I0(duty[8]), .I1(n51409), .I2(n17), .I3(n39286), 
            .O(pwm_setpoint_22__N_11[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_10_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 add_29_20_lut (.I0(GND_net), .I1(delay_counter[18]), .I2(GND_net), 
            .I3(n39007), .O(n672)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_20 (.CI(n39007), .I0(delay_counter[18]), .I1(GND_net), 
            .CO(n39008));
    SB_LUT4 encoder0_position_31__I_0_add_1905_17_lut (.I0(GND_net), .I1(n2819), 
            .I2(VCC_net), .I3(n40176), .O(n2886)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_17 (.CI(n40176), .I0(n2819), 
            .I1(VCC_net), .CO(n40177));
    SB_LUT4 encoder0_position_31__I_0_add_1905_16_lut (.I0(GND_net), .I1(n2820), 
            .I2(VCC_net), .I3(n40175), .O(n2887)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_29_19_lut (.I0(GND_net), .I1(delay_counter[17]), .I2(GND_net), 
            .I3(n39006), .O(n673)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_16 (.CI(n40175), .I0(n2820), 
            .I1(VCC_net), .CO(n40176));
    SB_LUT4 encoder0_position_31__I_0_add_1905_15_lut (.I0(GND_net), .I1(n2821), 
            .I2(VCC_net), .I3(n40174), .O(n2888)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_29_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(GND_net), 
            .I3(n38994), .O(n685)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_15 (.CI(n40174), .I0(n2821), 
            .I1(VCC_net), .CO(n40175));
    SB_LUT4 encoder0_position_31__I_0_add_1905_14_lut (.I0(GND_net), .I1(n2822), 
            .I2(VCC_net), .I3(n40173), .O(n2889)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_14 (.CI(n40173), .I0(n2822), 
            .I1(VCC_net), .CO(n40174));
    SB_CARRY add_673_10 (.CI(n39286), .I0(n51409), .I1(n17), .CO(n39287));
    SB_LUT4 encoder0_position_31__I_0_i1993_3_lut (.I0(n2926), .I1(n2993), 
            .I2(n2940), .I3(GND_net), .O(n3025));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1993_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_673_9_lut (.I0(duty[7]), .I1(n51409), .I2(n18), .I3(n39285), 
            .O(pwm_setpoint_22__N_11[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_9_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_i1987_3_lut (.I0(n2920), .I1(n2987), 
            .I2(n2940), .I3(GND_net), .O(n3019));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1987_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1990_3_lut (.I0(n2923), .I1(n2990), 
            .I2(n2940), .I3(GND_net), .O(n3022));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1990_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1905_13_lut (.I0(GND_net), .I1(n2823), 
            .I2(VCC_net), .I3(n40172), .O(n2890)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_13 (.CI(n40172), .I0(n2823), 
            .I1(VCC_net), .CO(n40173));
    SB_LUT4 encoder0_position_31__I_0_add_1905_12_lut (.I0(GND_net), .I1(n2824), 
            .I2(VCC_net), .I3(n40171), .O(n2891)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_12 (.CI(n40171), .I0(n2824), 
            .I1(VCC_net), .CO(n40172));
    SB_LUT4 encoder0_position_31__I_0_add_1905_11_lut (.I0(GND_net), .I1(n2825), 
            .I2(VCC_net), .I3(n40170), .O(n2892)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1991_3_lut (.I0(n2924), .I1(n2991), 
            .I2(n2940), .I3(GND_net), .O(n3023));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1991_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1905_11 (.CI(n40170), .I0(n2825), 
            .I1(VCC_net), .CO(n40171));
    SB_LUT4 encoder0_position_31__I_0_i1996_3_lut (.I0(n2929), .I1(n2996), 
            .I2(n2940), .I3(GND_net), .O(n3028));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1996_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1905_10_lut (.I0(GND_net), .I1(n2826), 
            .I2(VCC_net), .I3(n40169), .O(n2893)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_10 (.CI(n40169), .I0(n2826), 
            .I1(VCC_net), .CO(n40170));
    SB_LUT4 encoder0_position_31__I_0_add_1905_9_lut (.I0(GND_net), .I1(n2827), 
            .I2(VCC_net), .I3(n40168), .O(n2894)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_9 (.CI(n40168), .I0(n2827), 
            .I1(VCC_net), .CO(n40169));
    SB_LUT4 encoder0_position_31__I_0_add_1905_8_lut (.I0(GND_net), .I1(n2828), 
            .I2(VCC_net), .I3(n40167), .O(n2895)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_8 (.CI(n40167), .I0(n2828), 
            .I1(VCC_net), .CO(n40168));
    SB_LUT4 encoder0_position_31__I_0_add_1905_7_lut (.I0(GND_net), .I1(n2829), 
            .I2(GND_net), .I3(n40166), .O(n2896)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_7 (.CI(n40166), .I0(n2829), 
            .I1(GND_net), .CO(n40167));
    SB_LUT4 encoder0_position_31__I_0_add_1905_6_lut (.I0(GND_net), .I1(n2830), 
            .I2(GND_net), .I3(n40165), .O(n2897)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_6 (.CI(n40165), .I0(n2830), 
            .I1(GND_net), .CO(n40166));
    SB_LUT4 encoder0_position_31__I_0_add_1905_5_lut (.I0(GND_net), .I1(n2831), 
            .I2(VCC_net), .I3(n40164), .O(n2898)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_5 (.CI(n40164), .I0(n2831), 
            .I1(VCC_net), .CO(n40165));
    SB_LUT4 encoder0_position_31__I_0_add_1905_4_lut (.I0(GND_net), .I1(n2832), 
            .I2(GND_net), .I3(n40163), .O(n2899)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_4 (.CI(n40163), .I0(n2832), 
            .I1(GND_net), .CO(n40164));
    SB_LUT4 encoder0_position_31__I_0_add_1905_3_lut (.I0(GND_net), .I1(n2833), 
            .I2(VCC_net), .I3(n40162), .O(n2900)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1248_3_lut (.I0(n1829), .I1(n1896), 
            .I2(n1851), .I3(GND_net), .O(n1928));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1248_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1905_3 (.CI(n40162), .I0(n2833), 
            .I1(VCC_net), .CO(n40163));
    SB_LUT4 encoder0_position_31__I_0_add_1905_2_lut (.I0(GND_net), .I1(n953), 
            .I2(GND_net), .I3(VCC_net), .O(n2901)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1905_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1905_2 (.CI(VCC_net), .I0(n953), 
            .I1(GND_net), .CO(n40162));
    SB_LUT4 encoder0_position_31__I_0_i1988_3_lut (.I0(n2921), .I1(n2988), 
            .I2(n2940), .I3(GND_net), .O(n3020));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1988_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1999_3_lut (.I0(n2932), .I1(n2999), 
            .I2(n2940), .I3(GND_net), .O(n3031));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1999_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1998_3_lut (.I0(n2931), .I1(n2998), 
            .I2(n2940), .I3(GND_net), .O(n3030));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1998_3_lut.LUT_INIT = 16'hacac;
    SB_DFF \ID_READOUT_FSM.state__i1  (.Q(\ID_READOUT_FSM.state [1]), .C(CLK_c), 
           .D(n17_adj_4890));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFF \ID_READOUT_FSM.state__i0  (.Q(\ID_READOUT_FSM.state [0]), .C(CLK_c), 
           .D(n43285));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFF ID_i0_i7 (.Q(ID[7]), .C(CLK_c), .D(n28771));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFF ID_i0_i6 (.Q(ID[6]), .C(CLK_c), .D(n28770));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFF ID_i0_i5 (.Q(ID[5]), .C(CLK_c), .D(n28769));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFF ID_i0_i4 (.Q(ID[4]), .C(CLK_c), .D(n28768));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFF ID_i0_i3 (.Q(ID[3]), .C(CLK_c), .D(n28767));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFF ID_i0_i2 (.Q(ID[2]), .C(CLK_c), .D(n28766));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_DFF ID_i0_i1 (.Q(ID[1]), .C(CLK_c), .D(n28765));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_i1997_3_lut (.I0(n2930), .I1(n2997), 
            .I2(n2940), .I3(GND_net), .O(n3029));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1997_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1986_3_lut (.I0(n2919), .I1(n2986), 
            .I2(n2940), .I3(GND_net), .O(n3018));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1986_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1985_3_lut (.I0(n2918), .I1(n2985), 
            .I2(n2940), .I3(GND_net), .O(n3017));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1985_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1989_3_lut (.I0(n2922), .I1(n2989), 
            .I2(n2940), .I3(GND_net), .O(n3021));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1989_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1995_3_lut (.I0(n2928), .I1(n2995), 
            .I2(n2940), .I3(GND_net), .O(n3027));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1995_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1994_3_lut (.I0(n2927), .I1(n2994), 
            .I2(n2940), .I3(GND_net), .O(n3026));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1994_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1992_3_lut (.I0(n2925), .I1(n2992), 
            .I2(n2940), .I3(GND_net), .O(n3024));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1992_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1739 (.I0(n3024), .I1(n3026), .I2(n3027), .I3(n3021), 
            .O(n47499));
    defparam i1_4_lut_adj_1739.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1740 (.I0(n3020), .I1(n3028), .I2(n3023), .I3(n3022), 
            .O(n47497));
    defparam i1_4_lut_adj_1740.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1741 (.I0(n47499), .I1(n3019), .I2(n3025), .I3(GND_net), 
            .O(n47501));
    defparam i1_3_lut_adj_1741.LUT_INIT = 16'hfefe;
    SB_LUT4 i21534_3_lut (.I0(n955), .I1(n3032), .I2(n3033), .I3(GND_net), 
            .O(n34599));
    defparam i21534_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1742 (.I0(n3017), .I1(n47501), .I2(n3018), .I3(n47497), 
            .O(n47507));
    defparam i1_4_lut_adj_1742.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1743 (.I0(n3029), .I1(n34599), .I2(n3030), .I3(n3031), 
            .O(n45174));
    defparam i1_4_lut_adj_1743.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1744 (.I0(n3015), .I1(n3016), .I2(n45174), .I3(n47507), 
            .O(n47513));
    defparam i1_4_lut_adj_1744.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1745 (.I0(n3012), .I1(n3013), .I2(n3014), .I3(n47513), 
            .O(n47519));
    defparam i1_4_lut_adj_1745.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1746 (.I0(n3009), .I1(n3010), .I2(n3011), .I3(n47519), 
            .O(n47525));
    defparam i1_4_lut_adj_1746.LUT_INIT = 16'hfffe;
    SB_LUT4 i36253_4_lut (.I0(n3007), .I1(n3006), .I2(n3008), .I3(n47525), 
            .O(n3039));
    defparam i36253_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i10_1_lut (.I0(encoder1_position_scaled[9]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n16_adj_4902));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1909_3_lut (.I0(n2810), .I1(n2877), 
            .I2(n2841), .I3(GND_net), .O(n2909));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1909_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1908_3_lut (.I0(n2809), .I1(n2876), 
            .I2(n2841), .I3(GND_net), .O(n2908));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1908_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1911_3_lut (.I0(n2812), .I1(n2879), 
            .I2(n2841), .I3(GND_net), .O(n2911));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1911_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1910_3_lut (.I0(n2811), .I1(n2878), 
            .I2(n2841), .I3(GND_net), .O(n2910));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1910_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1915_3_lut (.I0(n2816), .I1(n2883), 
            .I2(n2841), .I3(GND_net), .O(n2915));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1915_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1913_3_lut (.I0(n2814), .I1(n2881), 
            .I2(n2841), .I3(GND_net), .O(n2913));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1913_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1918_3_lut (.I0(n2819), .I1(n2886), 
            .I2(n2841), .I3(GND_net), .O(n2918));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1918_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1917_3_lut (.I0(n2818), .I1(n2885), 
            .I2(n2841), .I3(GND_net), .O(n2917));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1917_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1916_3_lut (.I0(n2817), .I1(n2884), 
            .I2(n2841), .I3(GND_net), .O(n2916));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1916_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1921_3_lut (.I0(n2822), .I1(n2889), 
            .I2(n2841), .I3(GND_net), .O(n2921));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1921_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1923_3_lut (.I0(n2824), .I1(n2891), 
            .I2(n2841), .I3(GND_net), .O(n2923));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1923_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1912_3_lut (.I0(n2813), .I1(n2880), 
            .I2(n2841), .I3(GND_net), .O(n2912));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1912_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1914_3_lut (.I0(n2815), .I1(n2882), 
            .I2(n2841), .I3(GND_net), .O(n2914));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1914_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1931_3_lut (.I0(n2832), .I1(n2899), 
            .I2(n2841), .I3(GND_net), .O(n2931));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1931_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1930_3_lut (.I0(n2831), .I1(n2898), 
            .I2(n2841), .I3(GND_net), .O(n2930));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1930_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1929_3_lut (.I0(n2830), .I1(n2897), 
            .I2(n2841), .I3(GND_net), .O(n2929));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1929_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1925_3_lut (.I0(n2826), .I1(n2893), 
            .I2(n2841), .I3(GND_net), .O(n2925));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1925_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1919_3_lut (.I0(n2820), .I1(n2887), 
            .I2(n2841), .I3(GND_net), .O(n2919));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1919_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1928_3_lut (.I0(n2829), .I1(n2896), 
            .I2(n2841), .I3(GND_net), .O(n2928));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1928_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1920_3_lut (.I0(n2821), .I1(n2888), 
            .I2(n2841), .I3(GND_net), .O(n2920));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1920_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1933_3_lut (.I0(n953), .I1(n2901), 
            .I2(n2841), .I3(GND_net), .O(n2933));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1933_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1932_3_lut (.I0(n2833), .I1(n2900), 
            .I2(n2841), .I3(GND_net), .O(n2932));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1932_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i5_3_lut (.I0(encoder0_position[4]), 
            .I1(n29), .I2(encoder0_position[31]), .I3(GND_net), .O(n954));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1926_3_lut (.I0(n2827), .I1(n2894), 
            .I2(n2841), .I3(GND_net), .O(n2926));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1926_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35559_3_lut (.I0(n2724), .I1(n2791), .I2(n2742), .I3(GND_net), 
            .O(n2823));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i35559_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35263_3_lut (.I0(n2823), .I1(n2890), .I2(n2841), .I3(GND_net), 
            .O(n2922));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i35263_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1924_3_lut (.I0(n2825), .I1(n2892), 
            .I2(n2841), .I3(GND_net), .O(n2924));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1924_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1927_3_lut (.I0(n2828), .I1(n2895), 
            .I2(n2841), .I3(GND_net), .O(n2927));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1927_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1747 (.I0(n2920), .I1(n2928), .I2(GND_net), .I3(GND_net), 
            .O(n46895));
    defparam i1_2_lut_adj_1747.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1748 (.I0(n2927), .I1(n2924), .I2(n2922), .I3(n2926), 
            .O(n46899));
    defparam i1_4_lut_adj_1748.LUT_INIT = 16'hfffe;
    SB_LUT4 i21538_3_lut (.I0(n954), .I1(n2932), .I2(n2933), .I3(GND_net), 
            .O(n34603));
    defparam i21538_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1749 (.I0(n2919), .I1(n46899), .I2(n46895), .I3(n2925), 
            .O(n46903));
    defparam i1_4_lut_adj_1749.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1750 (.I0(n2929), .I1(n34603), .I2(n2930), .I3(n2931), 
            .O(n45125));
    defparam i1_4_lut_adj_1750.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1751 (.I0(n2916), .I1(n2917), .I2(n2918), .I3(n46903), 
            .O(n46909));
    defparam i1_4_lut_adj_1751.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1752 (.I0(n2913), .I1(n2915), .I2(n46909), .I3(n45125), 
            .O(n46915));
    defparam i1_4_lut_adj_1752.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1753 (.I0(n2914), .I1(n2912), .I2(n2923), .I3(n2921), 
            .O(n45531));
    defparam i1_4_lut_adj_1753.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1754 (.I0(n2910), .I1(n45531), .I2(n2911), .I3(n46915), 
            .O(n46921));
    defparam i1_4_lut_adj_1754.LUT_INIT = 16'hfffe;
    SB_LUT4 i36220_4_lut (.I0(n2908), .I1(n2907), .I2(n2909), .I3(n46921), 
            .O(n2940));
    defparam i36220_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_1838_27_lut (.I0(n51102), .I1(n2709), 
            .I2(VCC_net), .I3(n40152), .O(n2808)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_i1172_3_lut (.I0(n1721), .I1(n1788), 
            .I2(n1752), .I3(GND_net), .O(n1820));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1172_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1842_3_lut (.I0(n2711), .I1(n2778), 
            .I2(n2742), .I3(GND_net), .O(n2810));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1842_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1841_3_lut (.I0(n2710), .I1(n2777), 
            .I2(n2742), .I3(GND_net), .O(n2809));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1841_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1845_3_lut (.I0(n2714), .I1(n2781), 
            .I2(n2742), .I3(GND_net), .O(n2813));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1845_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1844_3_lut (.I0(n2713), .I1(n2780), 
            .I2(n2742), .I3(GND_net), .O(n2812));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1844_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_26_lut (.I0(GND_net), .I1(n2710), 
            .I2(VCC_net), .I3(n40151), .O(n2777)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_3 (.CI(n38990), .I0(delay_counter[1]), .I1(GND_net), 
            .CO(n38991));
    SB_LUT4 encoder0_position_31__I_0_i1843_3_lut (.I0(n2712), .I1(n2779), 
            .I2(n2742), .I3(GND_net), .O(n2811));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1843_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1851_3_lut (.I0(n2720), .I1(n2787), 
            .I2(n2742), .I3(GND_net), .O(n2819));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1851_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_29_7 (.CI(n38994), .I0(delay_counter[5]), .I1(GND_net), 
            .CO(n38995));
    SB_CARRY encoder0_position_31__I_0_add_1838_26 (.CI(n40151), .I0(n2710), 
            .I1(VCC_net), .CO(n40152));
    SB_LUT4 encoder0_position_31__I_0_add_1838_25_lut (.I0(GND_net), .I1(n2711), 
            .I2(VCC_net), .I3(n40150), .O(n2778)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1850_3_lut (.I0(n2719), .I1(n2786), 
            .I2(n2742), .I3(GND_net), .O(n2818));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1850_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1849_3_lut (.I0(n2718), .I1(n2785), 
            .I2(n2742), .I3(GND_net), .O(n2817));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1849_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1838_25 (.CI(n40150), .I0(n2711), 
            .I1(VCC_net), .CO(n40151));
    SB_LUT4 encoder0_position_31__I_0_add_1838_24_lut (.I0(GND_net), .I1(n2712), 
            .I2(VCC_net), .I3(n40149), .O(n2779)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_24 (.CI(n40149), .I0(n2712), 
            .I1(VCC_net), .CO(n40150));
    SB_LUT4 encoder0_position_31__I_0_add_1838_23_lut (.I0(GND_net), .I1(n2713), 
            .I2(VCC_net), .I3(n40148), .O(n2780)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_23 (.CI(n40148), .I0(n2713), 
            .I1(VCC_net), .CO(n40149));
    SB_LUT4 encoder0_position_31__I_0_add_1838_22_lut (.I0(GND_net), .I1(n2714), 
            .I2(VCC_net), .I3(n40147), .O(n2781)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_22 (.CI(n40147), .I0(n2714), 
            .I1(VCC_net), .CO(n40148));
    SB_CARRY encoder0_position_31__I_0_add_1436_15 (.CI(n39813), .I0(n2121), 
            .I1(VCC_net), .CO(n39814));
    SB_LUT4 encoder0_position_31__I_0_add_1838_21_lut (.I0(GND_net), .I1(n2715), 
            .I2(VCC_net), .I3(n40146), .O(n2782)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_21 (.CI(n40146), .I0(n2715), 
            .I1(VCC_net), .CO(n40147));
    SB_DFFESR delay_counter_i0_i18 (.Q(delay_counter[18]), .C(CLK_c), .E(n5722), 
            .D(n672), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_add_1838_20_lut (.I0(GND_net), .I1(n2716), 
            .I2(VCC_net), .I3(n40145), .O(n2783)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_20 (.CI(n40145), .I0(n2716), 
            .I1(VCC_net), .CO(n40146));
    SB_LUT4 encoder0_position_31__I_0_add_1838_19_lut (.I0(GND_net), .I1(n2717), 
            .I2(VCC_net), .I3(n40144), .O(n2784)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1848_3_lut (.I0(n2717), .I1(n2784), 
            .I2(n2742), .I3(GND_net), .O(n2816));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1848_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1847_3_lut (.I0(n2716), .I1(n2783), 
            .I2(n2742), .I3(GND_net), .O(n2815));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1847_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_29_19 (.CI(n39006), .I0(delay_counter[17]), .I1(GND_net), 
            .CO(n39007));
    SB_LUT4 encoder0_position_31__I_0_i1846_3_lut (.I0(n2715), .I1(n2782), 
            .I2(n2742), .I3(GND_net), .O(n2814));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1846_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_673_9 (.CI(n39285), .I0(n51409), .I1(n18), .CO(n39286));
    SB_LUT4 add_673_8_lut (.I0(duty[6]), .I1(n51409), .I2(n19), .I3(n39284), 
            .O(pwm_setpoint_22__N_11[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_8_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_1034_10_lut (.I0(GND_net), .I1(n1526), 
            .I2(VCC_net), .I3(n39705), .O(n1593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_29_18_lut (.I0(GND_net), .I1(delay_counter[16]), .I2(GND_net), 
            .I3(n39005), .O(n674)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_19 (.CI(n40144), .I0(n2717), 
            .I1(VCC_net), .CO(n40145));
    SB_LUT4 encoder0_position_31__I_0_add_1436_14_lut (.I0(GND_net), .I1(n2122), 
            .I2(VCC_net), .I3(n39812), .O(n2189)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1838_18_lut (.I0(GND_net), .I1(n2718), 
            .I2(VCC_net), .I3(n40143), .O(n2785)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_29_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n690)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1865_3_lut (.I0(n952), .I1(n2801), 
            .I2(n2742), .I3(GND_net), .O(n2833));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1865_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1838_18 (.CI(n40143), .I0(n2718), 
            .I1(VCC_net), .CO(n40144));
    SB_LUT4 encoder0_position_31__I_0_i1864_3_lut (.I0(n2733), .I1(n2800), 
            .I2(n2742), .I3(GND_net), .O(n2832));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1864_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1863_3_lut (.I0(n2732), .I1(n2799), 
            .I2(n2742), .I3(GND_net), .O(n2831));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1863_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_17_lut (.I0(GND_net), .I1(n2719), 
            .I2(VCC_net), .I3(n40142), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i6_3_lut (.I0(encoder0_position[5]), 
            .I1(n28), .I2(encoder0_position[31]), .I3(GND_net), .O(n953));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1838_17 (.CI(n40142), .I0(n2719), 
            .I1(VCC_net), .CO(n40143));
    SB_LUT4 encoder0_position_31__I_0_i1859_3_lut (.I0(n2728), .I1(n2795), 
            .I2(n2742), .I3(GND_net), .O(n2827));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1859_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1854_3_lut (.I0(n2723), .I1(n2790), 
            .I2(n2742), .I3(GND_net), .O(n2822));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1854_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_29_18 (.CI(n39005), .I0(delay_counter[16]), .I1(GND_net), 
            .CO(n39006));
    SB_LUT4 encoder0_position_31__I_0_i1862_3_lut (.I0(n2731), .I1(n2798), 
            .I2(n2742), .I3(GND_net), .O(n2830));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1862_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1861_3_lut (.I0(n2730), .I1(n2797), 
            .I2(n2742), .I3(GND_net), .O(n2829));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1861_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_16_lut (.I0(GND_net), .I1(n2720), 
            .I2(VCC_net), .I3(n40141), .O(n2787)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1860_3_lut (.I0(n2729), .I1(n2796), 
            .I2(n2742), .I3(GND_net), .O(n2828));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1860_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35553_3_lut (.I0(n50505), .I1(pwm_setpoint[14]), .I2(n29_adj_4978), 
            .I3(GND_net), .O(n50506));   // verilog/pwm.v(21[8:24])
    defparam i35553_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1838_16 (.CI(n40141), .I0(n2720), 
            .I1(VCC_net), .CO(n40142));
    SB_LUT4 encoder0_position_31__I_0_add_1838_15_lut (.I0(GND_net), .I1(n2721), 
            .I2(VCC_net), .I3(n40140), .O(n2788)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35032_4_lut (.I0(n33_adj_4981), .I1(n31_adj_4980), .I2(n29_adj_4978), 
            .I3(n50013), .O(n49984));
    defparam i35032_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35580_4_lut (.I0(n30_adj_4979), .I1(n10_adj_4967), .I2(n35), 
            .I3(n49982), .O(n50533));   // verilog/pwm.v(21[8:24])
    defparam i35580_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY encoder0_position_31__I_0_add_1838_15 (.CI(n40140), .I0(n2721), 
            .I1(VCC_net), .CO(n40141));
    SB_LUT4 encoder0_position_31__I_0_add_1838_14_lut (.I0(GND_net), .I1(n2722), 
            .I2(VCC_net), .I3(n40139), .O(n2789)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35272_3_lut (.I0(n50506), .I1(pwm_setpoint[15]), .I2(n31_adj_4980), 
            .I3(GND_net), .O(n50224));   // verilog/pwm.v(21[8:24])
    defparam i35272_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1838_14 (.CI(n40139), .I0(n2722), 
            .I1(VCC_net), .CO(n40140));
    SB_LUT4 i35554_3_lut (.I0(n6_adj_4963), .I1(pwm_setpoint[10]), .I2(n21_adj_4974), 
            .I3(GND_net), .O(n50507));   // verilog/pwm.v(21[8:24])
    defparam i35554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35555_3_lut (.I0(n50507), .I1(pwm_setpoint[11]), .I2(n23_adj_4975), 
            .I3(GND_net), .O(n50508));   // verilog/pwm.v(21[8:24])
    defparam i35555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35320_4_lut (.I0(n23_adj_4975), .I1(n21_adj_4974), .I2(n19_adj_4973), 
            .I3(n50024), .O(n50273));
    defparam i35320_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 encoder0_position_31__I_0_add_1838_13_lut (.I0(GND_net), .I1(n2723), 
            .I2(VCC_net), .I3(n40138), .O(n2790)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35512_3_lut (.I0(n8_adj_4965), .I1(pwm_setpoint[9]), .I2(n19_adj_4973), 
            .I3(GND_net), .O(n50465));   // verilog/pwm.v(21[8:24])
    defparam i35512_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35270_3_lut (.I0(n50508), .I1(pwm_setpoint[12]), .I2(n25_adj_4976), 
            .I3(GND_net), .O(n50222));   // verilog/pwm.v(21[8:24])
    defparam i35270_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1838_13 (.CI(n40138), .I0(n2723), 
            .I1(VCC_net), .CO(n40139));
    SB_LUT4 encoder0_position_31__I_0_add_1838_12_lut (.I0(GND_net), .I1(n2724), 
            .I2(VCC_net), .I3(n40137), .O(n2791)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35556_4_lut (.I0(n33_adj_4981), .I1(n31_adj_4980), .I2(n29_adj_4978), 
            .I3(n50018), .O(n50509));
    defparam i35556_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1838_12 (.CI(n40137), .I0(n2724), 
            .I1(VCC_net), .CO(n40138));
    SB_LUT4 encoder0_position_31__I_0_add_1838_11_lut (.I0(GND_net), .I1(n2725), 
            .I2(VCC_net), .I3(n40136), .O(n2792)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_11 (.CI(n40136), .I0(n2725), 
            .I1(VCC_net), .CO(n40137));
    SB_LUT4 encoder0_position_31__I_0_add_1838_10_lut (.I0(GND_net), .I1(n2726), 
            .I2(VCC_net), .I3(n40135), .O(n2793)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35688_4_lut (.I0(n50224), .I1(n50533), .I2(n35), .I3(n49984), 
            .O(n50641));   // verilog/pwm.v(21[8:24])
    defparam i35688_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY encoder0_position_31__I_0_add_1838_10 (.CI(n40135), .I0(n2726), 
            .I1(VCC_net), .CO(n40136));
    SB_LUT4 i35578_4_lut (.I0(n50222), .I1(n50465), .I2(n25_adj_4976), 
            .I3(n50273), .O(n50531));   // verilog/pwm.v(21[8:24])
    defparam i35578_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35720_4_lut (.I0(n50531), .I1(n50641), .I2(n35), .I3(n50509), 
            .O(n50673));   // verilog/pwm.v(21[8:24])
    defparam i35720_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_add_1838_9_lut (.I0(GND_net), .I1(n2727), 
            .I2(VCC_net), .I3(n40134), .O(n2794)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35721_3_lut (.I0(n50673), .I1(pwm_setpoint[18]), .I2(pwm_counter[18]), 
            .I3(GND_net), .O(n50674));   // verilog/pwm.v(21[8:24])
    defparam i35721_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_31__I_0_add_1838_9 (.CI(n40134), .I0(n2727), 
            .I1(VCC_net), .CO(n40135));
    SB_LUT4 encoder0_position_31__I_0_add_1838_8_lut (.I0(GND_net), .I1(n2728), 
            .I2(VCC_net), .I3(n40133), .O(n2795)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35719_3_lut (.I0(n50674), .I1(pwm_setpoint[19]), .I2(pwm_counter[19]), 
            .I3(GND_net), .O(n50672));   // verilog/pwm.v(21[8:24])
    defparam i35719_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_31__I_0_add_1838_8 (.CI(n40133), .I0(n2728), 
            .I1(VCC_net), .CO(n40134));
    SB_LUT4 encoder0_position_31__I_0_i1857_3_lut (.I0(n2726), .I1(n2793), 
            .I2(n2742), .I3(GND_net), .O(n2825));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1857_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35640_3_lut (.I0(n50672), .I1(pwm_setpoint[20]), .I2(pwm_counter[20]), 
            .I3(GND_net), .O(n50593));   // verilog/pwm.v(21[8:24])
    defparam i35640_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_31__I_0_add_1838_7_lut (.I0(GND_net), .I1(n2729), 
            .I2(GND_net), .I3(n40132), .O(n2796)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_7 (.CI(n40132), .I0(n2729), 
            .I1(GND_net), .CO(n40133));
    SB_LUT4 encoder0_position_31__I_0_add_1838_6_lut (.I0(GND_net), .I1(n2730), 
            .I2(GND_net), .I3(n40131), .O(n2797)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_6 (.CI(n40131), .I0(n2730), 
            .I1(GND_net), .CO(n40132));
    SB_LUT4 encoder0_position_31__I_0_add_1838_5_lut (.I0(GND_net), .I1(n2731), 
            .I2(VCC_net), .I3(n40130), .O(n2798)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35641_3_lut (.I0(n50593), .I1(pwm_setpoint[21]), .I2(pwm_counter[21]), 
            .I3(GND_net), .O(n50594));   // verilog/pwm.v(21[8:24])
    defparam i35641_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_31__I_0_add_1838_5 (.CI(n40130), .I0(n2731), 
            .I1(VCC_net), .CO(n40131));
    SB_LUT4 i35607_3_lut (.I0(n50594), .I1(pwm_setpoint[22]), .I2(pwm_counter[22]), 
            .I3(GND_net), .O(n50560));   // verilog/pwm.v(21[8:24])
    defparam i35607_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i29922_3_lut (.I0(n3_adj_4952), .I1(n6535), .I2(n44804), .I3(GND_net), 
            .O(n44805));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i29922_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29923_3_lut (.I0(encoder0_position[30]), .I1(n44805), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n829));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i29923_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1838_4_lut (.I0(GND_net), .I1(n2732), 
            .I2(GND_net), .I3(n40129), .O(n2799)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_4 (.CI(n40129), .I0(n2732), 
            .I1(GND_net), .CO(n40130));
    SB_LUT4 encoder0_position_31__I_0_i1171_3_lut (.I0(n1720), .I1(n1787), 
            .I2(n1752), .I3(GND_net), .O(n1819));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1171_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1858_rep_14_3_lut (.I0(n2727), .I1(n2794), 
            .I2(n2742), .I3(GND_net), .O(n2826));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1858_rep_14_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1838_3_lut (.I0(GND_net), .I1(n2733), 
            .I2(VCC_net), .I3(n40128), .O(n2800)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_3 (.CI(n40128), .I0(n2733), 
            .I1(VCC_net), .CO(n40129));
    SB_LUT4 encoder0_position_31__I_0_i568_3_lut (.I0(n829), .I1(n896), 
            .I2(n861), .I3(GND_net), .O(n928));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i568_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1838_2_lut (.I0(GND_net), .I1(n952), 
            .I2(GND_net), .I3(VCC_net), .O(n2801)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1838_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1838_2 (.CI(VCC_net), .I0(n952), 
            .I1(GND_net), .CO(n40128));
    SB_LUT4 encoder0_position_31__I_0_add_1771_26_lut (.I0(n50740), .I1(n2610), 
            .I2(VCC_net), .I3(n40127), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_31__I_0_add_1436_14 (.CI(n39812), .I0(n2122), 
            .I1(VCC_net), .CO(n39813));
    SB_LUT4 encoder0_position_31__I_0_add_1771_25_lut (.I0(GND_net), .I1(n2611), 
            .I2(VCC_net), .I3(n40126), .O(n2678)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i635_3_lut (.I0(n928), .I1(n995), 
            .I2(n960), .I3(GND_net), .O(n1027));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i635_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1771_25 (.CI(n40126), .I0(n2611), 
            .I1(VCC_net), .CO(n40127));
    SB_LUT4 i29928_3_lut (.I0(n6_adj_4949), .I1(n6538), .I2(n44804), .I3(GND_net), 
            .O(n44811));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i29928_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1771_24_lut (.I0(GND_net), .I1(n2612), 
            .I2(VCC_net), .I3(n40125), .O(n2679)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35442_3_lut (.I0(n2623), .I1(n2690), .I2(n2643), .I3(GND_net), 
            .O(n2722));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i35442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35443_3_lut (.I0(n2722), .I1(n2789), .I2(n2742), .I3(GND_net), 
            .O(n2821));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i35443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29929_3_lut (.I0(encoder0_position[27]), .I1(n44811), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n832));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i29929_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1771_24 (.CI(n40125), .I0(n2612), 
            .I1(VCC_net), .CO(n40126));
    SB_LUT4 encoder0_position_31__I_0_add_1771_23_lut (.I0(GND_net), .I1(n2613), 
            .I2(VCC_net), .I3(n40124), .O(n2680)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_23 (.CI(n40124), .I0(n2613), 
            .I1(VCC_net), .CO(n40125));
    SB_LUT4 encoder0_position_31__I_0_add_1771_22_lut (.I0(GND_net), .I1(n2614), 
            .I2(VCC_net), .I3(n40123), .O(n2681)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_22 (.CI(n40123), .I0(n2614), 
            .I1(VCC_net), .CO(n40124));
    SB_LUT4 encoder0_position_31__I_0_add_1771_21_lut (.I0(GND_net), .I1(n2615), 
            .I2(VCC_net), .I3(n40122), .O(n2682)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_21 (.CI(n40122), .I0(n2615), 
            .I1(VCC_net), .CO(n40123));
    SB_LUT4 encoder0_position_31__I_0_i571_3_lut (.I0(n832), .I1(n899), 
            .I2(n861), .I3(GND_net), .O(n931));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i571_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i27_3_lut (.I0(encoder0_position[26]), 
            .I1(n7_adj_4948), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n731));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i27_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1771_20_lut (.I0(GND_net), .I1(n2616), 
            .I2(VCC_net), .I3(n40121), .O(n2683)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1755 (.I0(n4_adj_4951), .I1(n5_adj_4950), .I2(n731), 
            .I3(n6_adj_4949), .O(n5_adj_4912));
    defparam i1_4_lut_adj_1755.LUT_INIT = 16'heeea;
    SB_LUT4 i1_3_lut_adj_1756 (.I0(n3_adj_4952), .I1(n2_adj_4953), .I2(n5_adj_4912), 
            .I3(GND_net), .O(n44804));
    defparam i1_3_lut_adj_1756.LUT_INIT = 16'h8080;
    SB_CARRY encoder0_position_31__I_0_add_1771_20 (.CI(n40121), .I0(n2616), 
            .I1(VCC_net), .CO(n40122));
    SB_LUT4 encoder0_position_31__I_0_add_1771_19_lut (.I0(GND_net), .I1(n2617), 
            .I2(VCC_net), .I3(n40120), .O(n2684)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i29930_3_lut (.I0(n7_adj_4948), .I1(n6539), .I2(n44804), .I3(GND_net), 
            .O(n44813));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i29930_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1771_19 (.CI(n40120), .I0(n2617), 
            .I1(VCC_net), .CO(n40121));
    SB_LUT4 i35440_3_lut (.I0(n2622), .I1(n2689), .I2(n2643), .I3(GND_net), 
            .O(n2721));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i35440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i29931_3_lut (.I0(encoder0_position[26]), .I1(n44813), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n833));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i29931_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1771_18_lut (.I0(GND_net), .I1(n2618), 
            .I2(VCC_net), .I3(n40119), .O(n2685)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_18 (.CI(n40119), .I0(n2618), 
            .I1(VCC_net), .CO(n40120));
    SB_LUT4 encoder0_position_31__I_0_add_1771_17_lut (.I0(GND_net), .I1(n2619), 
            .I2(VCC_net), .I3(n40118), .O(n2686)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_17 (.CI(n40118), .I0(n2619), 
            .I1(VCC_net), .CO(n40119));
    SB_LUT4 encoder0_position_31__I_0_add_1771_16_lut (.I0(GND_net), .I1(n2620), 
            .I2(VCC_net), .I3(n40117), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_16 (.CI(n40117), .I0(n2620), 
            .I1(VCC_net), .CO(n40118));
    SB_LUT4 encoder0_position_31__I_0_add_1771_15_lut (.I0(GND_net), .I1(n2621), 
            .I2(VCC_net), .I3(n40116), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_15 (.CI(n40116), .I0(n2621), 
            .I1(VCC_net), .CO(n40117));
    SB_CARRY add_673_8 (.CI(n39284), .I0(n51409), .I1(n19), .CO(n39285));
    SB_LUT4 encoder0_position_31__I_0_add_1771_14_lut (.I0(GND_net), .I1(n2622), 
            .I2(VCC_net), .I3(n40115), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_14 (.CI(n40115), .I0(n2622), 
            .I1(VCC_net), .CO(n40116));
    SB_LUT4 add_673_7_lut (.I0(duty[5]), .I1(n51409), .I2(n20), .I3(n39283), 
            .O(pwm_setpoint_22__N_11[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_7_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_1771_13_lut (.I0(GND_net), .I1(n2623), 
            .I2(VCC_net), .I3(n40114), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_13 (.CI(n40114), .I0(n2623), 
            .I1(VCC_net), .CO(n40115));
    SB_LUT4 i35441_3_lut (.I0(n2721), .I1(n2788), .I2(n2742), .I3(GND_net), 
            .O(n2820));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i35441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1771_12_lut (.I0(GND_net), .I1(n2624), 
            .I2(VCC_net), .I3(n40113), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_12 (.CI(n40113), .I0(n2624), 
            .I1(VCC_net), .CO(n40114));
    SB_LUT4 encoder0_position_31__I_0_add_1771_11_lut (.I0(GND_net), .I1(n2625), 
            .I2(VCC_net), .I3(n40112), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_11 (.CI(n40112), .I0(n2625), 
            .I1(VCC_net), .CO(n40113));
    SB_LUT4 encoder0_position_31__I_0_add_1771_10_lut (.I0(GND_net), .I1(n2626), 
            .I2(VCC_net), .I3(n40111), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_10 (.CI(n40111), .I0(n2626), 
            .I1(VCC_net), .CO(n40112));
    SB_LUT4 encoder0_position_31__I_0_add_1771_9_lut (.I0(GND_net), .I1(n2627), 
            .I2(VCC_net), .I3(n40110), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_9 (.CI(n40110), .I0(n2627), 
            .I1(VCC_net), .CO(n40111));
    SB_LUT4 encoder0_position_31__I_0_add_1771_8_lut (.I0(GND_net), .I1(n2628), 
            .I2(VCC_net), .I3(n40109), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_8 (.CI(n40109), .I0(n2628), 
            .I1(VCC_net), .CO(n40110));
    SB_LUT4 encoder0_position_31__I_0_add_1771_7_lut (.I0(GND_net), .I1(n2629), 
            .I2(GND_net), .I3(n40108), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_7 (.CI(n40108), .I0(n2629), 
            .I1(GND_net), .CO(n40109));
    SB_LUT4 encoder0_position_31__I_0_i572_3_lut (.I0(n833), .I1(n900), 
            .I2(n861), .I3(GND_net), .O(n932));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i572_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1771_6_lut (.I0(GND_net), .I1(n2630), 
            .I2(GND_net), .I3(n40107), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_6 (.CI(n40107), .I0(n2630), 
            .I1(GND_net), .CO(n40108));
    SB_LUT4 encoder0_position_31__I_0_add_1771_5_lut (.I0(GND_net), .I1(n2631), 
            .I2(VCC_net), .I3(n40106), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_5 (.CI(n40106), .I0(n2631), 
            .I1(VCC_net), .CO(n40107));
    SB_LUT4 encoder0_position_31__I_0_add_1771_4_lut (.I0(GND_net), .I1(n2632), 
            .I2(GND_net), .I3(n40105), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_4 (.CI(n40105), .I0(n2632), 
            .I1(GND_net), .CO(n40106));
    SB_LUT4 encoder0_position_31__I_0_add_1436_13_lut (.I0(GND_net), .I1(n2123), 
            .I2(VCC_net), .I3(n39811), .O(n2190)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1771_3_lut (.I0(GND_net), .I1(n2633), 
            .I2(VCC_net), .I3(n40104), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_3 (.CI(n40104), .I0(n2633), 
            .I1(VCC_net), .CO(n40105));
    SB_LUT4 encoder0_position_31__I_0_add_1771_2_lut (.I0(GND_net), .I1(n951), 
            .I2(GND_net), .I3(VCC_net), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1771_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1771_2 (.CI(VCC_net), .I0(n951), 
            .I1(GND_net), .CO(n40104));
    SB_LUT4 encoder0_position_31__I_0_add_1704_25_lut (.I0(n51390), .I1(n2511), 
            .I2(VCC_net), .I3(n40103), .O(n2610)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1704_24_lut (.I0(GND_net), .I1(n2512), 
            .I2(VCC_net), .I3(n40102), .O(n2579)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_24 (.CI(n40102), .I0(n2512), 
            .I1(VCC_net), .CO(n40103));
    SB_LUT4 encoder0_position_31__I_0_i1174_3_lut (.I0(n1723), .I1(n1790), 
            .I2(n1752), .I3(GND_net), .O(n1822));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1174_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_23_lut (.I0(GND_net), .I1(n2513), 
            .I2(VCC_net), .I3(n40101), .O(n2580)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1856_3_lut (.I0(n2725), .I1(n2792), 
            .I2(n2742), .I3(GND_net), .O(n2824));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1856_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1436_13 (.CI(n39811), .I0(n2123), 
            .I1(VCC_net), .CO(n39812));
    SB_CARRY encoder0_position_31__I_0_add_1034_10 (.CI(n39705), .I0(n1526), 
            .I1(VCC_net), .CO(n39706));
    SB_LUT4 encoder0_position_31__I_0_add_1034_9_lut (.I0(GND_net), .I1(n1527), 
            .I2(VCC_net), .I3(n39704), .O(n1594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_3_lut_adj_1757 (.I0(n2824), .I1(n2820), .I2(n2821), .I3(GND_net), 
            .O(n47451));
    defparam i1_3_lut_adj_1757.LUT_INIT = 16'hfefe;
    SB_LUT4 add_29_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(GND_net), 
            .I3(n39004), .O(n675)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_23 (.CI(n40101), .I0(n2513), 
            .I1(VCC_net), .CO(n40102));
    SB_LUT4 i1_4_lut_adj_1758 (.I0(n2826), .I1(n2825), .I2(n2823), .I3(n2828), 
            .O(n47453));
    defparam i1_4_lut_adj_1758.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1704_22_lut (.I0(GND_net), .I1(n2514), 
            .I2(VCC_net), .I3(n40100), .O(n2581)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_22 (.CI(n40100), .I0(n2514), 
            .I1(VCC_net), .CO(n40101));
    SB_LUT4 encoder0_position_31__I_0_add_1704_21_lut (.I0(GND_net), .I1(n2515), 
            .I2(VCC_net), .I3(n40099), .O(n2582)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1759 (.I0(n47453), .I1(n47451), .I2(n2822), .I3(n2827), 
            .O(n47457));
    defparam i1_4_lut_adj_1759.LUT_INIT = 16'hfffe;
    SB_LUT4 i21639_4_lut (.I0(n953), .I1(n2831), .I2(n2832), .I3(n2833), 
            .O(n34707));
    defparam i21639_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1760 (.I0(n2817), .I1(n2818), .I2(n47457), .I3(n2819), 
            .O(n47463));
    defparam i1_4_lut_adj_1760.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1173_3_lut (.I0(n1722), .I1(n1789), 
            .I2(n1752), .I3(GND_net), .O(n1821));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1173_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_21 (.CI(n40099), .I0(n2515), 
            .I1(VCC_net), .CO(n40100));
    SB_LUT4 encoder0_position_31__I_0_add_1704_20_lut (.I0(GND_net), .I1(n2516), 
            .I2(VCC_net), .I3(n40098), .O(n2583)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1761 (.I0(n47463), .I1(n2829), .I2(n34707), .I3(n2830), 
            .O(n47465));
    defparam i1_4_lut_adj_1761.LUT_INIT = 16'heaaa;
    SB_CARRY encoder0_position_31__I_0_add_1704_20 (.CI(n40098), .I0(n2516), 
            .I1(VCC_net), .CO(n40099));
    SB_LUT4 i1_4_lut_adj_1762 (.I0(n2814), .I1(n2815), .I2(n2816), .I3(n47465), 
            .O(n47471));
    defparam i1_4_lut_adj_1762.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1763 (.I0(n2811), .I1(n2812), .I2(n2813), .I3(n47471), 
            .O(n47477));
    defparam i1_4_lut_adj_1763.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1183_3_lut (.I0(n1732), .I1(n1799), 
            .I2(n1752), .I3(GND_net), .O(n1831));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1183_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_19_lut (.I0(GND_net), .I1(n2517), 
            .I2(VCC_net), .I3(n40097), .O(n2584)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_19 (.CI(n40097), .I0(n2517), 
            .I1(VCC_net), .CO(n40098));
    SB_CARRY add_673_7 (.CI(n39283), .I0(n51409), .I1(n20), .CO(n39284));
    SB_LUT4 encoder0_position_31__I_0_add_1436_12_lut (.I0(GND_net), .I1(n2124), 
            .I2(VCC_net), .I3(n39810), .O(n2191)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_12 (.CI(n39810), .I0(n2124), 
            .I1(VCC_net), .CO(n39811));
    SB_LUT4 add_673_6_lut (.I0(duty[4]), .I1(n51409), .I2(n21), .I3(n39282), 
            .O(pwm_setpoint_22__N_11[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_6_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_1034_9 (.CI(n39704), .I0(n1527), 
            .I1(VCC_net), .CO(n39705));
    SB_LUT4 i36188_4_lut (.I0(n2809), .I1(n2808), .I2(n2810), .I3(n47477), 
            .O(n2841));
    defparam i36188_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_1436_11_lut (.I0(GND_net), .I1(n2125), 
            .I2(VCC_net), .I3(n39809), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_83_i10_4_lut (.I0(encoder1_position_scaled[9]), .I1(displacement[9]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[9]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i10_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_add_1034_8_lut (.I0(GND_net), .I1(n1528), 
            .I2(VCC_net), .I3(n39703), .O(n1595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_18_lut (.I0(GND_net), .I1(n2518), 
            .I2(VCC_net), .I3(n40096), .O(n2585)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_673_6 (.CI(n39282), .I0(n51409), .I1(n21), .CO(n39283));
    SB_LUT4 add_673_5_lut (.I0(duty[3]), .I1(n51409), .I2(n22), .I3(n39281), 
            .O(pwm_setpoint_22__N_11[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_5_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_673_5 (.CI(n39281), .I0(n51409), .I1(n22), .CO(n39282));
    SB_CARRY encoder0_position_31__I_0_add_1704_18 (.CI(n40096), .I0(n2518), 
            .I1(VCC_net), .CO(n40097));
    SB_LUT4 add_673_4_lut (.I0(duty[2]), .I1(n51409), .I2(n23), .I3(n39280), 
            .O(pwm_setpoint_22__N_11[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_4_lut.LUT_INIT = 16'h8BB8;
    SB_LUT4 encoder0_position_31__I_0_add_1704_17_lut (.I0(GND_net), .I1(n2519), 
            .I2(VCC_net), .I3(n40095), .O(n2586)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1182_3_lut (.I0(n1731), .I1(n1798), 
            .I2(n1752), .I3(GND_net), .O(n1830));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1182_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_17 (.CI(n40095), .I0(n2519), 
            .I1(VCC_net), .CO(n40096));
    SB_LUT4 encoder0_position_31__I_0_i1181_3_lut (.I0(n1730), .I1(n1797), 
            .I2(n1752), .I3(GND_net), .O(n1829));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1181_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_16_lut (.I0(GND_net), .I1(n2520), 
            .I2(VCC_net), .I3(n40094), .O(n2587)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_16 (.CI(n40094), .I0(n2520), 
            .I1(VCC_net), .CO(n40095));
    SB_CARRY encoder0_position_31__I_0_add_1034_8 (.CI(n39703), .I0(n1528), 
            .I1(VCC_net), .CO(n39704));
    SB_LUT4 add_1890_7_lut (.I0(GND_net), .I1(n621), .I2(GND_net), .I3(n39380), 
            .O(n6534)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1890_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_673_4 (.CI(n39280), .I0(n51409), .I1(n23), .CO(n39281));
    SB_LUT4 encoder0_position_31__I_0_add_1704_15_lut (.I0(GND_net), .I1(n2521), 
            .I2(VCC_net), .I3(n40093), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_15 (.CI(n40093), .I0(n2521), 
            .I1(VCC_net), .CO(n40094));
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i11_1_lut (.I0(encoder1_position_scaled[10]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n15_adj_4901));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_add_1704_14_lut (.I0(GND_net), .I1(n2522), 
            .I2(VCC_net), .I3(n40092), .O(n2589)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1890_6_lut (.I0(GND_net), .I1(n622), .I2(GND_net), .I3(n39379), 
            .O(n6535)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1890_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_11 (.CI(n39809), .I0(n2125), 
            .I1(VCC_net), .CO(n39810));
    SB_LUT4 add_673_3_lut (.I0(duty[1]), .I1(n51409), .I2(n24), .I3(n39279), 
            .O(pwm_setpoint_22__N_11[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_3_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY add_1890_6 (.CI(n39379), .I0(n622), .I1(GND_net), .CO(n39380));
    SB_CARRY encoder0_position_31__I_0_add_1704_14 (.CI(n40092), .I0(n2522), 
            .I1(VCC_net), .CO(n40093));
    SB_LUT4 encoder0_position_31__I_0_add_1704_13_lut (.I0(GND_net), .I1(n2523), 
            .I2(VCC_net), .I3(n40091), .O(n2590)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_673_3 (.CI(n39279), .I0(n51409), .I1(n24), .CO(n39280));
    SB_CARRY encoder0_position_31__I_0_add_1704_13 (.CI(n40091), .I0(n2523), 
            .I1(VCC_net), .CO(n40092));
    SB_LUT4 encoder0_position_31__I_0_add_1704_12_lut (.I0(GND_net), .I1(n2524), 
            .I2(VCC_net), .I3(n40090), .O(n2591)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_1890_5_lut (.I0(GND_net), .I1(n623), .I2(VCC_net), .I3(n39378), 
            .O(n6536)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1890_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1778_3_lut (.I0(n2615), .I1(n2682), 
            .I2(n2643), .I3(GND_net), .O(n2714));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1778_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_12 (.CI(n40090), .I0(n2524), 
            .I1(VCC_net), .CO(n40091));
    SB_LUT4 encoder0_position_31__I_0_i1104_3_lut (.I0(n1621), .I1(n1688), 
            .I2(n1653), .I3(GND_net), .O(n1720));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1104_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_11_lut (.I0(GND_net), .I1(n2525), 
            .I2(VCC_net), .I3(n40089), .O(n2592)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_673_2_lut (.I0(duty[0]), .I1(n51409), .I2(n25), .I3(VCC_net), 
            .O(pwm_setpoint_22__N_11[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_673_2_lut.LUT_INIT = 16'h8BB8;
    SB_CARRY encoder0_position_31__I_0_add_1704_11 (.CI(n40089), .I0(n2525), 
            .I1(VCC_net), .CO(n40090));
    SB_LUT4 encoder0_position_31__I_0_add_1034_7_lut (.I0(GND_net), .I1(n1529), 
            .I2(GND_net), .I3(n39702), .O(n1596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1704_10_lut (.I0(GND_net), .I1(n2526), 
            .I2(VCC_net), .I3(n40088), .O(n2593)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1777_3_lut (.I0(n2614), .I1(n2681), 
            .I2(n2643), .I3(GND_net), .O(n2713));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1777_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_10 (.CI(n40088), .I0(n2526), 
            .I1(VCC_net), .CO(n40089));
    SB_LUT4 encoder0_position_31__I_0_add_1704_9_lut (.I0(GND_net), .I1(n2527), 
            .I2(VCC_net), .I3(n40087), .O(n2594)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_29_17 (.CI(n39004), .I0(delay_counter[15]), .I1(GND_net), 
            .CO(n39005));
    SB_LUT4 encoder0_position_31__I_0_i1176_3_lut (.I0(n1725), .I1(n1792), 
            .I2(n1752), .I3(GND_net), .O(n1824));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1176_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1436_10_lut (.I0(GND_net), .I1(n2126), 
            .I2(VCC_net), .I3(n39808), .O(n2193)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1776_3_lut (.I0(n2613), .I1(n2680), 
            .I2(n2643), .I3(GND_net), .O(n2712));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1776_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_29_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(GND_net), 
            .I3(n38993), .O(n686)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1775_3_lut (.I0(n2612), .I1(n2679), 
            .I2(n2643), .I3(GND_net), .O(n2711));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1775_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_9 (.CI(n40087), .I0(n2527), 
            .I1(VCC_net), .CO(n40088));
    SB_LUT4 encoder0_position_31__I_0_i1774_3_lut (.I0(n2611), .I1(n2678), 
            .I2(n2643), .I3(GND_net), .O(n2710));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1774_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_8_lut (.I0(GND_net), .I1(n2528), 
            .I2(VCC_net), .I3(n40086), .O(n2595)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_22_lut (.I0(GND_net), .I1(n2214), 
            .I2(VCC_net), .I3(n39920), .O(n2281)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1780_3_lut (.I0(n2617), .I1(n2684), 
            .I2(n2643), .I3(GND_net), .O(n2716));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1780_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1034_7 (.CI(n39702), .I0(n1529), 
            .I1(GND_net), .CO(n39703));
    SB_CARRY add_1890_5 (.CI(n39378), .I0(n623), .I1(VCC_net), .CO(n39379));
    SB_LUT4 add_29_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(GND_net), 
            .I3(n39003), .O(n676)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_8 (.CI(n40086), .I0(n2528), 
            .I1(VCC_net), .CO(n40087));
    SB_LUT4 encoder0_position_31__I_0_i1779_3_lut (.I0(n2616), .I1(n2683), 
            .I2(n2643), .I3(GND_net), .O(n2715));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1779_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1890_4_lut (.I0(GND_net), .I1(n516), .I2(GND_net), .I3(n39377), 
            .O(n6537)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1890_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1175_3_lut (.I0(n1724), .I1(n1791), 
            .I2(n1752), .I3(GND_net), .O(n1823));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1175_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1034_6_lut (.I0(GND_net), .I1(n1530), 
            .I2(GND_net), .I3(n39701), .O(n1597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1783_3_lut (.I0(n2620), .I1(n2687), 
            .I2(n2643), .I3(GND_net), .O(n2719));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1783_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1704_7_lut (.I0(GND_net), .I1(n2529), 
            .I2(GND_net), .I3(n40085), .O(n2596)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1782_3_lut (.I0(n2619), .I1(n2686), 
            .I2(n2643), .I3(GND_net), .O(n2718));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1782_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1436_10 (.CI(n39808), .I0(n2126), 
            .I1(VCC_net), .CO(n39809));
    SB_DFFESR delay_counter_i0_i17 (.Q(delay_counter[17]), .C(CLK_c), .E(n5722), 
            .D(n673), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY encoder0_position_31__I_0_add_1704_7 (.CI(n40085), .I0(n2529), 
            .I1(GND_net), .CO(n40086));
    SB_LUT4 encoder0_position_31__I_0_add_1704_6_lut (.I0(GND_net), .I1(n2530), 
            .I2(GND_net), .I3(n40084), .O(n2597)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1781_3_lut (.I0(n2618), .I1(n2685), 
            .I2(n2643), .I3(GND_net), .O(n2717));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1781_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_673_2 (.CI(VCC_net), .I0(n51409), .I1(n25), .CO(n39279));
    SB_LUT4 encoder0_position_31__I_0_i1795_3_lut (.I0(n2632), .I1(n2699), 
            .I2(n2643), .I3(GND_net), .O(n2731));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1795_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1890_4 (.CI(n39377), .I0(n516), .I1(GND_net), .CO(n39378));
    SB_LUT4 encoder0_position_31__I_0_i1794_3_lut (.I0(n2631), .I1(n2698), 
            .I2(n2643), .I3(GND_net), .O(n2730));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1794_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1793_3_lut (.I0(n2630), .I1(n2697), 
            .I2(n2643), .I3(GND_net), .O(n2729));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1793_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1436_9_lut (.I0(GND_net), .I1(n2127), 
            .I2(VCC_net), .I3(n39807), .O(n2194)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1790_3_lut (.I0(n2627), .I1(n2694), 
            .I2(n2643), .I3(GND_net), .O(n2726));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1790_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1791_3_lut (.I0(n2628), .I1(n2695), 
            .I2(n2643), .I3(GND_net), .O(n2727));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1791_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 add_1890_3_lut (.I0(GND_net), .I1(n625), .I2(VCC_net), .I3(n39376), 
            .O(n6538)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1890_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1797_3_lut (.I0(n951), .I1(n2701), 
            .I2(n2643), .I3(GND_net), .O(n2733));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1797_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1704_6 (.CI(n40084), .I0(n2530), 
            .I1(GND_net), .CO(n40085));
    SB_LUT4 encoder0_position_31__I_0_i1796_3_lut (.I0(n2633), .I1(n2700), 
            .I2(n2643), .I3(GND_net), .O(n2732));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1796_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1436_9 (.CI(n39807), .I0(n2127), 
            .I1(VCC_net), .CO(n39808));
    SB_LUT4 encoder0_position_31__I_0_add_1503_21_lut (.I0(GND_net), .I1(n2215), 
            .I2(VCC_net), .I3(n39919), .O(n2282)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_21_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i16 (.Q(delay_counter[16]), .C(CLK_c), .E(n5722), 
            .D(n674), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY encoder0_position_31__I_0_add_1503_21 (.CI(n39919), .I0(n2215), 
            .I1(VCC_net), .CO(n39920));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i7_3_lut (.I0(encoder0_position[6]), 
            .I1(n27), .I2(encoder0_position[31]), .I3(GND_net), .O(n952));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n5722), 
            .D(n675), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY add_29_2 (.CI(VCC_net), .I0(delay_counter[0]), .I1(GND_net), 
            .CO(n38990));
    SB_CARRY encoder0_position_31__I_0_add_1034_6 (.CI(n39701), .I0(n1530), 
            .I1(GND_net), .CO(n39702));
    SB_LUT4 encoder0_position_31__I_0_add_1704_5_lut (.I0(GND_net), .I1(n2531), 
            .I2(VCC_net), .I3(n40083), .O(n2598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n5722), 
            .D(n676), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_add_1503_20_lut (.I0(GND_net), .I1(n2216), 
            .I2(VCC_net), .I3(n39918), .O(n2283)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_20 (.CI(n39918), .I0(n2216), 
            .I1(VCC_net), .CO(n39919));
    SB_LUT4 encoder0_position_31__I_0_add_1436_8_lut (.I0(GND_net), .I1(n2128), 
            .I2(VCC_net), .I3(n39806), .O(n2195)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1792_rep_17_3_lut (.I0(n2629), .I1(n2696), 
            .I2(n2643), .I3(GND_net), .O(n2728));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1792_rep_17_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1503_19_lut (.I0(GND_net), .I1(n2217), 
            .I2(VCC_net), .I3(n39917), .O(n2284)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1034_5_lut (.I0(GND_net), .I1(n1531), 
            .I2(VCC_net), .I3(n39700), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_8 (.CI(n39806), .I0(n2128), 
            .I1(VCC_net), .CO(n39807));
    SB_CARRY encoder0_position_31__I_0_add_1704_5 (.CI(n40083), .I0(n2531), 
            .I1(VCC_net), .CO(n40084));
    SB_LUT4 encoder0_position_31__I_0_add_1704_4_lut (.I0(GND_net), .I1(n2532), 
            .I2(GND_net), .I3(n40082), .O(n2599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_4 (.CI(n40082), .I0(n2532), 
            .I1(GND_net), .CO(n40083));
    SB_LUT4 encoder0_position_31__I_0_add_1704_3_lut (.I0(GND_net), .I1(n2533), 
            .I2(VCC_net), .I3(n40081), .O(n2600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1704_3 (.CI(n40081), .I0(n2533), 
            .I1(VCC_net), .CO(n40082));
    SB_LUT4 encoder0_position_31__I_0_add_1704_2_lut (.I0(GND_net), .I1(n950), 
            .I2(GND_net), .I3(VCC_net), .O(n2601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1704_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n5722), 
            .D(n677), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_CARRY encoder0_position_31__I_0_add_1704_2 (.CI(VCC_net), .I0(n950), 
            .I1(GND_net), .CO(n40081));
    SB_CARRY add_29_6 (.CI(n38993), .I0(delay_counter[4]), .I1(GND_net), 
            .CO(n38994));
    SB_LUT4 encoder0_position_31__I_0_add_1436_7_lut (.I0(GND_net), .I1(n2129), 
            .I2(GND_net), .I3(n39805), .O(n2196)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_7_lut.LUT_INIT = 16'hC33C;
    \quadrature_decoder(1,500000)_U0  quad_counter0 (.b_prev(b_prev), .GND_net(GND_net), 
            .a_new({a_new[1], Open_0}), .direction_N_3807(direction_N_3807), 
            .ENCODER0_B_N_keep(ENCODER0_B_N), .n1188(CLK_c), .ENCODER0_A_N_keep(ENCODER0_A_N), 
            .encoder0_position({encoder0_position}), .VCC_net(VCC_net), 
            .n28241(n28241), .n1152(n1152)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(187[57] 194[6])
    SB_LUT4 encoder0_position_31__I_0_i1109_3_lut (.I0(n1626), .I1(n1693), 
            .I2(n1653), .I3(GND_net), .O(n1725));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1109_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1788_3_lut (.I0(n2625), .I1(n2692), 
            .I2(n2643), .I3(GND_net), .O(n2724));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1788_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_24_lut (.I0(n51356), .I1(n2412), 
            .I2(VCC_net), .I3(n40080), .O(n2511)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1637_23_lut (.I0(GND_net), .I1(n2413), 
            .I2(VCC_net), .I3(n40079), .O(n2480)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_19 (.CI(n39917), .I0(n2217), 
            .I1(VCC_net), .CO(n39918));
    SB_CARRY encoder0_position_31__I_0_add_1637_23 (.CI(n40079), .I0(n2413), 
            .I1(VCC_net), .CO(n40080));
    SB_LUT4 encoder0_position_31__I_0_i1789_3_lut (.I0(n2626), .I1(n2693), 
            .I2(n2643), .I3(GND_net), .O(n2725));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1789_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1637_22_lut (.I0(GND_net), .I1(n2414), 
            .I2(VCC_net), .I3(n40078), .O(n2481)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_22 (.CI(n40078), .I0(n2414), 
            .I1(VCC_net), .CO(n40079));
    SB_LUT4 encoder0_position_31__I_0_add_1637_21_lut (.I0(GND_net), .I1(n2415), 
            .I2(VCC_net), .I3(n40077), .O(n2482_adj_4959)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1436_7 (.CI(n39805), .I0(n2129), 
            .I1(GND_net), .CO(n39806));
    SB_CARRY encoder0_position_31__I_0_add_1637_21 (.CI(n40077), .I0(n2415), 
            .I1(VCC_net), .CO(n40078));
    SB_LUT4 encoder0_position_31__I_0_i1784_3_lut (.I0(n2621), .I1(n2688), 
            .I2(n2643), .I3(GND_net), .O(n2720));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1784_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1787_3_lut (.I0(n2624), .I1(n2691), 
            .I2(n2643), .I3(GND_net), .O(n2723));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1787_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1034_5 (.CI(n39700), .I0(n1531), 
            .I1(VCC_net), .CO(n39701));
    SB_LUT4 encoder0_position_31__I_0_add_1436_6_lut (.I0(GND_net), .I1(n2130), 
            .I2(GND_net), .I3(n39804), .O(n2197)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i21542_3_lut (.I0(n952), .I1(n2732), .I2(n2733), .I3(GND_net), 
            .O(n34607));
    defparam i21542_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_3_lut_adj_1764 (.I0(n2723), .I1(n2720), .I2(n2725), .I3(GND_net), 
            .O(n47179));
    defparam i1_3_lut_adj_1764.LUT_INIT = 16'hfefe;
    SB_LUT4 encoder0_position_31__I_0_add_1503_18_lut (.I0(GND_net), .I1(n2218), 
            .I2(VCC_net), .I3(n39916), .O(n2285)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1765 (.I0(n2724), .I1(n2722), .I2(n2721), .I3(n2728), 
            .O(n47181));
    defparam i1_4_lut_adj_1765.LUT_INIT = 16'hfffe;
    SB_CARRY add_1890_3 (.CI(n39376), .I0(n625), .I1(VCC_net), .CO(n39377));
    SB_LUT4 i1_4_lut_adj_1766 (.I0(n47181), .I1(n47179), .I2(n2727), .I3(n2726), 
            .O(n47185));
    defparam i1_4_lut_adj_1766.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1767 (.I0(n2729), .I1(n34607), .I2(n2730), .I3(n2731), 
            .O(n45111));
    defparam i1_4_lut_adj_1767.LUT_INIT = 16'ha080;
    SB_CARRY encoder0_position_31__I_0_add_1436_6 (.CI(n39804), .I0(n2130), 
            .I1(GND_net), .CO(n39805));
    SB_LUT4 encoder0_position_31__I_0_add_1034_4_lut (.I0(GND_net), .I1(n1532), 
            .I2(GND_net), .I3(n39699), .O(n1599)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_18 (.CI(n39916), .I0(n2218), 
            .I1(VCC_net), .CO(n39917));
    SB_LUT4 encoder0_position_31__I_0_add_1503_17_lut (.I0(GND_net), .I1(n2219), 
            .I2(VCC_net), .I3(n39915), .O(n2286)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1637_20_lut (.I0(GND_net), .I1(n2416), 
            .I2(VCC_net), .I3(n40076), .O(n2483)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_17 (.CI(n39915), .I0(n2219), 
            .I1(VCC_net), .CO(n39916));
    SB_CARRY encoder0_position_31__I_0_add_1637_20 (.CI(n40076), .I0(n2416), 
            .I1(VCC_net), .CO(n40077));
    SB_CARRY add_29_16 (.CI(n39003), .I0(delay_counter[14]), .I1(GND_net), 
            .CO(n39004));
    SB_LUT4 encoder0_position_31__I_0_add_1637_19_lut (.I0(GND_net), .I1(n2417), 
            .I2(VCC_net), .I3(n40075), .O(n2484)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_19 (.CI(n40075), .I0(n2417), 
            .I1(VCC_net), .CO(n40076));
    SB_LUT4 i1_4_lut_adj_1768 (.I0(n2717), .I1(n2718), .I2(n47185), .I3(n2719), 
            .O(n47191));
    defparam i1_4_lut_adj_1768.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1637_18_lut (.I0(GND_net), .I1(n2418), 
            .I2(VCC_net), .I3(n40074), .O(n2485)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_18 (.CI(n40074), .I0(n2418), 
            .I1(VCC_net), .CO(n40075));
    SB_LUT4 i1_4_lut_adj_1769 (.I0(n2715), .I1(n2716), .I2(n47191), .I3(n45111), 
            .O(n47197));
    defparam i1_4_lut_adj_1769.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1637_17_lut (.I0(GND_net), .I1(n2419), 
            .I2(VCC_net), .I3(n40073), .O(n2486)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_17 (.CI(n40073), .I0(n2419), 
            .I1(VCC_net), .CO(n40074));
    SB_LUT4 encoder0_position_31__I_0_add_1637_16_lut (.I0(GND_net), .I1(n2420), 
            .I2(VCC_net), .I3(n40072), .O(n2487)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_16 (.CI(n40072), .I0(n2420), 
            .I1(VCC_net), .CO(n40073));
    SB_LUT4 encoder0_position_31__I_0_add_1637_15_lut (.I0(GND_net), .I1(n2421), 
            .I2(VCC_net), .I3(n40071), .O(n2488)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_15 (.CI(n40071), .I0(n2421), 
            .I1(VCC_net), .CO(n40072));
    SB_LUT4 i1_4_lut_adj_1770 (.I0(n2712), .I1(n2713), .I2(n2714), .I3(n47197), 
            .O(n47203));
    defparam i1_4_lut_adj_1770.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1637_14_lut (.I0(GND_net), .I1(n2422), 
            .I2(VCC_net), .I3(n40070), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_14 (.CI(n40070), .I0(n2422), 
            .I1(VCC_net), .CO(n40071));
    SB_LUT4 encoder0_position_31__I_0_add_1637_13_lut (.I0(GND_net), .I1(n2423), 
            .I2(VCC_net), .I3(n40069), .O(n2490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_4 (.CI(n39699), .I0(n1532), 
            .I1(GND_net), .CO(n39700));
    SB_LUT4 i36157_4_lut (.I0(n2710), .I1(n2709), .I2(n2711), .I3(n47203), 
            .O(n2742));
    defparam i36157_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1708_3_lut (.I0(n2513), .I1(n2580), 
            .I2(n2544), .I3(GND_net), .O(n2612));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1707_3_lut (.I0(n2512), .I1(n2579), 
            .I2(n2544), .I3(GND_net), .O(n2611));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1711_3_lut (.I0(n2516), .I1(n2583), 
            .I2(n2544), .I3(GND_net), .O(n2615));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1711_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i639_3_lut (.I0(n932), .I1(n999), 
            .I2(n960), .I3(GND_net), .O(n1031));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i639_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1710_3_lut (.I0(n2515), .I1(n2582), 
            .I2(n2544), .I3(GND_net), .O(n2614));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1710_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1709_3_lut (.I0(n2514), .I1(n2581), 
            .I2(n2544), .I3(GND_net), .O(n2613));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1713_3_lut (.I0(n2518), .I1(n2585), 
            .I2(n2544), .I3(GND_net), .O(n2617));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1713_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1637_13 (.CI(n40069), .I0(n2423), 
            .I1(VCC_net), .CO(n40070));
    SB_LUT4 encoder0_position_31__I_0_add_1637_12_lut (.I0(GND_net), .I1(n2424), 
            .I2(VCC_net), .I3(n40068), .O(n2491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_12 (.CI(n40068), .I0(n2424), 
            .I1(VCC_net), .CO(n40069));
    SB_LUT4 encoder0_position_31__I_0_add_1637_11_lut (.I0(GND_net), .I1(n2425), 
            .I2(VCC_net), .I3(n40067), .O(n2492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_11 (.CI(n40067), .I0(n2425), 
            .I1(VCC_net), .CO(n40068));
    SB_LUT4 encoder0_position_31__I_0_add_1637_10_lut (.I0(GND_net), .I1(n2426), 
            .I2(VCC_net), .I3(n40066), .O(n2493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_10 (.CI(n40066), .I0(n2426), 
            .I1(VCC_net), .CO(n40067));
    SB_LUT4 encoder0_position_31__I_0_add_1637_9_lut (.I0(GND_net), .I1(n2427), 
            .I2(VCC_net), .I3(n40065), .O(n2494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_9 (.CI(n40065), .I0(n2427), 
            .I1(VCC_net), .CO(n40066));
    SB_LUT4 encoder0_position_31__I_0_add_1637_8_lut (.I0(GND_net), .I1(n2428), 
            .I2(VCC_net), .I3(n40064), .O(n2495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_8 (.CI(n40064), .I0(n2428), 
            .I1(VCC_net), .CO(n40065));
    SB_LUT4 encoder0_position_31__I_0_add_1637_7_lut (.I0(GND_net), .I1(n2429), 
            .I2(GND_net), .I3(n40063), .O(n2496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_7 (.CI(n40063), .I0(n2429), 
            .I1(GND_net), .CO(n40064));
    SB_LUT4 encoder0_position_31__I_0_add_1637_6_lut (.I0(GND_net), .I1(n2430), 
            .I2(GND_net), .I3(n40062), .O(n2497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_6 (.CI(n40062), .I0(n2430), 
            .I1(GND_net), .CO(n40063));
    SB_LUT4 encoder0_position_31__I_0_add_1637_5_lut (.I0(GND_net), .I1(n2431), 
            .I2(VCC_net), .I3(n40061), .O(n2498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_5 (.CI(n40061), .I0(n2431), 
            .I1(VCC_net), .CO(n40062));
    SB_LUT4 encoder0_position_31__I_0_add_1637_4_lut (.I0(GND_net), .I1(n2432), 
            .I2(GND_net), .I3(n40060), .O(n2499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_4 (.CI(n40060), .I0(n2432), 
            .I1(GND_net), .CO(n40061));
    SB_LUT4 encoder0_position_31__I_0_add_1637_3_lut (.I0(GND_net), .I1(n2433), 
            .I2(VCC_net), .I3(n40059), .O(n2500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_3 (.CI(n40059), .I0(n2433), 
            .I1(VCC_net), .CO(n40060));
    SB_LUT4 encoder0_position_31__I_0_add_1637_2_lut (.I0(GND_net), .I1(n949), 
            .I2(GND_net), .I3(VCC_net), .O(n2501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1637_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1637_2 (.CI(VCC_net), .I0(n949), 
            .I1(GND_net), .CO(n40059));
    SB_LUT4 encoder0_position_31__I_0_add_1570_23_lut (.I0(n51327), .I1(n2313), 
            .I2(VCC_net), .I3(n40058), .O(n2412)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1570_22_lut (.I0(GND_net), .I1(n2314), 
            .I2(VCC_net), .I3(n40057), .O(n2381)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_22 (.CI(n40057), .I0(n2314), 
            .I1(VCC_net), .CO(n40058));
    SB_LUT4 encoder0_position_31__I_0_i1712_3_lut (.I0(n2517), .I1(n2584), 
            .I2(n2544), .I3(GND_net), .O(n2616));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1712_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1570_21_lut (.I0(GND_net), .I1(n2315), 
            .I2(VCC_net), .I3(n40056), .O(n2382)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_21 (.CI(n40056), .I0(n2315), 
            .I1(VCC_net), .CO(n40057));
    SB_LUT4 encoder0_position_31__I_0_add_1570_20_lut (.I0(GND_net), .I1(n2316), 
            .I2(VCC_net), .I3(n40055), .O(n2383)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_20 (.CI(n40055), .I0(n2316), 
            .I1(VCC_net), .CO(n40056));
    SB_LUT4 encoder0_position_31__I_0_i1722_rep_20_3_lut (.I0(n2527), .I1(n2594), 
            .I2(n2544), .I3(GND_net), .O(n2626));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1722_rep_20_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1717_rep_25_3_lut (.I0(n2522), .I1(n2589), 
            .I2(n2544), .I3(GND_net), .O(n2621));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1717_rep_25_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1570_19_lut (.I0(GND_net), .I1(n2317), 
            .I2(VCC_net), .I3(n40054), .O(n2384)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1720_rep_24_3_lut (.I0(n2525), .I1(n2592), 
            .I2(n2544), .I3(GND_net), .O(n2624));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1720_rep_24_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1570_19 (.CI(n40054), .I0(n2317), 
            .I1(VCC_net), .CO(n40055));
    SB_LUT4 encoder0_position_31__I_0_i1724_rep_21_3_lut (.I0(n2529), .I1(n2596), 
            .I2(n2544), .I3(GND_net), .O(n2628));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1724_rep_21_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1729_3_lut (.I0(n950), .I1(n2601), 
            .I2(n2544), .I3(GND_net), .O(n2633));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1729_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1570_18_lut (.I0(GND_net), .I1(n2318), 
            .I2(VCC_net), .I3(n40053), .O(n2385)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1728_3_lut (.I0(n2533), .I1(n2600), 
            .I2(n2544), .I3(GND_net), .O(n2632));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1728_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1570_18 (.CI(n40053), .I0(n2318), 
            .I1(VCC_net), .CO(n40054));
    SB_LUT4 encoder0_position_31__I_0_add_1570_17_lut (.I0(GND_net), .I1(n2319), 
            .I2(VCC_net), .I3(n40052), .O(n2386)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1436_5_lut (.I0(GND_net), .I1(n2131), 
            .I2(VCC_net), .I3(n39803), .O(n2198)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1034_3_lut (.I0(GND_net), .I1(n1533), 
            .I2(VCC_net), .I3(n39698), .O(n1600)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_3 (.CI(n39698), .I0(n1533), 
            .I1(VCC_net), .CO(n39699));
    SB_CARRY encoder0_position_31__I_0_add_1436_5 (.CI(n39803), .I0(n2131), 
            .I1(VCC_net), .CO(n39804));
    SB_LUT4 add_1890_2_lut (.I0(GND_net), .I1(n731), .I2(GND_net), .I3(VCC_net), 
            .O(n6539)) /* synthesis syn_instantiated=1 */ ;
    defparam add_1890_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_17 (.CI(n40052), .I0(n2319), 
            .I1(VCC_net), .CO(n40053));
    SB_LUT4 encoder0_position_31__I_0_mux_3_i8_3_lut (.I0(encoder0_position[7]), 
            .I1(n26), .I2(encoder0_position[31]), .I3(GND_net), .O(n951));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1436_4_lut (.I0(GND_net), .I1(n2132), 
            .I2(GND_net), .I3(n39802), .O(n2199)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_16_lut (.I0(GND_net), .I1(n2320), 
            .I2(VCC_net), .I3(n40051), .O(n2387)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_16_lut (.I0(GND_net), .I1(n2220), 
            .I2(VCC_net), .I3(n39914), .O(n2287)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1716_3_lut (.I0(n2521), .I1(n2588), 
            .I2(n2544), .I3(GND_net), .O(n2620));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1716_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1715_3_lut (.I0(n2520), .I1(n2587), 
            .I2(n2544), .I3(GND_net), .O(n2619));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1715_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1714_3_lut (.I0(n2519), .I1(n2586), 
            .I2(n2544), .I3(GND_net), .O(n2618));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1714_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1727_3_lut (.I0(n2532), .I1(n2599), 
            .I2(n2544), .I3(GND_net), .O(n2631));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1727_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY add_1890_2 (.CI(VCC_net), .I0(n731), .I1(GND_net), .CO(n39376));
    SB_LUT4 encoder0_position_31__I_0_i1726_3_lut (.I0(n2531), .I1(n2598), 
            .I2(n2544), .I3(GND_net), .O(n2630));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1726_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1725_3_lut (.I0(n2530), .I1(n2597), 
            .I2(n2544), .I3(GND_net), .O(n2629));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1725_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1503_16 (.CI(n39914), .I0(n2220), 
            .I1(VCC_net), .CO(n39915));
    SB_LUT4 LessThan_699_i6_3_lut_3_lut (.I0(pwm_setpoint[2]), .I1(pwm_setpoint[3]), 
            .I2(pwm_counter[3]), .I3(GND_net), .O(n6_adj_4963));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i6_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY encoder0_position_31__I_0_add_1436_4 (.CI(n39802), .I0(n2132), 
            .I1(GND_net), .CO(n39803));
    SB_LUT4 encoder0_position_31__I_0_add_1436_3_lut (.I0(GND_net), .I1(n2133), 
            .I2(VCC_net), .I3(n39801), .O(n2200)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1719_3_lut (.I0(n2524), .I1(n2591), 
            .I2(n2544), .I3(GND_net), .O(n2623));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1719_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1723_rep_29_3_lut (.I0(n2528), .I1(n2595), 
            .I2(n2544), .I3(GND_net), .O(n2627));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1723_rep_29_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1436_3 (.CI(n39801), .I0(n2133), 
            .I1(VCC_net), .CO(n39802));
    SB_LUT4 encoder0_position_31__I_0_add_1503_15_lut (.I0(GND_net), .I1(n2221), 
            .I2(VCC_net), .I3(n39913), .O(n2288)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1718_3_lut (.I0(n2523), .I1(n2590), 
            .I2(n2544), .I3(GND_net), .O(n2622));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1718_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1034_2_lut (.I0(GND_net), .I1(n940), 
            .I2(GND_net), .I3(VCC_net), .O(n1601)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1034_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1034_2 (.CI(VCC_net), .I0(n940), 
            .I1(GND_net), .CO(n39698));
    SB_LUT4 encoder0_position_31__I_0_add_967_14_lut (.I0(n50904), .I1(n1422), 
            .I2(VCC_net), .I3(n39697), .O(n1521)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1436_2_lut (.I0(GND_net), .I1(n946), 
            .I2(GND_net), .I3(VCC_net), .O(n2201)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1436_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_15 (.CI(n39913), .I0(n2221), 
            .I1(VCC_net), .CO(n39914));
    SB_CARRY encoder0_position_31__I_0_add_1570_16 (.CI(n40051), .I0(n2320), 
            .I1(VCC_net), .CO(n40052));
    SB_LUT4 encoder0_position_31__I_0_add_1570_15_lut (.I0(GND_net), .I1(n2321), 
            .I2(VCC_net), .I3(n40050), .O(n2388)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_13_lut (.I0(GND_net), .I1(n1423), 
            .I2(VCC_net), .I3(n39696), .O(n1490)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1721_3_lut (.I0(n2526), .I1(n2593), 
            .I2(n2544), .I3(GND_net), .O(n2625));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1721_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_967_13 (.CI(n39696), .I0(n1423), 
            .I1(VCC_net), .CO(n39697));
    SB_CARRY encoder0_position_31__I_0_add_1436_2 (.CI(VCC_net), .I0(n946), 
            .I1(GND_net), .CO(n39801));
    SB_LUT4 encoder0_position_31__I_0_add_1369_20_lut (.I0(n51045), .I1(n2016), 
            .I2(VCC_net), .I3(n39800), .O(n2115)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i21546_3_lut (.I0(n951), .I1(n2632), .I2(n2633), .I3(GND_net), 
            .O(n34611));
    defparam i21546_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_31__I_0_add_1503_14_lut (.I0(GND_net), .I1(n2222), 
            .I2(VCC_net), .I3(n39912), .O(n2289)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_12_lut (.I0(GND_net), .I1(n1424), 
            .I2(VCC_net), .I3(n39695), .O(n1491)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_12 (.CI(n39695), .I0(n1424), 
            .I1(VCC_net), .CO(n39696));
    SB_LUT4 encoder0_position_31__I_0_add_967_11_lut (.I0(GND_net), .I1(n1425), 
            .I2(VCC_net), .I3(n39694), .O(n1492)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_14 (.CI(n39912), .I0(n2222), 
            .I1(VCC_net), .CO(n39913));
    SB_CARRY encoder0_position_31__I_0_add_967_11 (.CI(n39694), .I0(n1425), 
            .I1(VCC_net), .CO(n39695));
    SB_LUT4 encoder0_position_31__I_0_add_1369_19_lut (.I0(GND_net), .I1(n2017), 
            .I2(VCC_net), .I3(n39799), .O(n2084)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_13_lut (.I0(GND_net), .I1(n2223), 
            .I2(VCC_net), .I3(n39911), .O(n2290)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_15 (.CI(n40050), .I0(n2321), 
            .I1(VCC_net), .CO(n40051));
    SB_LUT4 encoder0_position_31__I_0_add_967_10_lut (.I0(GND_net), .I1(n1426), 
            .I2(VCC_net), .I3(n39693), .O(n1493)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_19 (.CI(n39799), .I0(n2017), 
            .I1(VCC_net), .CO(n39800));
    SB_CARRY encoder0_position_31__I_0_add_1503_13 (.CI(n39911), .I0(n2223), 
            .I1(VCC_net), .CO(n39912));
    SB_LUT4 i1_2_lut_adj_1771 (.I0(n2628), .I1(n2624), .I2(GND_net), .I3(GND_net), 
            .O(n47411));
    defparam i1_2_lut_adj_1771.LUT_INIT = 16'heeee;
    SB_LUT4 encoder0_position_31__I_0_add_1503_12_lut (.I0(GND_net), .I1(n2224), 
            .I2(VCC_net), .I3(n39910), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_10 (.CI(n39693), .I0(n1426), 
            .I1(VCC_net), .CO(n39694));
    SB_LUT4 i1_4_lut_adj_1772 (.I0(n2625), .I1(n2622), .I2(n2627), .I3(n2623), 
            .O(n47415));
    defparam i1_4_lut_adj_1772.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1503_12 (.CI(n39910), .I0(n2224), 
            .I1(VCC_net), .CO(n39911));
    SB_LUT4 i1_4_lut_adj_1773 (.I0(n2621), .I1(n47415), .I2(n47411), .I3(n2626), 
            .O(n47419));
    defparam i1_4_lut_adj_1773.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1369_18_lut (.I0(GND_net), .I1(n2018), 
            .I2(VCC_net), .I3(n39798), .O(n2085)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_9_lut (.I0(GND_net), .I1(n1427), 
            .I2(VCC_net), .I3(n39692), .O(n1494)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1774 (.I0(n2629), .I1(n34611), .I2(n2630), .I3(n2631), 
            .O(n45146));
    defparam i1_4_lut_adj_1774.LUT_INIT = 16'ha080;
    SB_CARRY encoder0_position_31__I_0_add_1369_18 (.CI(n39798), .I0(n2018), 
            .I1(VCC_net), .CO(n39799));
    SB_LUT4 encoder0_position_31__I_0_add_1369_17_lut (.I0(GND_net), .I1(n2019), 
            .I2(VCC_net), .I3(n39797), .O(n2086)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_9 (.CI(n39692), .I0(n1427), 
            .I1(VCC_net), .CO(n39693));
    SB_LUT4 encoder0_position_31__I_0_add_967_8_lut (.I0(GND_net), .I1(n1428), 
            .I2(VCC_net), .I3(n39691), .O(n1495)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_17 (.CI(n39797), .I0(n2019), 
            .I1(VCC_net), .CO(n39798));
    SB_LUT4 encoder0_position_31__I_0_add_1503_11_lut (.I0(GND_net), .I1(n2225), 
            .I2(VCC_net), .I3(n39909), .O(n2292)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_14_lut (.I0(GND_net), .I1(n2322), 
            .I2(VCC_net), .I3(n40049), .O(n2389)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_8 (.CI(n39691), .I0(n1428), 
            .I1(VCC_net), .CO(n39692));
    SB_CARRY encoder0_position_31__I_0_add_1570_14 (.CI(n40049), .I0(n2322), 
            .I1(VCC_net), .CO(n40050));
    SB_LUT4 encoder0_position_31__I_0_add_1369_16_lut (.I0(GND_net), .I1(n2020), 
            .I2(VCC_net), .I3(n39796), .O(n2087)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_11 (.CI(n39909), .I0(n2225), 
            .I1(VCC_net), .CO(n39910));
    SB_LUT4 encoder0_position_31__I_0_add_1503_10_lut (.I0(GND_net), .I1(n2226), 
            .I2(VCC_net), .I3(n39908), .O(n2293)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_13_lut (.I0(GND_net), .I1(n2323), 
            .I2(VCC_net), .I3(n40048), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_10 (.CI(n39908), .I0(n2226), 
            .I1(VCC_net), .CO(n39909));
    SB_LUT4 add_29_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(GND_net), 
            .I3(n39002), .O(n677)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_7_lut (.I0(GND_net), .I1(n1429), 
            .I2(GND_net), .I3(n39690), .O(n1496)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_16 (.CI(n39796), .I0(n2020), 
            .I1(VCC_net), .CO(n39797));
    SB_LUT4 encoder0_position_31__I_0_add_1369_15_lut (.I0(GND_net), .I1(n2021), 
            .I2(VCC_net), .I3(n39795), .O(n2088)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_15 (.CI(n39795), .I0(n2021), 
            .I1(VCC_net), .CO(n39796));
    SB_LUT4 encoder0_position_31__I_0_add_1369_14_lut (.I0(GND_net), .I1(n2022), 
            .I2(VCC_net), .I3(n39794), .O(n2089)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_14 (.CI(n39794), .I0(n2022), 
            .I1(VCC_net), .CO(n39795));
    SB_LUT4 encoder0_position_31__I_0_add_1503_9_lut (.I0(GND_net), .I1(n2227), 
            .I2(VCC_net), .I3(n39907), .O(n2294)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1369_13_lut (.I0(GND_net), .I1(n2023), 
            .I2(VCC_net), .I3(n39793), .O(n2090)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_9 (.CI(n39907), .I0(n2227), 
            .I1(VCC_net), .CO(n39908));
    SB_CARRY add_29_15 (.CI(n39002), .I0(delay_counter[13]), .I1(GND_net), 
            .CO(n39003));
    SB_CARRY encoder0_position_31__I_0_add_967_7 (.CI(n39690), .I0(n1429), 
            .I1(GND_net), .CO(n39691));
    SB_LUT4 encoder0_position_31__I_0_add_967_6_lut (.I0(GND_net), .I1(n1430), 
            .I2(GND_net), .I3(n39689), .O(n1497)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_6 (.CI(n39689), .I0(n1430), 
            .I1(GND_net), .CO(n39690));
    SB_LUT4 encoder0_position_31__I_0_add_1503_8_lut (.I0(GND_net), .I1(n2228), 
            .I2(VCC_net), .I3(n39906), .O(n2295)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_5_lut (.I0(GND_net), .I1(n1431), 
            .I2(VCC_net), .I3(n39688), .O(n1498)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_8 (.CI(n39906), .I0(n2228), 
            .I1(VCC_net), .CO(n39907));
    SB_LUT4 encoder0_position_31__I_0_add_1503_7_lut (.I0(GND_net), .I1(n2229), 
            .I2(GND_net), .I3(n39905), .O(n2296)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_7 (.CI(n39905), .I0(n2229), 
            .I1(GND_net), .CO(n39906));
    SB_CARRY encoder0_position_31__I_0_add_1570_13 (.CI(n40048), .I0(n2323), 
            .I1(VCC_net), .CO(n40049));
    SB_LUT4 encoder0_position_31__I_0_add_1570_12_lut (.I0(GND_net), .I1(n2324), 
            .I2(VCC_net), .I3(n40047), .O(n2391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_12 (.CI(n40047), .I0(n2324), 
            .I1(VCC_net), .CO(n40048));
    SB_LUT4 encoder0_position_31__I_0_add_1570_11_lut (.I0(GND_net), .I1(n2325), 
            .I2(VCC_net), .I3(n40046), .O(n2392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_11 (.CI(n40046), .I0(n2325), 
            .I1(VCC_net), .CO(n40047));
    SB_LUT4 i1_4_lut_adj_1775 (.I0(n2618), .I1(n2619), .I2(n2620), .I3(n47419), 
            .O(n47425));
    defparam i1_4_lut_adj_1775.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_add_1570_10_lut (.I0(GND_net), .I1(n2326), 
            .I2(VCC_net), .I3(n40045), .O(n2393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_10 (.CI(n40045), .I0(n2326), 
            .I1(VCC_net), .CO(n40046));
    SB_CARRY encoder0_position_31__I_0_add_1369_13 (.CI(n39793), .I0(n2023), 
            .I1(VCC_net), .CO(n39794));
    SB_LUT4 encoder0_position_31__I_0_add_1570_9_lut (.I0(GND_net), .I1(n2327), 
            .I2(VCC_net), .I3(n40044), .O(n2394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1503_6_lut (.I0(GND_net), .I1(n2230), 
            .I2(GND_net), .I3(n39904), .O(n2297)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1776 (.I0(n2616), .I1(n2617), .I2(n47425), .I3(n45146), 
            .O(n47431));
    defparam i1_4_lut_adj_1776.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1777 (.I0(n2613), .I1(n2614), .I2(n2615), .I3(n47431), 
            .O(n47437));
    defparam i1_4_lut_adj_1777.LUT_INIT = 16'hfffe;
    SB_CARRY encoder0_position_31__I_0_add_1570_9 (.CI(n40044), .I0(n2327), 
            .I1(VCC_net), .CO(n40045));
    SB_LUT4 i35793_4_lut (.I0(n2611), .I1(n2610), .I2(n2612), .I3(n47437), 
            .O(n2643));
    defparam i35793_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_1570_8_lut (.I0(GND_net), .I1(n2328), 
            .I2(VCC_net), .I3(n40043), .O(n2395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_8 (.CI(n40043), .I0(n2328), 
            .I1(VCC_net), .CO(n40044));
    SB_LUT4 encoder0_position_31__I_0_add_1570_7_lut (.I0(GND_net), .I1(n2329), 
            .I2(GND_net), .I3(n40042), .O(n2396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1641_3_lut (.I0(n2414), .I1(n2481), 
            .I2(n2445), .I3(GND_net), .O(n2513));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1641_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1570_7 (.CI(n40042), .I0(n2329), 
            .I1(GND_net), .CO(n40043));
    SB_CARRY encoder0_position_31__I_0_add_1503_6 (.CI(n39904), .I0(n2230), 
            .I1(GND_net), .CO(n39905));
    SB_LUT4 encoder0_position_31__I_0_add_1570_6_lut (.I0(GND_net), .I1(n2330), 
            .I2(GND_net), .I3(n40041), .O(n2397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1640_3_lut (.I0(n2413), .I1(n2480), 
            .I2(n2445), .I3(GND_net), .O(n2512));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1640_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1570_6 (.CI(n40041), .I0(n2330), 
            .I1(GND_net), .CO(n40042));
    SB_LUT4 encoder0_position_31__I_0_add_1570_5_lut (.I0(GND_net), .I1(n2331), 
            .I2(VCC_net), .I3(n40040), .O(n2398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_5 (.CI(n40040), .I0(n2331), 
            .I1(VCC_net), .CO(n40041));
    SB_CARRY encoder0_position_31__I_0_add_967_5 (.CI(n39688), .I0(n1431), 
            .I1(VCC_net), .CO(n39689));
    SB_LUT4 encoder0_position_31__I_0_add_1570_4_lut (.I0(GND_net), .I1(n2332), 
            .I2(GND_net), .I3(n40039), .O(n2399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_967_4_lut (.I0(GND_net), .I1(n1432), 
            .I2(GND_net), .I3(n39687), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_4 (.CI(n40039), .I0(n2332), 
            .I1(GND_net), .CO(n40040));
    SB_LUT4 encoder0_position_31__I_0_add_1570_3_lut (.I0(GND_net), .I1(n2333), 
            .I2(VCC_net), .I3(n40038), .O(n2400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1570_3 (.CI(n40038), .I0(n2333), 
            .I1(VCC_net), .CO(n40039));
    SB_LUT4 encoder0_position_31__I_0_add_1503_5_lut (.I0(GND_net), .I1(n2231), 
            .I2(VCC_net), .I3(n39903), .O(n2298)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1570_2_lut (.I0(GND_net), .I1(n948), 
            .I2(GND_net), .I3(VCC_net), .O(n2401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1570_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1644_3_lut (.I0(n2417), .I1(n2484), 
            .I2(n2445), .I3(GND_net), .O(n2516));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1644_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1570_2 (.CI(VCC_net), .I0(n948), 
            .I1(GND_net), .CO(n40038));
    SB_LUT4 encoder0_position_31__I_0_i1643_3_lut (.I0(n2416), .I1(n2483), 
            .I2(n2445), .I3(GND_net), .O(n2515));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1643_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_967_4 (.CI(n39687), .I0(n1432), 
            .I1(GND_net), .CO(n39688));
    SB_CARRY encoder0_position_31__I_0_add_1503_5 (.CI(n39903), .I0(n2231), 
            .I1(VCC_net), .CO(n39904));
    SB_LUT4 encoder0_position_31__I_0_i1642_3_lut (.I0(n2415), .I1(n2482_adj_4959), 
            .I2(n2445), .I3(GND_net), .O(n2514));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1642_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1661_3_lut (.I0(n949), .I1(n2501), 
            .I2(n2445), .I3(GND_net), .O(n2533));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1661_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1503_4_lut (.I0(GND_net), .I1(n2232), 
            .I2(GND_net), .I3(n39902), .O(n2299)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1660_3_lut (.I0(n2433), .I1(n2500), 
            .I2(n2445), .I3(GND_net), .O(n2532));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1660_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1369_12_lut (.I0(GND_net), .I1(n2024), 
            .I2(VCC_net), .I3(n39792), .O(n2091)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i9_3_lut (.I0(encoder0_position[8]), 
            .I1(n25_adj_4917), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n950));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY encoder0_position_31__I_0_add_1369_12 (.CI(n39792), .I0(n2024), 
            .I1(VCC_net), .CO(n39793));
    SB_LUT4 encoder0_position_31__I_0_add_1369_11_lut (.I0(GND_net), .I1(n2025), 
            .I2(VCC_net), .I3(n39791), .O(n2092)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_11 (.CI(n39791), .I0(n2025), 
            .I1(VCC_net), .CO(n39792));
    SB_LUT4 encoder0_position_31__I_0_add_967_3_lut (.I0(GND_net), .I1(n1433), 
            .I2(VCC_net), .I3(n39686), .O(n1500)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1369_10_lut (.I0(GND_net), .I1(n2026), 
            .I2(VCC_net), .I3(n39790), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_10 (.CI(n39790), .I0(n2026), 
            .I1(VCC_net), .CO(n39791));
    SB_LUT4 encoder0_position_31__I_0_add_1369_9_lut (.I0(GND_net), .I1(n2027), 
            .I2(VCC_net), .I3(n39789), .O(n2094)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_967_3 (.CI(n39686), .I0(n1433), 
            .I1(VCC_net), .CO(n39687));
    SB_LUT4 encoder0_position_31__I_0_add_967_2_lut (.I0(GND_net), .I1(n939), 
            .I2(GND_net), .I3(VCC_net), .O(n1501)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_967_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_9 (.CI(n39789), .I0(n2027), 
            .I1(VCC_net), .CO(n39790));
    SB_LUT4 encoder0_position_31__I_0_i1646_3_lut (.I0(n2419), .I1(n2486), 
            .I2(n2445), .I3(GND_net), .O(n2518));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1646_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1369_8_lut (.I0(GND_net), .I1(n2028), 
            .I2(VCC_net), .I3(n39788), .O(n2095)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1645_3_lut (.I0(n2418), .I1(n2485), 
            .I2(n2445), .I3(GND_net), .O(n2517));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1645_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1656_3_lut (.I0(n2429), .I1(n2496), 
            .I2(n2445), .I3(GND_net), .O(n2528));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1656_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1651_3_lut (.I0(n2424), .I1(n2491), 
            .I2(n2445), .I3(GND_net), .O(n2523));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1651_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1653_3_lut (.I0(n2426), .I1(n2493), 
            .I2(n2445), .I3(GND_net), .O(n2525));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1653_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_967_2 (.CI(VCC_net), .I0(n939), 
            .I1(GND_net), .CO(n39686));
    SB_CARRY encoder0_position_31__I_0_add_1369_8 (.CI(n39788), .I0(n2028), 
            .I1(VCC_net), .CO(n39789));
    SB_DFF h1_56 (.Q(INLA_c), .C(CLK_c), .D(hall1));   // verilog/TinyFPGA_B.v(96[10] 109[6])
    SB_LUT4 encoder0_position_31__I_0_add_900_13_lut (.I0(n50832), .I1(n1323), 
            .I2(VCC_net), .I3(n39685), .O(n1422)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY encoder0_position_31__I_0_add_1503_4 (.CI(n39902), .I0(n2232), 
            .I1(GND_net), .CO(n39903));
    SB_LUT4 encoder0_position_31__I_0_add_1503_3_lut (.I0(GND_net), .I1(n2233), 
            .I2(VCC_net), .I3(n39901), .O(n2300)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_900_12_lut (.I0(GND_net), .I1(n1324), 
            .I2(VCC_net), .I3(n39684), .O(n1391)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1369_7_lut (.I0(GND_net), .I1(n2029), 
            .I2(GND_net), .I3(n39787), .O(n2096)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1503_3 (.CI(n39901), .I0(n2233), 
            .I1(VCC_net), .CO(n39902));
    SB_LUT4 encoder0_position_31__I_0_add_1503_2_lut (.I0(GND_net), .I1(n947), 
            .I2(GND_net), .I3(VCC_net), .O(n2301)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1503_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_7 (.CI(n39787), .I0(n2029), 
            .I1(GND_net), .CO(n39788));
    SB_CARRY encoder0_position_31__I_0_add_1503_2 (.CI(VCC_net), .I0(n947), 
            .I1(GND_net), .CO(n39901));
    SB_CARRY encoder0_position_31__I_0_add_900_12 (.CI(n39684), .I0(n1324), 
            .I1(VCC_net), .CO(n39685));
    SB_LUT4 add_29_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(GND_net), 
            .I3(n39001), .O(n678)) /* synthesis syn_instantiated=1 */ ;
    defparam add_29_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1369_6_lut (.I0(GND_net), .I1(n2030), 
            .I2(GND_net), .I3(n39786), .O(n2097)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_900_11_lut (.I0(GND_net), .I1(n1325), 
            .I2(VCC_net), .I3(n39683), .O(n1392)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_6 (.CI(n39786), .I0(n2030), 
            .I1(GND_net), .CO(n39787));
    SB_CARRY encoder0_position_31__I_0_add_900_11 (.CI(n39683), .I0(n1325), 
            .I1(VCC_net), .CO(n39684));
    SB_LUT4 encoder0_position_31__I_0_i1654_3_lut (.I0(n2427), .I1(n2494), 
            .I2(n2445), .I3(GND_net), .O(n2526));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1654_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1369_5_lut (.I0(GND_net), .I1(n2031), 
            .I2(VCC_net), .I3(n39785), .O(n2098)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1659_3_lut (.I0(n2432), .I1(n2499), 
            .I2(n2445), .I3(GND_net), .O(n2531));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1659_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1658_3_lut (.I0(n2431), .I1(n2498), 
            .I2(n2445), .I3(GND_net), .O(n2530));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1658_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1369_5 (.CI(n39785), .I0(n2031), 
            .I1(VCC_net), .CO(n39786));
    SB_LUT4 encoder0_position_31__I_0_add_1369_4_lut (.I0(GND_net), .I1(n2032), 
            .I2(GND_net), .I3(n39784), .O(n2099)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1657_3_lut (.I0(n2430), .I1(n2497), 
            .I2(n2445), .I3(GND_net), .O(n2529));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1657_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1369_4 (.CI(n39784), .I0(n2032), 
            .I1(GND_net), .CO(n39785));
    SB_LUT4 encoder0_position_31__I_0_add_900_10_lut (.I0(GND_net), .I1(n1326), 
            .I2(VCC_net), .I3(n39682), .O(n1393)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1369_3_lut (.I0(GND_net), .I1(n2033), 
            .I2(VCC_net), .I3(n39783), .O(n2100)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_10 (.CI(n39682), .I0(n1326), 
            .I1(VCC_net), .CO(n39683));
    SB_CARRY encoder0_position_31__I_0_add_1369_3 (.CI(n39783), .I0(n2033), 
            .I1(VCC_net), .CO(n39784));
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n5722), 
            .D(n678), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_i1648_3_lut (.I0(n2421), .I1(n2488), 
            .I2(n2445), .I3(GND_net), .O(n2520));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1648_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_1369_2_lut (.I0(GND_net), .I1(n945), 
            .I2(GND_net), .I3(VCC_net), .O(n2101)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1369_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_900_9_lut (.I0(GND_net), .I1(n1327), 
            .I2(VCC_net), .I3(n39681), .O(n1394)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1369_2 (.CI(VCC_net), .I0(n945), 
            .I1(GND_net), .CO(n39783));
    SB_LUT4 encoder0_position_31__I_0_i1647_3_lut (.I0(n2420), .I1(n2487), 
            .I2(n2445), .I3(GND_net), .O(n2519));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1647_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_900_9 (.CI(n39681), .I0(n1327), 
            .I1(VCC_net), .CO(n39682));
    SB_LUT4 encoder0_position_31__I_0_i1650_3_lut (.I0(n2423), .I1(n2490), 
            .I2(n2445), .I3(GND_net), .O(n2522));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1650_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_900_8_lut (.I0(GND_net), .I1(n1328), 
            .I2(VCC_net), .I3(n39680), .O(n1395)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_1302_19_lut (.I0(n51019), .I1(n1917), 
            .I2(VCC_net), .I3(n39782), .O(n2016)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_add_1302_18_lut (.I0(GND_net), .I1(n1918), 
            .I2(VCC_net), .I3(n39781), .O(n1985)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1655_3_lut (.I0(n2428), .I1(n2495), 
            .I2(n2445), .I3(GND_net), .O(n2527));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1655_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_900_8 (.CI(n39680), .I0(n1328), 
            .I1(VCC_net), .CO(n39681));
    SB_LUT4 encoder0_position_31__I_0_i1652_3_lut (.I0(n2425), .I1(n2492), 
            .I2(n2445), .I3(GND_net), .O(n2524));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1652_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_add_900_7_lut (.I0(GND_net), .I1(n1329), 
            .I2(GND_net), .I3(n39679), .O(n1396)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_18 (.CI(n39781), .I0(n1918), 
            .I1(VCC_net), .CO(n39782));
    SB_LUT4 encoder0_position_31__I_0_i1185_3_lut (.I0(n942), .I1(n1801), 
            .I2(n1752), .I3(GND_net), .O(n1833));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1185_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_900_7 (.CI(n39679), .I0(n1329), 
            .I1(GND_net), .CO(n39680));
    SB_LUT4 encoder0_position_31__I_0_add_1302_17_lut (.I0(GND_net), .I1(n1919), 
            .I2(VCC_net), .I3(n39780), .O(n1986)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_900_6_lut (.I0(GND_net), .I1(n1330), 
            .I2(GND_net), .I3(n39678), .O(n1397)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_17 (.CI(n39780), .I0(n1919), 
            .I1(VCC_net), .CO(n39781));
    SB_CARRY encoder0_position_31__I_0_add_900_6 (.CI(n39678), .I0(n1330), 
            .I1(GND_net), .CO(n39679));
    SB_CARRY add_29_14 (.CI(n39001), .I0(delay_counter[12]), .I1(GND_net), 
            .CO(n39002));
    SB_LUT4 encoder0_position_31__I_0_add_1302_16_lut (.I0(GND_net), .I1(n1920), 
            .I2(VCC_net), .I3(n39779), .O(n1987)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_16 (.CI(n39779), .I0(n1920), 
            .I1(VCC_net), .CO(n39780));
    SB_LUT4 encoder0_position_31__I_0_add_1302_15_lut (.I0(GND_net), .I1(n1921), 
            .I2(VCC_net), .I3(n39778), .O(n1988)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1649_rep_32_3_lut (.I0(n2422), .I1(n2489), 
            .I2(n2445), .I3(GND_net), .O(n2521));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1649_rep_32_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1302_15 (.CI(n39778), .I0(n1921), 
            .I1(VCC_net), .CO(n39779));
    SB_LUT4 encoder0_position_31__I_0_add_1302_14_lut (.I0(GND_net), .I1(n1922), 
            .I2(VCC_net), .I3(n39777), .O(n1989)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_900_5_lut (.I0(GND_net), .I1(n1331), 
            .I2(VCC_net), .I3(n39677), .O(n1398)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_14 (.CI(n39777), .I0(n1922), 
            .I1(VCC_net), .CO(n39778));
    SB_LUT4 encoder0_position_31__I_0_add_1302_13_lut (.I0(GND_net), .I1(n1923), 
            .I2(VCC_net), .I3(n39776), .O(n1990)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_5 (.CI(n39677), .I0(n1331), 
            .I1(VCC_net), .CO(n39678));
    SB_CARRY encoder0_position_31__I_0_add_1302_13 (.CI(n39776), .I0(n1923), 
            .I1(VCC_net), .CO(n39777));
    SB_LUT4 encoder0_position_31__I_0_add_1302_12_lut (.I0(GND_net), .I1(n1924), 
            .I2(VCC_net), .I3(n39775), .O(n1991)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_900_4_lut (.I0(GND_net), .I1(n1332), 
            .I2(GND_net), .I3(n39676), .O(n1399)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_12 (.CI(n39775), .I0(n1924), 
            .I1(VCC_net), .CO(n39776));
    SB_LUT4 i1_4_lut_adj_1778 (.I0(n2526), .I1(n2525), .I2(n2523), .I3(n2528), 
            .O(n47119));
    defparam i1_4_lut_adj_1778.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1184_3_lut (.I0(n1733), .I1(n1800), 
            .I2(n1752), .I3(GND_net), .O(n1832));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1184_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1779 (.I0(n2521), .I1(n2524), .I2(n2527), .I3(n2522), 
            .O(n47121));
    defparam i1_4_lut_adj_1779.LUT_INIT = 16'hfffe;
    SB_LUT4 i21550_3_lut (.I0(n950), .I1(n2532), .I2(n2533), .I3(GND_net), 
            .O(n34615));
    defparam i21550_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1780 (.I0(n2519), .I1(n2520), .I2(n47121), .I3(n47119), 
            .O(n47127));
    defparam i1_4_lut_adj_1780.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1781 (.I0(n2529), .I1(n34615), .I2(n2530), .I3(n2531), 
            .O(n45105));
    defparam i1_4_lut_adj_1781.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1782 (.I0(n2517), .I1(n2518), .I2(n45105), .I3(n47127), 
            .O(n47133));
    defparam i1_4_lut_adj_1782.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1783 (.I0(n2514), .I1(n2515), .I2(n2516), .I3(n47133), 
            .O(n47139));
    defparam i1_4_lut_adj_1783.LUT_INIT = 16'hfffe;
    GND i1 (.Y(GND_net));
    SB_LUT4 encoder0_position_31__I_0_add_1302_11_lut (.I0(GND_net), .I1(n1925), 
            .I2(VCC_net), .I3(n39774), .O(n1992)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_4 (.CI(n39676), .I0(n1332), 
            .I1(GND_net), .CO(n39677));
    SB_LUT4 i36440_4_lut (.I0(n2512), .I1(n2511), .I2(n2513), .I3(n47139), 
            .O(n2544));
    defparam i36440_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_add_900_3_lut (.I0(GND_net), .I1(n1333), 
            .I2(VCC_net), .I3(n39675), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_1302_11 (.CI(n39774), .I0(n1925), 
            .I1(VCC_net), .CO(n39775));
    SB_LUT4 encoder0_position_31__I_0_i1593_rep_33_3_lut (.I0(n948), .I1(n2401), 
            .I2(n2346), .I3(GND_net), .O(n2433));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1593_rep_33_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1592_3_lut (.I0(n2333), .I1(n2400), 
            .I2(n2346), .I3(GND_net), .O(n2432));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1592_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i10_3_lut (.I0(encoder0_position[9]), 
            .I1(n24_adj_4918), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n949));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_add_1302_10_lut (.I0(GND_net), .I1(n1926), 
            .I2(VCC_net), .I3(n39773), .O(n1993)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_i1574_3_lut (.I0(n2315), .I1(n2382), 
            .I2(n2346), .I3(GND_net), .O(n2414));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1574_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1573_3_lut (.I0(n2314), .I1(n2381), 
            .I2(n2346), .I3(GND_net), .O(n2413));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1573_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1577_3_lut (.I0(n2318), .I1(n2385), 
            .I2(n2346), .I3(GND_net), .O(n2417));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1577_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1576_3_lut (.I0(n2317), .I1(n2384), 
            .I2(n2346), .I3(GND_net), .O(n2416));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1576_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1575_3_lut (.I0(n2316), .I1(n2383), 
            .I2(n2346), .I3(GND_net), .O(n2415));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1575_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_1302_10 (.CI(n39773), .I0(n1926), 
            .I1(VCC_net), .CO(n39774));
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n5722), 
            .D(n679), .R(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    SB_LUT4 encoder0_position_31__I_0_i1579_3_lut (.I0(n2320), .I1(n2387), 
            .I2(n2346), .I3(GND_net), .O(n2419));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1579_3_lut.LUT_INIT = 16'hacac;
    SB_CARRY encoder0_position_31__I_0_add_900_3 (.CI(n39675), .I0(n1333), 
            .I1(VCC_net), .CO(n39676));
    SB_LUT4 encoder0_position_31__I_0_add_1302_9_lut (.I0(GND_net), .I1(n1927), 
            .I2(VCC_net), .I3(n39772), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_1302_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 encoder0_position_31__I_0_add_900_2_lut (.I0(GND_net), .I1(n938), 
            .I2(GND_net), .I3(VCC_net), .O(n1401)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_900_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY encoder0_position_31__I_0_add_900_2 (.CI(VCC_net), .I0(n938), 
            .I1(GND_net), .CO(n39675));
    SB_LUT4 encoder0_position_31__I_0_add_833_12_lut (.I0(n50817), .I1(n1224), 
            .I2(VCC_net), .I3(n39674), .O(n1323)) /* synthesis syn_instantiated=1 */ ;
    defparam encoder0_position_31__I_0_add_833_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i16_3_lut (.I0(encoder0_position[15]), 
            .I1(n18_adj_4924), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n943));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1110_3_lut (.I0(n1627), .I1(n1694), 
            .I2(n1653), .I3(GND_net), .O(n1726));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1110_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1578_3_lut (.I0(n2319), .I1(n2386), 
            .I2(n2346), .I3(GND_net), .O(n2418));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1578_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1591_3_lut (.I0(n2332), .I1(n2399), 
            .I2(n2346), .I3(GND_net), .O(n2431));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1591_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1590_3_lut (.I0(n2331), .I1(n2398), 
            .I2(n2346), .I3(GND_net), .O(n2430));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1590_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1589_3_lut (.I0(n2330), .I1(n2397), 
            .I2(n2346), .I3(GND_net), .O(n2429));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1589_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1581_3_lut (.I0(n2322), .I1(n2389), 
            .I2(n2346), .I3(GND_net), .O(n2421));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1581_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1580_3_lut (.I0(n2321), .I1(n2388), 
            .I2(n2346), .I3(GND_net), .O(n2420));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1580_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1583_3_lut (.I0(n2324), .I1(n2391), 
            .I2(n2346), .I3(GND_net), .O(n2423));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1583_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1582_3_lut (.I0(n2323), .I1(n2390), 
            .I2(n2346), .I3(GND_net), .O(n2422));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1582_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1585_3_lut (.I0(n2326), .I1(n2393), 
            .I2(n2346), .I3(GND_net), .O(n2425));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1585_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1588_3_lut (.I0(n2329), .I1(n2396), 
            .I2(n2346), .I3(GND_net), .O(n2428));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1588_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1584_3_lut (.I0(n2325), .I1(n2392), 
            .I2(n2346), .I3(GND_net), .O(n2424));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1584_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1587_3_lut (.I0(n2328), .I1(n2395), 
            .I2(n2346), .I3(GND_net), .O(n2427));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1587_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1586_3_lut (.I0(n2327), .I1(n2394), 
            .I2(n2346), .I3(GND_net), .O(n2426));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1586_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1784 (.I0(n2426), .I1(n2427), .I2(n2424), .I3(n2428), 
            .O(n47379));
    defparam i1_4_lut_adj_1784.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_3_lut_adj_1785 (.I0(n2425), .I1(n2422), .I2(n2423), .I3(GND_net), 
            .O(n47377));
    defparam i1_3_lut_adj_1785.LUT_INIT = 16'hfefe;
    SB_LUT4 i21552_3_lut (.I0(n949), .I1(n2432), .I2(n2433), .I3(GND_net), 
            .O(n34617));
    defparam i21552_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1786 (.I0(n2420), .I1(n2421), .I2(n47377), .I3(n47379), 
            .O(n47385));
    defparam i1_4_lut_adj_1786.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1787 (.I0(n2429), .I1(n34617), .I2(n2430), .I3(n2431), 
            .O(n45131));
    defparam i1_4_lut_adj_1787.LUT_INIT = 16'ha080;
    SB_LUT4 encoder0_position_31__I_0_i638_3_lut (.I0(n931), .I1(n998), 
            .I2(n960), .I3(GND_net), .O(n1030));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i638_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1788 (.I0(n2418), .I1(n2419), .I2(n45131), .I3(n47385), 
            .O(n47391));
    defparam i1_4_lut_adj_1788.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1789 (.I0(n2415), .I1(n2416), .I2(n2417), .I3(n47391), 
            .O(n47397));
    defparam i1_4_lut_adj_1789.LUT_INIT = 16'hfffe;
    SB_LUT4 i36407_4_lut (.I0(n2413), .I1(n2412), .I2(n2414), .I3(n47397), 
            .O(n2445));
    defparam i36407_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 i3_4_lut_adj_1790 (.I0(n74), .I1(n46759), .I2(n771), .I3(n8_adj_5037), 
            .O(n8_adj_5034));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1790.LUT_INIT = 16'hff37;
    SB_LUT4 i2_4_lut_adj_1791 (.I0(\FRAME_MATCHER.i_31__N_2524 ), .I1(\FRAME_MATCHER.i_31__N_2526 ), 
            .I2(n3303), .I3(n4452), .O(n7_adj_5035));   // verilog/coms.v(127[12] 300[6])
    defparam i2_4_lut_adj_1791.LUT_INIT = 16'h0ace;
    SB_LUT4 i2_2_lut (.I0(n33298), .I1(\FRAME_MATCHER.state [3]), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_5026));
    defparam i2_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_4_lut_adj_1792 (.I0(n7_adj_5035), .I1(\FRAME_MATCHER.state [0]), 
            .I2(n8_adj_5034), .I3(n23831), .O(n40_adj_5036));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1792.LUT_INIT = 16'hc8fa;
    SB_LUT4 LessThan_699_i10_3_lut_3_lut (.I0(pwm_setpoint[5]), .I1(pwm_setpoint[6]), 
            .I2(pwm_counter[6]), .I3(GND_net), .O(n10_adj_4967));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i10_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35030_2_lut_4_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[7]), .I3(pwm_setpoint[7]), .O(n49982));
    defparam i35030_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_4_lut_adj_1793 (.I0(\FRAME_MATCHER.state [0]), .I1(n40_adj_5036), 
            .I2(n6_adj_5026), .I3(n73), .O(n43485));   // verilog/coms.v(127[12] 300[6])
    defparam i1_4_lut_adj_1793.LUT_INIT = 16'hcdcc;
    SB_LUT4 LessThan_699_i12_3_lut_3_lut (.I0(pwm_setpoint[7]), .I1(pwm_setpoint[16]), 
            .I2(pwm_counter[16]), .I3(GND_net), .O(n12_adj_4969));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i12_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_31__I_0_i1507_3_lut (.I0(n2216), .I1(n2283), 
            .I2(n2247), .I3(GND_net), .O(n2315));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1507_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1505_3_lut (.I0(n2214), .I1(n2281), 
            .I2(n2247), .I3(GND_net), .O(n2313));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1505_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1506_3_lut (.I0(n2215), .I1(n2282), 
            .I2(n2247), .I3(GND_net), .O(n2314));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1506_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1510_3_lut (.I0(n2219), .I1(n2286), 
            .I2(n2247), .I3(GND_net), .O(n2318));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1510_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1509_3_lut (.I0(n2218), .I1(n2285), 
            .I2(n2247), .I3(GND_net), .O(n2317));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1509_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1508_3_lut (.I0(n2217), .I1(n2284), 
            .I2(n2247), .I3(GND_net), .O(n2316));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1508_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1513_3_lut (.I0(n2222), .I1(n2289), 
            .I2(n2247), .I3(GND_net), .O(n2321));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1513_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1512_3_lut (.I0(n2221), .I1(n2288), 
            .I2(n2247), .I3(GND_net), .O(n2320));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1512_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1511_3_lut (.I0(n2220), .I1(n2287), 
            .I2(n2247), .I3(GND_net), .O(n2319));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1511_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1522_3_lut (.I0(n2231), .I1(n2298), 
            .I2(n2247), .I3(GND_net), .O(n2330));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1522_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1521_3_lut (.I0(n2230), .I1(n2297), 
            .I2(n2247), .I3(GND_net), .O(n2329));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1521_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1525_3_lut (.I0(n947), .I1(n2301), 
            .I2(n2247), .I3(GND_net), .O(n2333));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1525_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1524_3_lut (.I0(n2233), .I1(n2300), 
            .I2(n2247), .I3(GND_net), .O(n2332));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1524_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1523_3_lut (.I0(n2232), .I1(n2299), 
            .I2(n2247), .I3(GND_net), .O(n2331));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1523_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i11_3_lut (.I0(encoder0_position[10]), 
            .I1(n23_adj_4919), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n948));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1518_rep_34_3_lut (.I0(n2227), .I1(n2294), 
            .I2(n2247), .I3(GND_net), .O(n2326));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1518_rep_34_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1514_3_lut (.I0(n2223), .I1(n2290), 
            .I2(n2247), .I3(GND_net), .O(n2322));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1514_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1515_rep_39_3_lut (.I0(n2224), .I1(n2291), 
            .I2(n2247), .I3(GND_net), .O(n2323));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1515_rep_39_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1520_rep_38_3_lut (.I0(n2229), .I1(n2296), 
            .I2(n2247), .I3(GND_net), .O(n2328));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1520_rep_38_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1517_rep_35_3_lut (.I0(n2226), .I1(n2293), 
            .I2(n2247), .I3(GND_net), .O(n2325));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1517_rep_35_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1516_rep_36_3_lut (.I0(n2225), .I1(n2292), 
            .I2(n2247), .I3(GND_net), .O(n2324));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1516_rep_36_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1519_rep_37_3_lut (.I0(n2228), .I1(n2295), 
            .I2(n2247), .I3(GND_net), .O(n2327));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1519_rep_37_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1794 (.I0(n2327), .I1(n2324), .I2(n2325), .I3(n2328), 
            .O(n47017));
    defparam i1_4_lut_adj_1794.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1795 (.I0(n2323), .I1(n47017), .I2(n2322), .I3(n2326), 
            .O(n47019));
    defparam i1_4_lut_adj_1795.LUT_INIT = 16'hfffe;
    SB_LUT4 i21655_4_lut (.I0(n948), .I1(n2331), .I2(n2332), .I3(n2333), 
            .O(n34723));
    defparam i21655_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1796 (.I0(n2319), .I1(n2320), .I2(n2321), .I3(n47019), 
            .O(n47025));
    defparam i1_4_lut_adj_1796.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1797 (.I0(n47025), .I1(n2329), .I2(n34723), .I3(n2330), 
            .O(n47027));
    defparam i1_4_lut_adj_1797.LUT_INIT = 16'heaaa;
    SB_LUT4 i1_4_lut_adj_1798 (.I0(n2316), .I1(n2317), .I2(n2318), .I3(n47027), 
            .O(n47033));
    defparam i1_4_lut_adj_1798.LUT_INIT = 16'hfffe;
    SB_LUT4 i36378_4_lut (.I0(n2314), .I1(n2313), .I2(n2315), .I3(n47033), 
            .O(n2346));
    defparam i36378_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i12_1_lut (.I0(encoder1_position_scaled[11]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n14_adj_4900));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i1439_3_lut (.I0(n2116), .I1(n2183), 
            .I2(n2148), .I3(GND_net), .O(n2215));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1439_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1444_3_lut (.I0(n2121), .I1(n2188), 
            .I2(n2148), .I3(GND_net), .O(n2220));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1444_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1443_3_lut (.I0(n2120), .I1(n2187), 
            .I2(n2148), .I3(GND_net), .O(n2219));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1443_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1451_3_lut (.I0(n2128), .I1(n2195), 
            .I2(n2148), .I3(GND_net), .O(n2227));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1451_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1447_3_lut (.I0(n2124), .I1(n2191), 
            .I2(n2148), .I3(GND_net), .O(n2223));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1447_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1452_3_lut (.I0(n2129), .I1(n2196), 
            .I2(n2148), .I3(GND_net), .O(n2228));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1452_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1445_3_lut (.I0(n2122), .I1(n2189), 
            .I2(n2148), .I3(GND_net), .O(n2221));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1445_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1457_3_lut (.I0(n946), .I1(n2201), 
            .I2(n2148), .I3(GND_net), .O(n2233));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1457_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1456_3_lut (.I0(n2133), .I1(n2200), 
            .I2(n2148), .I3(GND_net), .O(n2232));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1456_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i12_3_lut (.I0(encoder0_position[11]), 
            .I1(n22_adj_4920), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n947));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1442_3_lut (.I0(n2119), .I1(n2186), 
            .I2(n2148), .I3(GND_net), .O(n2218));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1442_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1441_3_lut (.I0(n2118), .I1(n2185), 
            .I2(n2148), .I3(GND_net), .O(n2217));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1441_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1440_3_lut (.I0(n2117), .I1(n2184), 
            .I2(n2148), .I3(GND_net), .O(n2216));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1440_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1455_3_lut (.I0(n2132), .I1(n2199), 
            .I2(n2148), .I3(GND_net), .O(n2231));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1455_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1454_3_lut (.I0(n2131), .I1(n2198), 
            .I2(n2148), .I3(GND_net), .O(n2230));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1454_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1453_3_lut (.I0(n2130), .I1(n2197), 
            .I2(n2148), .I3(GND_net), .O(n2229));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1453_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1449_3_lut (.I0(n2126), .I1(n2193), 
            .I2(n2148), .I3(GND_net), .O(n2225));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1449_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1450_3_lut (.I0(n2127), .I1(n2194), 
            .I2(n2148), .I3(GND_net), .O(n2226));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1450_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1448_3_lut (.I0(n2125), .I1(n2192), 
            .I2(n2148), .I3(GND_net), .O(n2224));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1448_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1446_3_lut (.I0(n2123), .I1(n2190), 
            .I2(n2148), .I3(GND_net), .O(n2222));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1446_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36349_1_lut (.I0(n2247), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51302));
    defparam i36349_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1799 (.I0(n2222), .I1(n2224), .I2(n2226), .I3(n2225), 
            .O(n47357));
    defparam i1_4_lut_adj_1799.LUT_INIT = 16'hfffe;
    SB_LUT4 i21564_3_lut (.I0(n947), .I1(n2232), .I2(n2233), .I3(GND_net), 
            .O(n34631));
    defparam i21564_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1800 (.I0(n2221), .I1(n2228), .I2(n2223), .I3(n2227), 
            .O(n47345));
    defparam i1_4_lut_adj_1800.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1801 (.I0(n2229), .I1(n34631), .I2(n2230), .I3(n2231), 
            .O(n45116));
    defparam i1_4_lut_adj_1801.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1802 (.I0(n2216), .I1(n2217), .I2(n2218), .I3(n47357), 
            .O(n47363));
    defparam i1_4_lut_adj_1802.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1803 (.I0(n2219), .I1(n2220), .I2(n45116), .I3(n47345), 
            .O(n47351));
    defparam i1_4_lut_adj_1803.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1112_3_lut (.I0(n1629), .I1(n1696), 
            .I2(n1653), .I3(GND_net), .O(n1728));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1112_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i36352_4_lut (.I0(n2214), .I1(n47351), .I2(n47363), .I3(n2215), 
            .O(n2247));
    defparam i36352_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1373_3_lut (.I0(n2018), .I1(n2085), 
            .I2(n2049), .I3(GND_net), .O(n2117));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1373_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1372_3_lut (.I0(n2017), .I1(n2084), 
            .I2(n2049), .I3(GND_net), .O(n2116));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1372_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1386_3_lut (.I0(n2031), .I1(n2098), 
            .I2(n2049), .I3(GND_net), .O(n2130));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1386_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1385_3_lut (.I0(n2030), .I1(n2097), 
            .I2(n2049), .I3(GND_net), .O(n2129));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1385_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1376_3_lut (.I0(n2021), .I1(n2088), 
            .I2(n2049), .I3(GND_net), .O(n2120));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1376_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1375_3_lut (.I0(n2020), .I1(n2087), 
            .I2(n2049), .I3(GND_net), .O(n2119));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1375_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1374_3_lut (.I0(n2019), .I1(n2086), 
            .I2(n2049), .I3(GND_net), .O(n2118));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1374_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1382_3_lut (.I0(n2027), .I1(n2094), 
            .I2(n2049), .I3(GND_net), .O(n2126));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1382_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1384_3_lut (.I0(n2029), .I1(n2096), 
            .I2(n2049), .I3(GND_net), .O(n2128));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1384_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1383_3_lut (.I0(n2028), .I1(n2095), 
            .I2(n2049), .I3(GND_net), .O(n2127));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1383_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1381_3_lut (.I0(n2026), .I1(n2093), 
            .I2(n2049), .I3(GND_net), .O(n2125));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1381_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1380_3_lut (.I0(n2025), .I1(n2092), 
            .I2(n2049), .I3(GND_net), .O(n2124));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1380_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1379_3_lut (.I0(n2024), .I1(n2091), 
            .I2(n2049), .I3(GND_net), .O(n2123));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1379_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1378_3_lut (.I0(n2023), .I1(n2090), 
            .I2(n2049), .I3(GND_net), .O(n2122));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1378_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1377_3_lut (.I0(n2022), .I1(n2089), 
            .I2(n2049), .I3(GND_net), .O(n2121));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1377_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1389_rep_40_3_lut (.I0(n945), .I1(n2101), 
            .I2(n2049), .I3(GND_net), .O(n2133));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1389_rep_40_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1388_3_lut (.I0(n2033), .I1(n2100), 
            .I2(n2049), .I3(GND_net), .O(n2132));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1388_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1387_3_lut (.I0(n2032), .I1(n2099), 
            .I2(n2049), .I3(GND_net), .O(n2131));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1387_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i13_3_lut (.I0(encoder0_position[12]), 
            .I1(n21_adj_4921), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n946));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1804 (.I0(n2123), .I1(n2124), .I2(GND_net), .I3(GND_net), 
            .O(n47043));
    defparam i1_2_lut_adj_1804.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1805 (.I0(n2125), .I1(n2127), .I2(n2128), .I3(n2126), 
            .O(n47045));
    defparam i1_4_lut_adj_1805.LUT_INIT = 16'hfffe;
    SB_LUT4 i21667_4_lut (.I0(n946), .I1(n2131), .I2(n2132), .I3(n2133), 
            .O(n34735));
    defparam i21667_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_4_lut_adj_1806 (.I0(n2121), .I1(n2122), .I2(n47045), .I3(n47043), 
            .O(n47051));
    defparam i1_4_lut_adj_1806.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1807 (.I0(n2129), .I1(n47051), .I2(n34735), .I3(n2130), 
            .O(n47053));
    defparam i1_4_lut_adj_1807.LUT_INIT = 16'heccc;
    SB_LUT4 i1_4_lut_adj_1808 (.I0(n2118), .I1(n2119), .I2(n47053), .I3(n2120), 
            .O(n47059));
    defparam i1_4_lut_adj_1808.LUT_INIT = 16'hfffe;
    SB_LUT4 i36126_4_lut (.I0(n2116), .I1(n2115), .I2(n2117), .I3(n47059), 
            .O(n2148));
    defparam i36126_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1306_3_lut (.I0(n1919), .I1(n1986), 
            .I2(n1950), .I3(GND_net), .O(n2018));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1306_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1305_3_lut (.I0(n1918), .I1(n1985), 
            .I2(n1950), .I3(GND_net), .O(n2017));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1305_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1308_3_lut (.I0(n1921), .I1(n1988), 
            .I2(n1950), .I3(GND_net), .O(n2020));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1308_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 LessThan_699_i8_3_lut_3_lut (.I0(pwm_setpoint[4]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[8]), .I3(GND_net), .O(n8_adj_4965));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 encoder0_position_31__I_0_i1307_3_lut (.I0(n1920), .I1(n1987), 
            .I2(n1950), .I3(GND_net), .O(n2019));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1307_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1311_3_lut (.I0(n1924), .I1(n1991), 
            .I2(n1950), .I3(GND_net), .O(n2023));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1311_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1310_3_lut (.I0(n1923), .I1(n1990), 
            .I2(n1950), .I3(GND_net), .O(n2022));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1310_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1309_3_lut (.I0(n1922), .I1(n1989), 
            .I2(n1950), .I3(GND_net), .O(n2021));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1309_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1315_3_lut (.I0(n1928), .I1(n1995), 
            .I2(n1950), .I3(GND_net), .O(n2027));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1315_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35258_3_lut (.I0(n1927), .I1(n1994), .I2(n1950), .I3(GND_net), 
            .O(n2026));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i35258_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1319_3_lut (.I0(n1932), .I1(n1999), 
            .I2(n1950), .I3(GND_net), .O(n2031));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1319_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1318_3_lut (.I0(n1931), .I1(n1998), 
            .I2(n1950), .I3(GND_net), .O(n2030));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1318_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1317_3_lut (.I0(n1930), .I1(n1997), 
            .I2(n1950), .I3(GND_net), .O(n2029));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1317_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1313_rep_41_3_lut (.I0(n1926), .I1(n1993), 
            .I2(n1950), .I3(GND_net), .O(n2025));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1313_rep_41_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35255_3_lut (.I0(n1826), .I1(n1893), .I2(n1851), .I3(GND_net), 
            .O(n1925));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i35255_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35256_3_lut (.I0(n1925), .I1(n1992), .I2(n1950), .I3(GND_net), 
            .O(n2024));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i35256_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1316_rep_42_3_lut (.I0(n1929), .I1(n1996), 
            .I2(n1950), .I3(GND_net), .O(n2028));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1316_rep_42_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1321_3_lut (.I0(n944), .I1(n2001), 
            .I2(n1950), .I3(GND_net), .O(n2033));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1321_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1320_3_lut (.I0(n1933), .I1(n2000), 
            .I2(n1950), .I3(GND_net), .O(n2032));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1320_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i14_3_lut (.I0(encoder0_position[13]), 
            .I1(n20_adj_4922), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n945));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21570_3_lut (.I0(n945), .I1(n2032), .I2(n2033), .I3(GND_net), 
            .O(n34637));
    defparam i21570_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_2_lut_adj_1809 (.I0(n2026), .I1(n2027), .I2(GND_net), .I3(GND_net), 
            .O(n47317));
    defparam i1_2_lut_adj_1809.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1810 (.I0(n2028), .I1(n47317), .I2(n2024), .I3(n2025), 
            .O(n47321));
    defparam i1_4_lut_adj_1810.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1811 (.I0(n2029), .I1(n34637), .I2(n2030), .I3(n2031), 
            .O(n45109));
    defparam i1_4_lut_adj_1811.LUT_INIT = 16'ha080;
    SB_LUT4 i35072_2_lut_4_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(pwm_counter[4]), .I3(pwm_setpoint[4]), .O(n50024));
    defparam i35072_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i1_4_lut_adj_1812 (.I0(n2021), .I1(n2022), .I2(n2023), .I3(n47321), 
            .O(n47327));
    defparam i1_4_lut_adj_1812.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1813 (.I0(n2019), .I1(n2020), .I2(n47327), .I3(n45109), 
            .O(n47333));
    defparam i1_4_lut_adj_1813.LUT_INIT = 16'hfffe;
    SB_LUT4 i36096_4_lut (.I0(n2017), .I1(n2016), .I2(n2018), .I3(n47333), 
            .O(n2049));
    defparam i36096_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_83_i11_4_lut (.I0(encoder1_position_scaled[10]), .I1(displacement[10]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[10]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i11_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_31__I_0_i1239_3_lut (.I0(n1820), .I1(n1887), 
            .I2(n1851), .I3(GND_net), .O(n1919));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1239_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1238_3_lut (.I0(n1819), .I1(n1886), 
            .I2(n1851), .I3(GND_net), .O(n1918));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1244_3_lut (.I0(n1825), .I1(n1892), 
            .I2(n1851), .I3(GND_net), .O(n1924));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1244_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1241_3_lut (.I0(n1822), .I1(n1889), 
            .I2(n1851), .I3(GND_net), .O(n1921));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1241_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1240_3_lut (.I0(n1821), .I1(n1888), 
            .I2(n1851), .I3(GND_net), .O(n1920));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1246_3_lut (.I0(n1827), .I1(n1894), 
            .I2(n1851), .I3(GND_net), .O(n1926));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1246_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1243_3_lut (.I0(n1824), .I1(n1891), 
            .I2(n1851), .I3(GND_net), .O(n1923));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1243_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1242_3_lut (.I0(n1823), .I1(n1890), 
            .I2(n1851), .I3(GND_net), .O(n1922));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1242_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1814 (.I0(n1926), .I1(n1928), .I2(GND_net), .I3(GND_net), 
            .O(n46929));
    defparam i1_2_lut_adj_1814.LUT_INIT = 16'heeee;
    SB_LUT4 i1_3_lut_adj_1815 (.I0(n1925), .I1(n1924), .I2(n1927), .I3(GND_net), 
            .O(n46931));
    defparam i1_3_lut_adj_1815.LUT_INIT = 16'hfefe;
    SB_LUT4 i21574_3_lut (.I0(n944), .I1(n1932), .I2(n1933), .I3(GND_net), 
            .O(n34641));
    defparam i21574_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i1_4_lut_adj_1816 (.I0(n1922), .I1(n1923), .I2(n46931), .I3(n46929), 
            .O(n46937));
    defparam i1_4_lut_adj_1816.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1817 (.I0(n1929), .I1(n34641), .I2(n1930), .I3(n1931), 
            .O(n45073));
    defparam i1_4_lut_adj_1817.LUT_INIT = 16'ha080;
    SB_LUT4 i1_4_lut_adj_1818 (.I0(n1920), .I1(n45073), .I2(n1921), .I3(n46937), 
            .O(n46943));
    defparam i1_4_lut_adj_1818.LUT_INIT = 16'hfffe;
    SB_LUT4 i36071_4_lut (.I0(n1918), .I1(n1917), .I2(n1919), .I3(n46943), 
            .O(n1950));
    defparam i36071_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i1108_3_lut (.I0(n1625), .I1(n1692), 
            .I2(n1653), .I3(GND_net), .O(n1724));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1108_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15238_3_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(timer[15]), 
            .I2(n43085), .I3(GND_net), .O(n28301));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15238_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1107_3_lut (.I0(n1624), .I1(n1691), 
            .I2(n1653), .I3(GND_net), .O(n1723));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1107_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1037_3_lut (.I0(n1522), .I1(n1589), 
            .I2(n1554), .I3(GND_net), .O(n1621));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1037_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15239_3_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(timer[14]), 
            .I2(n43085), .I3(GND_net), .O(n28302));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15239_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1038_3_lut (.I0(n1523), .I1(n1590), 
            .I2(n1554), .I3(GND_net), .O(n1622));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1038_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1252_3_lut (.I0(n1833), .I1(n1900), 
            .I2(n1851), .I3(GND_net), .O(n1932));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1252_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_adj_1819 (.I0(delay_counter[12]), .I1(delay_counter[11]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_4985));
    defparam i1_2_lut_adj_1819.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_1820 (.I0(delay_counter[9]), .I1(n4_adj_4985), 
            .I2(delay_counter[10]), .I3(n26508), .O(n46246));
    defparam i2_4_lut_adj_1820.LUT_INIT = 16'hfcec;
    SB_LUT4 i2_4_lut_adj_1821 (.I0(n46246), .I1(n26502), .I2(delay_counter[13]), 
            .I3(delay_counter[14]), .O(n45439));
    defparam i2_4_lut_adj_1821.LUT_INIT = 16'hffec;
    SB_LUT4 i3_3_lut (.I0(delay_counter[20]), .I1(delay_counter[21]), .I2(delay_counter[23]), 
            .I3(GND_net), .O(n8_adj_5023));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i2_4_lut_adj_1822 (.I0(delay_counter[22]), .I1(n45439), .I2(delay_counter[19]), 
            .I3(delay_counter[18]), .O(n7_adj_5024));
    defparam i2_4_lut_adj_1822.LUT_INIT = 16'ha8a0;
    SB_LUT4 i20809_4_lut (.I0(n7_adj_5024), .I1(delay_counter[31]), .I2(n26505), 
            .I3(n8_adj_5023), .O(n777));   // verilog/TinyFPGA_B.v(280[14:38])
    defparam i20809_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i35864_1_lut (.I0(n1257), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50817));
    defparam i35864_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_4_lut (.I0(delay_counter[27]), .I1(delay_counter[29]), .I2(delay_counter[24]), 
            .I3(delay_counter[26]), .O(n12_adj_4888));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35830_1_lut (.I0(n1059), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n50783));
    defparam i35830_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i6_4_lut (.I0(delay_counter[28]), .I1(n12_adj_4888), .I2(delay_counter[25]), 
            .I3(delay_counter[30]), .O(n26505));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_3_lut_adj_1823 (.I0(delay_counter[3]), .I1(delay_counter[5]), 
            .I2(delay_counter[4]), .I3(GND_net), .O(n14_adj_4946));
    defparam i5_3_lut_adj_1823.LUT_INIT = 16'hfefe;
    SB_LUT4 i6_4_lut_adj_1824 (.I0(delay_counter[8]), .I1(delay_counter[7]), 
            .I2(delay_counter[1]), .I3(delay_counter[0]), .O(n15_adj_4945));
    defparam i6_4_lut_adj_1824.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n15_adj_4945), .I1(delay_counter[2]), .I2(n14_adj_4946), 
            .I3(delay_counter[6]), .O(n26508));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i2_3_lut_adj_1825 (.I0(delay_counter[17]), .I1(delay_counter[16]), 
            .I2(delay_counter[15]), .I3(GND_net), .O(n26502));
    defparam i2_3_lut_adj_1825.LUT_INIT = 16'hfefe;
    SB_LUT4 i3760_4_lut (.I0(n26508), .I1(delay_counter[11]), .I2(delay_counter[10]), 
            .I3(delay_counter[9]), .O(n24_adj_4960));
    defparam i3760_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i2_4_lut_adj_1826 (.I0(n24_adj_4960), .I1(delay_counter[14]), 
            .I2(delay_counter[12]), .I3(delay_counter[13]), .O(n45377));
    defparam i2_4_lut_adj_1826.LUT_INIT = 16'hc800;
    SB_LUT4 i2_3_lut_adj_1827 (.I0(n45377), .I1(delay_counter[18]), .I2(n26502), 
            .I3(GND_net), .O(n45435));
    defparam i2_3_lut_adj_1827.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_4_lut_adj_1828 (.I0(enable_slow_N_4090), .I1(data_ready), 
            .I2(state_adj_5100[1]), .I3(state_adj_5100[0]), .O(n43797));   // verilog/eeprom.v(26[8] 58[4])
    defparam i1_4_lut_adj_1828.LUT_INIT = 16'hccd0;
    SB_LUT4 i15154_4_lut (.I0(rw), .I1(state_adj_5100[0]), .I2(state_adj_5100[1]), 
            .I3(n4227), .O(n28217));   // verilog/eeprom.v(26[8] 58[4])
    defparam i15154_4_lut.LUT_INIT = 16'hacaa;
    SB_LUT4 i2_4_lut_adj_1829 (.I0(delay_counter[23]), .I1(n45435), .I2(delay_counter[20]), 
            .I3(delay_counter[19]), .O(n7));
    defparam i2_4_lut_adj_1829.LUT_INIT = 16'heaaa;
    SB_LUT4 i4_4_lut_adj_1830 (.I0(n7), .I1(delay_counter[21]), .I2(delay_counter[22]), 
            .I3(n26505), .O(n62));
    defparam i4_4_lut_adj_1830.LUT_INIT = 16'hfffe;
    SB_LUT4 i20808_2_lut (.I0(n62), .I1(delay_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(read_N_321));   // verilog/TinyFPGA_B.v(265[12:35])
    defparam i20808_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_2_lut_adj_1831 (.I0(ID[2]), .I1(ID[4]), .I2(GND_net), .I3(GND_net), 
            .O(n10_adj_4987));   // verilog/TinyFPGA_B.v(278[12:17])
    defparam i2_2_lut_adj_1831.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1832 (.I0(ID[7]), .I1(ID[5]), .I2(ID[1]), .I3(ID[0]), 
            .O(n14_adj_4986));   // verilog/TinyFPGA_B.v(278[12:17])
    defparam i6_4_lut_adj_1832.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(ID[3]), .I1(n14_adj_4986), .I2(n10_adj_4987), 
            .I3(ID[6]), .O(n26483));   // verilog/TinyFPGA_B.v(278[12:17])
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 \ID_READOUT_FSM.state_2__I_0_i5_2_lut  (.I0(\ID_READOUT_FSM.state [0]), 
            .I1(\ID_READOUT_FSM.state [1]), .I2(GND_net), .I3(GND_net), 
            .O(n5_adj_4947));   // verilog/TinyFPGA_B.v(277[7:11])
    defparam \ID_READOUT_FSM.state_2__I_0_i5_2_lut .LUT_INIT = 16'hbbbb;
    SB_LUT4 i15155_4_lut (.I0(r_Rx_Data), .I1(rx_data[3]), .I2(n4_adj_4916), 
            .I3(n26624), .O(n28218));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15155_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i15156_4_lut (.I0(r_Rx_Data), .I1(rx_data[4]), .I2(n4_adj_4942), 
            .I3(n26629), .O(n28219));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15156_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i14981_4_lut (.I0(n5722), .I1(n777), .I2(n49714), .I3(n26484), 
            .O(n28044));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i14981_4_lut.LUT_INIT = 16'ha088;
    SB_LUT4 i15240_3_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(timer[13]), 
            .I2(n43085), .I3(GND_net), .O(n28303));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15240_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15241_3_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(timer[12]), 
            .I2(n43085), .I3(GND_net), .O(n28304));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15241_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_83_i12_4_lut (.I0(encoder1_position_scaled[11]), .I1(displacement[11]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[11]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i12_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1399_4_lut_4_lut (.I0(\ID_READOUT_FSM.state [0]), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(n777), .I3(n26483), .O(n5855));   // verilog/TinyFPGA_B.v(262[5] 286[12])
    defparam i1399_4_lut_4_lut.LUT_INIT = 16'hcc8c;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i13_1_lut (.I0(encoder1_position_scaled[12]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n13_adj_4899));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15242_3_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(timer[11]), 
            .I2(n43085), .I3(GND_net), .O(n28305));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15242_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1251_3_lut (.I0(n1832), .I1(n1899), 
            .I2(n1851), .I3(GND_net), .O(n1931));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1251_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_4_lut (.I0(data_ready), .I1(n62), .I2(delay_counter[31]), 
            .I3(\ID_READOUT_FSM.state [0]), .O(n6_adj_5041));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h080c;
    SB_LUT4 mux_83_i13_4_lut (.I0(encoder1_position_scaled[12]), .I1(displacement[12]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[12]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i13_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15243_3_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(timer[10]), 
            .I2(n43085), .I3(GND_net), .O(n28306));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15243_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1106_3_lut (.I0(n1623), .I1(n1690), 
            .I2(n1653), .I3(GND_net), .O(n1722));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1106_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15244_3_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(timer[9]), 
            .I2(n43085), .I3(GND_net), .O(n28307));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15244_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i15158_4_lut (.I0(r_Rx_Data), .I1(rx_data[5]), .I2(n4_adj_4942), 
            .I3(n26624), .O(n28221));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15158_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 encoder0_position_31__I_0_i706_3_lut (.I0(n1031), .I1(n1098), 
            .I2(n1059), .I3(GND_net), .O(n1130));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i706_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i705_3_lut (.I0(n1030), .I1(n1097), 
            .I2(n1059), .I3(GND_net), .O(n1129));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i705_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i701_3_lut (.I0(n1026), .I1(n1093), 
            .I2(n1059), .I3(GND_net), .O(n1125));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i701_3_lut.LUT_INIT = 16'hacac;
    \quadrature_decoder(1,500000)  quad_counter1 (.b_prev(b_prev_adj_4940), 
            .GND_net(GND_net), .a_new({a_new_adj_5076[1], Open_1}), .direction_N_3807(direction_N_3807_adj_4941), 
            .ENCODER1_B_N_keep(ENCODER1_B_N), .n1188(CLK_c), .ENCODER1_A_N_keep(ENCODER1_A_N), 
            .encoder1_position({encoder1_position}), .VCC_net(VCC_net), 
            .n28234(n28234), .n1193(n1193)) /* synthesis lattice_noprune=1 */ ;   // verilog/TinyFPGA_B.v(196[57] 203[6])
    SB_LUT4 encoder0_position_31__I_0_i1250_3_lut (.I0(n1831), .I1(n1898), 
            .I2(n1851), .I3(GND_net), .O(n1930));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1250_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i1105_3_lut (.I0(n1622), .I1(n1689), 
            .I2(n1653), .I3(GND_net), .O(n1721));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1105_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_2_lut_3_lut_adj_1833 (.I0(n5728), .I1(n33308), .I2(n61), 
            .I3(GND_net), .O(n44058));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1833.LUT_INIT = 16'h0e0e;
    SB_LUT4 i21610_4_lut (.I0(n834), .I1(n831), .I2(n832), .I3(n833), 
            .O(n34677));
    defparam i21610_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_4_lut (.I0(n44035), .I1(n33308), .I2(tx_transmit_N_3413), 
            .I3(n40), .O(n8_adj_5037));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h2220;
    SB_LUT4 i15178_3_lut_4_lut (.I0(n1152), .I1(b_prev), .I2(a_new[1]), 
            .I3(direction_N_3807), .O(n28241));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i15178_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 i12_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n27803), 
            .I3(rx_data_ready), .O(n43659));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i12_3_lut_4_lut.LUT_INIT = 16'h4f40;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main_2__N_3442[2]), .O(n44048));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h4000;
    SB_LUT4 i21751_4_lut (.I0(n829), .I1(n828), .I2(n34677), .I3(n830), 
            .O(n861));
    defparam i21751_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 mux_83_i14_4_lut (.I0(encoder1_position_scaled[13]), .I1(displacement[13]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[13]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i14_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i13_3_lut_4_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), 
            .I2(r_SM_Main[0]), .I3(r_SM_Main_2__N_3442[2]), .O(n27803));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i13_3_lut_4_lut_4_lut.LUT_INIT = 16'h4303;
    SB_LUT4 i29924_3_lut (.I0(n4_adj_4951), .I1(n6536), .I2(n44804), .I3(GND_net), 
            .O(n44807));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i29924_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i29925_3_lut (.I0(encoder0_position[29]), .I1(n44807), .I2(encoder0_position[31]), 
            .I3(GND_net), .O(n830));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam i29925_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i21608_4_lut (.I0(n934), .I1(n931), .I2(n932), .I3(n933), 
            .O(n34675));
    defparam i21608_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_2_lut_adj_1834 (.I0(n929), .I1(n930), .I2(GND_net), .I3(GND_net), 
            .O(n47213));
    defparam i1_2_lut_adj_1834.LUT_INIT = 16'h8888;
    pll32MHz pll32MHz_inst (.GND_net(GND_net), .CLK_c(CLK_c), .VCC_net(VCC_net), 
            .clk32MHz(clk32MHz)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    SB_LUT4 i1_4_lut_adj_1835 (.I0(n927), .I1(n47213), .I2(n928), .I3(n34675), 
            .O(n960));
    defparam i1_4_lut_adj_1835.LUT_INIT = 16'hfefa;
    SB_LUT4 encoder0_position_31__I_0_i569_3_lut (.I0(n830), .I1(n897), 
            .I2(n861), .I3(GND_net), .O(n929));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i569_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1115_3_lut (.I0(n1632), .I1(n1699), 
            .I2(n1653), .I3(GND_net), .O(n1731));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1115_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21477_3_lut (.I0(n935), .I1(n1032), .I2(n1033), .I3(GND_net), 
            .O(n34541));
    defparam i21477_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i14_1_lut (.I0(encoder1_position_scaled[13]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n12_adj_4898));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i15_1_lut (.I0(encoder1_position_scaled[14]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n11_adj_4897));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_83_i15_4_lut (.I0(encoder1_position_scaled[14]), .I1(displacement[14]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[14]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i15_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i1_2_lut_4_lut_adj_1836 (.I0(control_mode[0]), .I1(control_mode[6]), 
            .I2(n10_adj_5040), .I3(control_mode[2]), .O(n26480));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam i1_2_lut_4_lut_adj_1836.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i16_1_lut (.I0(encoder1_position_scaled[15]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n10_adj_4896));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i1_4_lut_adj_1837 (.I0(n1029), .I1(n34541), .I2(n1030), .I3(n1031), 
            .O(n45031));
    defparam i1_4_lut_adj_1837.LUT_INIT = 16'ha080;
    SB_LUT4 mux_83_i16_4_lut (.I0(encoder1_position_scaled[15]), .I1(displacement[15]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[15]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i16_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i35833_4_lut (.I0(n1026), .I1(n45031), .I2(n1027), .I3(n1028), 
            .O(n1059));
    defparam i35833_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 encoder0_position_31__I_0_i636_3_lut (.I0(n929), .I1(n996), 
            .I2(n960), .I3(GND_net), .O(n1028));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i636_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i704_3_lut (.I0(n1029), .I1(n1096), 
            .I2(n1059), .I3(GND_net), .O(n1128));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i704_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i703_3_lut (.I0(n1028), .I1(n1095), 
            .I2(n1059), .I3(GND_net), .O(n1127));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i703_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i709_3_lut (.I0(n935), .I1(n1101), 
            .I2(n1059), .I3(GND_net), .O(n1133));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i709_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i16_4_lut_4_lut (.I0(state_adj_5116[0]), .I1(n49785), .I2(n5538), 
            .I3(n10_adj_4935), .O(n8_adj_4958));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i16_4_lut_4_lut.LUT_INIT = 16'h3a7a;
    SB_LUT4 encoder0_position_31__I_0_i708_3_lut (.I0(n1033), .I1(n1100), 
            .I2(n1059), .I3(GND_net), .O(n1132));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i708_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i17_1_lut (.I0(encoder1_position_scaled[16]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n9_adj_4895));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i15171_3_lut_4_lut (.I0(n1193), .I1(b_prev_adj_4940), .I2(a_new_adj_5076[1]), 
            .I3(direction_N_3807_adj_4941), .O(n28234));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i15171_3_lut_4_lut.LUT_INIT = 16'h3caa;
    SB_LUT4 mux_83_i17_4_lut (.I0(encoder1_position_scaled[16]), .I1(displacement[16]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[16]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i17_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i18_1_lut (.I0(encoder1_position_scaled[17]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n8_adj_4894));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 encoder0_position_31__I_0_i707_3_lut (.I0(n1032), .I1(n1099), 
            .I2(n1059), .I3(GND_net), .O(n1131));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i707_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_83_i18_4_lut (.I0(encoder1_position_scaled[17]), .I1(displacement[17]), 
            .I2(n15), .I3(n15_adj_4885), .O(motor_state_23__N_106[17]));   // verilog/TinyFPGA_B.v(169[5] 171[10])
    defparam mux_83_i18_4_lut.LUT_INIT = 16'h0aca;
    SB_LUT4 i15159_4_lut (.I0(r_Rx_Data), .I1(rx_data[6]), .I2(n33765), 
            .I3(n26629), .O(n28222));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15159_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 encoder0_position_31__I_0_i1045_3_lut (.I0(n1530), .I1(n1597), 
            .I2(n1554), .I3(GND_net), .O(n1629));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1045_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_mux_3_i23_3_lut (.I0(encoder0_position[22]), 
            .I1(n11_adj_4931), .I2(encoder0_position[31]), .I3(GND_net), 
            .O(n936));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_mux_3_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 encoder0_position_31__I_0_i1114_3_lut (.I0(n1631), .I1(n1698), 
            .I2(n1653), .I3(GND_net), .O(n1730));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1114_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i21604_4_lut (.I0(n936), .I1(n1131), .I2(n1132), .I3(n1133), 
            .O(n34671));
    defparam i21604_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 i1_3_lut_adj_1838 (.I0(n1126), .I1(n1127), .I2(n1128), .I3(GND_net), 
            .O(n47167));
    defparam i1_3_lut_adj_1838.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1839 (.I0(n1129), .I1(n1130), .I2(GND_net), .I3(GND_net), 
            .O(n47219));
    defparam i1_2_lut_adj_1839.LUT_INIT = 16'h8888;
    SB_LUT4 encoder0_position_31__I_0_i1113_3_lut (.I0(n1630), .I1(n1697), 
            .I2(n1653), .I3(GND_net), .O(n1729));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1113_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i35849_4_lut (.I0(n47219), .I1(n1125), .I2(n47167), .I3(n34671), 
            .O(n1158));
    defparam i35849_4_lut.LUT_INIT = 16'h0103;
    SB_LUT4 encoder0_position_31__I_0_i702_3_lut (.I0(n1027), .I1(n1094), 
            .I2(n1059), .I3(GND_net), .O(n1126));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i702_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 encoder0_position_31__I_0_i769_3_lut (.I0(n1126), .I1(n1193_adj_4956), 
            .I2(n1158), .I3(GND_net), .O(n1225));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i769_3_lut.LUT_INIT = 16'hacac;
    motorControl control (.\Kp[3] (Kp[3]), .GND_net(GND_net), .\Ki[8] (Ki[8]), 
            .\Kp[13] (Kp[13]), .\Kp[4] (Kp[4]), .\Kp[14] (Kp[14]), .\Ki[9] (Ki[9]), 
            .\Kp[5] (Kp[5]), .PWMLimit({PWMLimit}), .\Ki[3] (Ki[3]), .\Kp[15] (Kp[15]), 
            .\Ki[10] (Ki[10]), .\Kp[6] (Kp[6]), .\Kp[7] (Kp[7]), .\Kp[8] (Kp[8]), 
            .\Kp[9] (Kp[9]), .\Ki[11] (Ki[11]), .\Kp[10] (Kp[10]), .\Ki[4] (Ki[4]), 
            .\Ki[5] (Ki[5]), .\Ki[0] (Ki[0]), .\Kp[0] (Kp[0]), .\Kp[11] (Kp[11]), 
            .\Ki[6] (Ki[6]), .\Ki[12] (Ki[12]), .\Kp[12] (Kp[12]), .\Ki[7] (Ki[7]), 
            .\Ki[13] (Ki[13]), .\Ki[14] (Ki[14]), .\Ki[15] (Ki[15]), .\Ki[1] (Ki[1]), 
            .\Ki[2] (Ki[2]), .\Kp[1] (Kp[1]), .\Kp[2] (Kp[2]), .IntegralLimit({IntegralLimit}), 
            .duty({duty}), .clk32MHz(clk32MHz), .VCC_net(VCC_net), .setpoint({setpoint}), 
            .motor_state({motor_state}), .n51409(n51409)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(173[16] 185[4])
    SB_LUT4 i15160_4_lut (.I0(r_Rx_Data), .I1(rx_data[7]), .I2(n33765), 
            .I3(n26624), .O(n28223));   // verilog/uart_rx.v(49[10] 144[8])
    defparam i15160_4_lut.LUT_INIT = 16'hccac;
    SB_LUT4 i15161_4_lut (.I0(saved_addr[0]), .I1(rw), .I2(state_7__N_3987[0]), 
            .I3(enable_slow_N_4090), .O(n28224));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i15161_4_lut.LUT_INIT = 16'haaca;
    SB_LUT4 encoder0_position_scaled_23__I_0_inv_0_i19_1_lut (.I0(encoder1_position_scaled[18]), 
            .I1(GND_net), .I2(GND_net), .I3(GND_net), .O(n7_adj_4893));   // verilog/TinyFPGA_B.v(224[21:72])
    defparam encoder0_position_scaled_23__I_0_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i2_2_lut_adj_1840 (.I0(pwm_counter[28]), .I1(pwm_counter[29]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_5044));
    defparam i2_2_lut_adj_1840.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1841 (.I0(pwm_counter[26]), .I1(pwm_counter[23]), 
            .I2(pwm_counter[27]), .I3(pwm_counter[25]), .O(n14_adj_5043));
    defparam i6_4_lut_adj_1841.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1842 (.I0(pwm_counter[30]), .I1(n14_adj_5043), 
            .I2(n10_adj_5044), .I3(pwm_counter[24]), .O(n26490));
    defparam i7_4_lut_adj_1842.LUT_INIT = 16'hfffe;
    SB_LUT4 encoder0_position_31__I_0_i1044_3_lut (.I0(n1529), .I1(n1596), 
            .I2(n1554), .I3(GND_net), .O(n1628));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1044_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_3_lut_adj_1843 (.I0(data_ready), .I1(\ID_READOUT_FSM.state [1]), 
            .I2(\ID_READOUT_FSM.state [0]), .I3(GND_net), .O(n46808));
    defparam i2_3_lut_adj_1843.LUT_INIT = 16'hdfdf;
    SB_LUT4 i15162_3_lut (.I0(ID[0]), .I1(data[0]), .I2(n46808), .I3(GND_net), 
            .O(n28225));   // verilog/TinyFPGA_B.v(259[10] 287[6])
    defparam i15162_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i1_4_lut_adj_1844 (.I0(n26881), .I1(n27546), .I2(\data_out_frame[20] [0]), 
            .I3(n44240), .O(n44436));
    defparam i1_4_lut_adj_1844.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1845 (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[20] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n44685));
    defparam i1_2_lut_adj_1845.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_699_i9_2_lut (.I0(pwm_counter[4]), .I1(pwm_setpoint[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4966));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_81_i1_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[0]), 
            .I3(encoder0_position_scaled[0]), .O(motor_state[0]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i1_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 LessThan_699_i11_2_lut (.I0(pwm_counter[5]), .I1(pwm_setpoint[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4968));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_699_i17_2_lut (.I0(pwm_counter[8]), .I1(pwm_setpoint[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4972));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_699_i27_2_lut (.I0(pwm_counter[13]), .I1(pwm_setpoint[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4977));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_699_i15_2_lut (.I0(pwm_counter[7]), .I1(pwm_setpoint[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4971));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_81_i2_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[1]), 
            .I3(encoder0_position_scaled[1]), .O(motor_state[1]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i2_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 LessThan_699_i13_2_lut (.I0(pwm_counter[6]), .I1(pwm_setpoint[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4970));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_699_i7_2_lut (.I0(pwm_counter[3]), .I1(pwm_setpoint[3]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4964));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i7_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_699_i21_2_lut (.I0(pwm_counter[10]), .I1(pwm_setpoint[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4974));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_699_i23_2_lut (.I0(pwm_counter[11]), .I1(pwm_setpoint[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4975));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_81_i3_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[2]), 
            .I3(encoder0_position_scaled[2]), .O(motor_state[2]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i3_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_81_i4_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[3]), 
            .I3(encoder0_position_scaled[3]), .O(motor_state[3]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i4_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_81_i5_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[4]), 
            .I3(encoder0_position_scaled[4]), .O(motor_state[4]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i5_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_81_i6_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[5]), 
            .I3(encoder0_position_scaled[5]), .O(motor_state[5]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i6_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_81_i7_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[6]), 
            .I3(encoder0_position_scaled[6]), .O(motor_state[6]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i7_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_81_i8_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[7]), 
            .I3(encoder0_position_scaled[7]), .O(motor_state[7]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i8_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 LessThan_699_i19_2_lut (.I0(pwm_counter[9]), .I1(pwm_setpoint[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4973));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_699_i29_2_lut (.I0(pwm_counter[14]), .I1(pwm_setpoint[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4978));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mux_81_i9_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[8]), 
            .I3(encoder0_position_scaled[8]), .O(motor_state[8]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i9_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_81_i10_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[9]), 
            .I3(encoder0_position_scaled[9]), .O(motor_state[9]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i10_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_81_i11_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[10]), 
            .I3(encoder0_position_scaled[10]), .O(motor_state[10]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i11_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_81_i12_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[11]), 
            .I3(encoder0_position_scaled[11]), .O(motor_state[11]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i12_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 LessThan_699_i31_2_lut (.I0(pwm_counter[15]), .I1(pwm_setpoint[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4980));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_699_i33_2_lut (.I0(pwm_counter[16]), .I1(pwm_setpoint[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4981));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_699_i35_2_lut (.I0(pwm_counter[17]), .I1(pwm_setpoint[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_699_i25_2_lut (.I0(pwm_counter[12]), .I1(pwm_setpoint[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4976));   // verilog/pwm.v(21[8:24])
    defparam LessThan_699_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1846 (.I0(n26490), .I1(pwm_counter[31]), .I2(GND_net), 
            .I3(GND_net), .O(n26492));
    defparam i1_2_lut_adj_1846.LUT_INIT = 16'heeee;
    SB_LUT4 mux_81_i13_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[12]), 
            .I3(encoder0_position_scaled[12]), .O(motor_state[12]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i13_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i19_3_lut (.I0(\data_out_frame[16] [6]), .I1(\data_out_frame[17] [6]), 
            .I2(byte_transmit_counter[0]), .I3(GND_net), .O(n15_adj_4913));   // verilog/coms.v(102[12:33])
    defparam i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35050_2_lut (.I0(\data_out_frame[23] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49819));
    defparam i35050_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35052_2_lut (.I0(\data_out_frame[20] [6]), .I1(byte_transmit_counter[0]), 
            .I2(GND_net), .I3(GND_net), .O(n49818));
    defparam i35052_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mux_81_i14_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[13]), 
            .I3(encoder0_position_scaled[13]), .O(motor_state[13]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i14_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_81_i15_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[14]), 
            .I3(encoder0_position_scaled[14]), .O(motor_state[14]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i15_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_81_i16_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[15]), 
            .I3(encoder0_position_scaled[15]), .O(motor_state[15]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i16_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_81_i17_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[16]), 
            .I3(encoder0_position_scaled[16]), .O(motor_state[16]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i17_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_81_i18_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[17]), 
            .I3(encoder0_position_scaled[17]), .O(motor_state[17]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i18_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    coms neopxl_color_23__I_0 (.rx_data({rx_data}), .CLK_c(CLK_c), .\data_out_frame[9] ({\data_out_frame[9] }), 
         .\data_out_frame[4] ({\data_out_frame[4] }), .GND_net(GND_net), 
         .\data_out_frame[8] ({\data_out_frame[8] }), .\data_out_frame[13] ({\data_out_frame[13] }), 
         .\data_out_frame[18] ({\data_out_frame[18] [7:3], Open_2, Open_3, 
         Open_4}), .\data_out_frame[16] ({\data_out_frame[16] }), .\data_out_frame[20] ({\data_out_frame[20] }), 
         .\data_out_frame[25] ({\data_out_frame[25] }), .\data_out_frame[11] ({\data_out_frame[11] }), 
         .\data_out_frame[15] ({\data_out_frame[15] }), .\data_out_frame[23] ({\data_out_frame[23] }), 
         .\data_out_frame[14] ({\data_out_frame[14] }), .\data_out_frame[7] ({\data_out_frame[7] }), 
         .\data_out_frame[12] ({\data_out_frame[12] }), .\data_out_frame[5] ({\data_out_frame[5] }), 
         .\data_out_frame[10] ({\data_out_frame[10] }), .\data_out_frame[17] ({\data_out_frame[17] }), 
         .\data_out_frame[19] ({\data_out_frame[19] }), .\data_out_frame[6] ({\data_out_frame[6] }), 
         .\byte_transmit_counter[2] (byte_transmit_counter[2]), .\FRAME_MATCHER.state ({Open_5, 
         Open_6, Open_7, Open_8, Open_9, Open_10, Open_11, Open_12, 
         Open_13, Open_14, Open_15, Open_16, Open_17, Open_18, Open_19, 
         Open_20, Open_21, Open_22, Open_23, Open_24, Open_25, Open_26, 
         Open_27, Open_28, Open_29, Open_30, Open_31, Open_32, \FRAME_MATCHER.state [3], 
         Open_33, Open_34, Open_35}), .\data_in_frame[2] ({\data_in_frame[2] }), 
         .\data_in_frame[1] ({\data_in_frame[1] }), .\data_in_frame[8] ({\data_in_frame[8] }), 
         .n44058(n44058), .n33302(n33302), .n23831(n23831), .n46759(n46759), 
         .n40(n40), .n33308(n33308), .n5728(n5728), .n44035(n44035), 
         .n61(n61), .n76(n76), .n2482(n2482), .n29985(n29985), .n63(n63), 
         .n51904(n51904), .\FRAME_MATCHER.i_31__N_2524 (\FRAME_MATCHER.i_31__N_2524 ), 
         .n3303(n3303), .n5(n5_adj_4982), .\FRAME_MATCHER.i_31__N_2526 (\FRAME_MATCHER.i_31__N_2526 ), 
         .n4452(n4452), .n7(n7_adj_4983), .\data_in_frame[9] ({\data_in_frame[9] }), 
         .\displacement[17] (displacement[17]), .n23935(n23935), .rx_data_ready(rx_data_ready), 
         .n33298(n33298), .\FRAME_MATCHER.state[0] (\FRAME_MATCHER.state [0]), 
         .n73(n73), .setpoint({setpoint}), .\byte_transmit_counter[0] (byte_transmit_counter[0]), 
         .tx_transmit_N_3413(tx_transmit_N_3413), .\data_in_frame[10] ({\data_in_frame[10] }), 
         .\FRAME_MATCHER.i[31] (\FRAME_MATCHER.i [31]), .\data_in_frame[11] ({\data_in_frame[11] }), 
         .n28284(n28284), .control_mode({control_mode}), .n28283(n28283), 
         .n28282(n28282), .n28281(n28281), .n28280(n28280), .n28279(n28279), 
         .n771(n771), .n26687(n26687), .n1476(n1476), .n28278(n28278), 
         .n28277(n28277), .PWMLimit({PWMLimit}), .n28276(n28276), .n28275(n28275), 
         .n28274(n28274), .n28273(n28273), .n26489(n26489), .\data_in[3] ({\data_in[3] }), 
         .\data_in[1] ({\data_in[1] }), .\data_in[0] ({\data_in[0] }), .\data_in[2] ({\data_in[2] }), 
         .n28272(n28272), .n28271(n28271), .\data_in_frame[12] ({\data_in_frame[12] }), 
         .\data_in_frame[3] ({\data_in_frame[3] }), .\data_in_frame[13] ({\data_in_frame[13] }), 
         .n28270(n28270), .n28269(n28269), .n28268(n28268), .n28267(n28267), 
         .n28266(n28266), .n28265(n28265), .n28264(n28264), .n28263(n28263), 
         .n28262(n28262), .n28261(n28261), .n28260(n28260), .n28259(n28259), 
         .n28258(n28258), .n28257(n28257), .n28256(n28256), .n28255(n28255), 
         .n51636(n51636), .n51637(n51637), .\state[2] (state_adj_5116[2]), 
         .\state[3] (state_adj_5116[3]), .n10(n10_adj_4955), .n27771(n27771), 
         .n43485(n43485), .n49817(n49817), .\data_out_frame[24] ({\data_out_frame[24] }), 
         .n51546(n51546), .\data_out_frame[18][0] (\data_out_frame[18] [0]), 
         .n28214(n28214), .n27546(n27546), .DE_c(DE_c), .LED_c(LED_c), 
         .n74(n74), .n28213(n28213), .n44240(n44240), .n28211(n28211), 
         .neopxl_color({neopxl_color}), .n28210(n28210), .\Ki[0] (Ki[0]), 
         .n28209(n28209), .\Kp[0] (Kp[0]), .n28208(n28208), .n28759(n28759), 
         .IntegralLimit({IntegralLimit}), .n28758(n28758), .n28757(n28757), 
         .n28756(n28756), .n28755(n28755), .n28754(n28754), .n28753(n28753), 
         .n28752(n28752), .n28751(n28751), .n28750(n28750), .n28749(n28749), 
         .n28748(n28748), .n28747(n28747), .n28746(n28746), .n28745(n28745), 
         .n28744(n28744), .n28743(n28743), .n28742(n28742), .n28741(n28741), 
         .n28740(n28740), .n28739(n28739), .n28738(n28738), .n28737(n28737), 
         .n28736(n28736), .n28735(n28735), .n28734(n28734), .n28733(n28733), 
         .n28732(n28732), .n28731(n28731), .n28730(n28730), .n28729(n28729), 
         .n28728(n28728), .n28727(n28727), .\data_in_frame[5] ({\data_in_frame[5] }), 
         .\data_in_frame[6] ({\data_in_frame[6] }), .\data_in_frame[4] ({\data_in_frame[4] }), 
         .n28726(n28726), .n28725(n28725), .n28724(n28724), .n28723(n28723), 
         .n28722(n28722), .n28721(n28721), .n28720(n28720), .n28719(n28719), 
         .n28718(n28718), .n28717(n28717), .n28716(n28716), .n28715(n28715), 
         .n28714(n28714), .n28713(n28713), .n28712(n28712), .n28711(n28711), 
         .n28710(n28710), .n28709(n28709), .n28708(n28708), .n28707(n28707), 
         .n28706(n28706), .n28705(n28705), .\Kp[1] (Kp[1]), .n28704(n28704), 
         .\Kp[2] (Kp[2]), .n28703(n28703), .\Kp[3] (Kp[3]), .n28702(n28702), 
         .\Kp[4] (Kp[4]), .n28701(n28701), .\Kp[5] (Kp[5]), .n28700(n28700), 
         .\Kp[6] (Kp[6]), .n28699(n28699), .\Kp[7] (Kp[7]), .n28698(n28698), 
         .\Kp[8] (Kp[8]), .n28697(n28697), .\Kp[9] (Kp[9]), .n28696(n28696), 
         .\Kp[10] (Kp[10]), .n28695(n28695), .\Kp[11] (Kp[11]), .n28694(n28694), 
         .\Kp[12] (Kp[12]), .n28693(n28693), .\Kp[13] (Kp[13]), .n28692(n28692), 
         .\Kp[14] (Kp[14]), .n28691(n28691), .\Kp[15] (Kp[15]), .n28690(n28690), 
         .\Ki[1] (Ki[1]), .n28689(n28689), .\Ki[2] (Ki[2]), .n28688(n28688), 
         .\Ki[3] (Ki[3]), .n28687(n28687), .\Ki[4] (Ki[4]), .n28686(n28686), 
         .\Ki[5] (Ki[5]), .n28685(n28685), .\Ki[6] (Ki[6]), .n28684(n28684), 
         .\Ki[7] (Ki[7]), .n28683(n28683), .\Ki[8] (Ki[8]), .n28682(n28682), 
         .\Ki[9] (Ki[9]), .n28681(n28681), .\Ki[10] (Ki[10]), .n28680(n28680), 
         .\Ki[11] (Ki[11]), .n28679(n28679), .\Ki[12] (Ki[12]), .n28678(n28678), 
         .\Ki[13] (Ki[13]), .n28677(n28677), .\Ki[14] (Ki[14]), .n28676(n28676), 
         .\Ki[15] (Ki[15]), .n28675(n28675), .n28674(n28674), .n28673(n28673), 
         .n28672(n28672), .n28671(n28671), .n28670(n28670), .n28669(n28669), 
         .n28668(n28668), .n28667(n28667), .n28666(n28666), .n28665(n28665), 
         .n28664(n28664), .n28663(n28663), .n28662(n28662), .n28661(n28661), 
         .n28660(n28660), .n28659(n28659), .n28658(n28658), .n28657(n28657), 
         .n28656(n28656), .n28655(n28655), .n28654(n28654), .n28653(n28653), 
         .n28652(n28652), .n28651(n28651), .n28650(n28650), .n28649(n28649), 
         .n28648(n28648), .n28647(n28647), .n28646(n28646), .n28645(n28645), 
         .n28644(n28644), .n28643(n28643), .n28642(n28642), .n28641(n28641), 
         .n28640(n28640), .n28639(n28639), .n28638(n28638), .n28637(n28637), 
         .n28636(n28636), .n28635(n28635), .n28634(n28634), .n28633(n28633), 
         .n28632(n28632), .n28631(n28631), .n28630(n28630), .n28629(n28629), 
         .n28628(n28628), .n28627(n28627), .n28626(n28626), .n28625(n28625), 
         .n28624(n28624), .n28623(n28623), .n28622(n28622), .n28621(n28621), 
         .n28620(n28620), .n28619(n28619), .n28618(n28618), .n28617(n28617), 
         .n28616(n28616), .n28615(n28615), .n28614(n28614), .n28613(n28613), 
         .n28612(n28612), .n28611(n28611), .n28610(n28610), .n28609(n28609), 
         .n28608(n28608), .n28607(n28607), .n28606(n28606), .n28605(n28605), 
         .n28604(n28604), .n28603(n28603), .n28602(n28602), .n28601(n28601), 
         .n28600(n28600), .n28599(n28599), .n28598(n28598), .n28597(n28597), 
         .n28596(n28596), .n28595(n28595), .n28594(n28594), .n28593(n28593), 
         .n28592(n28592), .n28591(n28591), .n28590(n28590), .n28589(n28589), 
         .n28588(n28588), .n28587(n28587), .n28586(n28586), .n28585(n28585), 
         .n28584(n28584), .n28583(n28583), .n28582(n28582), .n28581(n28581), 
         .n28580(n28580), .n28579(n28579), .n28578(n28578), .n28577(n28577), 
         .n28576(n28576), .n28575(n28575), .n28574(n28574), .n28573(n28573), 
         .n28572(n28572), .n28571(n28571), .n28570(n28570), .n28569(n28569), 
         .n28568(n28568), .n28567(n28567), .n28566(n28566), .n28565(n28565), 
         .n28564(n28564), .n28563(n28563), .n28561(n28561), .\data_out_frame[18][2] (\data_out_frame[18] [2]), 
         .n28560(n28560), .n28559(n28559), .n28558(n28558), .n28557(n28557), 
         .n28556(n28556), .n28555(n28555), .n28554(n28554), .n28553(n28553), 
         .n28552(n28552), .n28551(n28551), .n28550(n28550), .n28549(n28549), 
         .n28548(n28548), .n28547(n28547), .n28546(n28546), .n28545(n28545), 
         .n28544(n28544), .n28543(n28543), .n28542(n28542), .n28541(n28541), 
         .n28540(n28540), .n28539(n28539), .n28538(n28538), .n28537(n28537), 
         .n28536(n28536), .n28535(n28535), .n28534(n28534), .n28533(n28533), 
         .n28532(n28532), .n28531(n28531), .n28530(n28530), .n28529(n28529), 
         .n28528(n28528), .n28527(n28527), .n28526(n28526), .n28525(n28525), 
         .n28524(n28524), .n28523(n28523), .n28522(n28522), .n28189(n28189), 
         .n28521(n28521), .n28520(n28520), .n28519(n28519), .n28518(n28518), 
         .n28517(n28517), .n28516(n28516), .n28515(n28515), .n28514(n28514), 
         .n28513(n28513), .n28512(n28512), .n28511(n28511), .n28510(n28510), 
         .n28509(n28509), .n28508(n28508), .n28507(n28507), .n28506(n28506), 
         .n28505(n28505), .n28504(n28504), .n28503(n28503), .n28502(n28502), 
         .n28501(n28501), .n28500(n28500), .n28499(n28499), .n28498(n28498), 
         .n28497(n28497), .n28496(n28496), .n28495(n28495), .n28494(n28494), 
         .n28493(n28493), .n46360(n46360), .ID({ID}), .n39(n39), .\state[0] (state_adj_5116[0]), 
         .n6014(n6014), .n44092(n44092), .n44436(n44436), .n44685(n44685), 
         .n26881(n26881), .n49818(n49818), .n49819(n49819), .n15(n15_adj_4913), 
         .tx_o(tx_o), .VCC_net(VCC_net), .tx_enable(tx_enable), .r_SM_Main({r_SM_Main}), 
         .\r_SM_Main_2__N_3442[2] (r_SM_Main_2__N_3442[2]), .\r_Bit_Index[0] (r_Bit_Index[0]), 
         .n26629(n26629), .n4(n4_adj_4938), .r_Rx_Data(r_Rx_Data), .RX_N_10(RX_N_10), 
         .n27846(n27846), .n28246(n28246), .n43659(n43659), .n28250(n28250), 
         .n28223(n28223), .n28222(n28222), .n28221(n28221), .n28219(n28219), 
         .n28218(n28218), .n43968(n43968), .n28203(n28203), .n28202(n28202), 
         .n44048(n44048), .n4_adj_10(n4_adj_4916), .n4_adj_11(n4_adj_4942), 
         .n26624(n26624), .n33765(n33765)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(140[8] 163[4])
    SB_LUT4 mux_81_i19_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[18]), 
            .I3(encoder0_position_scaled[18]), .O(motor_state[18]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i19_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_81_i20_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[19]), 
            .I3(encoder0_position_scaled[19]), .O(motor_state[19]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i20_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_81_i21_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[20]), 
            .I3(encoder0_position_scaled[20]), .O(motor_state[20]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i21_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 encoder0_position_31__I_0_i1042_3_lut (.I0(n1527), .I1(n1594), 
            .I2(n1554), .I3(GND_net), .O(n1626));   // verilog/TinyFPGA_B.v(222[33:53])
    defparam encoder0_position_31__I_0_i1042_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mux_81_i24_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[23]), 
            .I3(encoder0_position_scaled[23]), .O(motor_state[23]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i24_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 i35061_4_lut (.I0(n27_adj_4977), .I1(n15_adj_4971), .I2(n13_adj_4970), 
            .I3(n11_adj_4968), .O(n50013));
    defparam i35061_4_lut.LUT_INIT = 16'haaab;
    EEPROM eeprom (.CLK_c(CLK_c), .n4226({n4227}), .\state[1] (state_adj_5100[1]), 
           .GND_net(GND_net), .\state[0] (state_adj_5100[0]), .read(read), 
           .\state[2] (state_adj_5116[2]), .n7(n7_adj_4961), .\state[3] (state_adj_5116[3]), 
           .n6(n6_adj_4984), .n28217(n28217), .rw(rw), .n43797(n43797), 
           .data_ready(data_ready), .enable_slow_N_4090(enable_slow_N_4090), 
           .n43693(n43693), .n43685(n43685), .n44859(n44859), .n44120(n44120), 
           .n34334(n34334), .VCC_net(VCC_net), .n5538(n5538), .n33769(n33769), 
           .n4(n4_adj_4915), .scl_enable(scl_enable), .\state_7__N_4003[3] (state_7__N_4003[3]), 
           .n6014(n6014), .\state_7__N_3987[0] (state_7__N_3987[0]), .sda_enable(sda_enable), 
           .n4_adj_4(n4_adj_4914), .\saved_addr[0] (saved_addr[0]), .\state[0]_adj_5 (state_adj_5116[0]), 
           .n10(n10_adj_5039), .n10_adj_6(n10_adj_4935), .n8(n8_adj_4958), 
           .n28230(n28230), .data({data}), .n10_adj_7(n10_adj_4955), .n28224(n28224), 
           .scl(scl), .sda_out(sda_out), .n28207(n28207), .n28206(n28206), 
           .n28205(n28205), .n28204(n28204), .n28200(n28200), .n28199(n28199), 
           .n28198(n28198), .n26650(n26650), .n26645(n26645), .n49785(n49785)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(289[10] 300[6])
    SB_LUT4 mux_81_i23_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[22]), 
            .I3(encoder0_position_scaled[22]), .O(motor_state[22]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i23_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    SB_LUT4 mux_81_i22_3_lut_4_lut (.I0(n26480), .I1(control_mode[1]), .I2(motor_state_23__N_106[21]), 
            .I3(encoder0_position_scaled[21]), .O(motor_state[21]));   // verilog/TinyFPGA_B.v(168[5:22])
    defparam mux_81_i22_3_lut_4_lut.LUT_INIT = 16'h0e1f;
    pwm PWM (.n50560(n50560), .VCC_net(VCC_net), .INHA_c(INHA_c), .clk32MHz(clk32MHz), 
        .n26492(n26492), .GND_net(GND_net), .pwm_counter({pwm_counter}), 
        .n26490(n26490)) /* synthesis syn_module_defined=1 */ ;   // verilog/TinyFPGA_B.v(89[6] 94[3])
    
endmodule
//
// Verilog Description of module \neopixel(CLOCK_SPEED_HZ=16000000) 
//

module \neopixel(CLOCK_SPEED_HZ=16000000)  (n28315, \neo_pixel_transmitter.t0 , 
            CLK_c, n28314, n28313, n28312, VCC_net, GND_net, \neo_pixel_transmitter.done , 
            n28311, n28310, n28309, \state[0] , n34525, \state[1] , 
            n28308, timer, n28307, n28306, n28305, n28304, n28303, 
            n28302, n28301, n28300, n28299, n28298, n28297, n28296, 
            n28295, n28294, n28293, n28292, n28291, n28290, n28289, 
            n28288, n28287, n28286, n28285, \state_3__N_428[1] , LED_c, 
            n34629, n44839, n27916, neopxl_color, start, n43085, 
            n42985, n28194, n28188, NEOPXL_c) /* synthesis syn_module_defined=1 */ ;
    input n28315;
    output [31:0]\neo_pixel_transmitter.t0 ;
    input CLK_c;
    input n28314;
    input n28313;
    input n28312;
    input VCC_net;
    input GND_net;
    output \neo_pixel_transmitter.done ;
    input n28311;
    input n28310;
    input n28309;
    output \state[0] ;
    output n34525;
    output \state[1] ;
    input n28308;
    output [31:0]timer;
    input n28307;
    input n28306;
    input n28305;
    input n28304;
    input n28303;
    input n28302;
    input n28301;
    input n28300;
    input n28299;
    input n28298;
    input n28297;
    input n28296;
    input n28295;
    input n28294;
    input n28293;
    input n28292;
    input n28291;
    input n28290;
    input n28289;
    input n28288;
    input n28287;
    input n28286;
    input n28285;
    output \state_3__N_428[1] ;
    input LED_c;
    output n34629;
    output n44839;
    output n27916;
    input [23:0]neopxl_color;
    output start;
    output n43085;
    input n42985;
    input n28194;
    input n28188;
    output NEOPXL_c;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [31:0]n2951;
    
    wire n2887, n40584;
    wire [31:0]n1;
    
    wire \neo_pixel_transmitter.done_N_636 , n51632, n2789;
    wire [31:0]n2852;
    
    wire n2819, n2888, n40998, n44851, n50261, n49769, n26525, 
        n44943, n50262, n44987, \neo_pixel_transmitter.done_N_642 ;
    wire [31:0]bit_ctr;   // verilog/neopixel.v(18[12:19])
    
    wire n1203, n1209, n12, n1208, n1205, n1207, n1204, n13, 
        n1206, n1202, n1235, n1999;
    wire [31:0]n2060;
    
    wire n2027, n2098, n1997, n2096, n1998, n2097, n1996, n2095, 
        n2109, n2009, n2108, n2007, n2106, n2006, n2105, n2008, 
        n2107, n2003, n2102, n2001, n2100, n2002, n2101, n2000, 
        n2099, n2005, n2104, n2004, n2103, n1995, n2094, n2093, 
        n18, n24_adj_4769, n30, n28, n29, n27, n2126;
    wire [31:0]n255;
    
    wire n27743, n28088, n40585, n40583, n2889, n40582;
    wire [31:0]one_wire_N_579;
    
    wire n39183, n39049, n39050;
    wire [31:0]n1961;
    
    wire n1928, n1898, n1906, n1897, n1896, n2890, n40581, n1908, 
        n1905, n1909, n1904, n1899, n1907, n1903, n1902, n1900, 
        n1901, n20, n28_adj_4771, n26, n27_adj_4772, n1994, n25_adj_4773, 
        n1808;
    wire [31:0]n1862;
    
    wire n1829, n1809, n1807, n1801, n1799, n1800, n1798, n1797, 
        n1805, n1803, n1804, n1802, n1806, n21, n39184, n2891, 
        n40580, n25_adj_4774, n1895, n16, n24_adj_4775, n28_adj_4776, 
        n34485, n2892, n40579, n18_adj_4777, n24_adj_4778, n1796, 
        n22, n39182, n26_adj_4780, n2893, n40578, n2894, n40577, 
        n1730, n51405, n1600;
    wire [31:0]n1664;
    
    wire n1631, n1699, n1603, n1702, n1599, n1698, n1709, n1609, 
        n1708, n1602, n1701, n1606, n1705, n1605, n1704, n1607, 
        n1706, n1601, n1700, n2895, n40576, n1608, n1707, n1604, 
        n1703, n16_adj_4781, n22_adj_4782, n20_adj_4783, n24_adj_4784, 
        n1697, n2896, n40575, n2897, n40574, n2898, n40573, n2899, 
        n40572, n2900, n40571, n2901, n40570, n1509;
    wire [31:0]n1565;
    
    wire n1532, n1503, n2902, n40569, n2903, n40568, n2904, n40567, 
        n1500, n2905, n40566, n1502, n1505, n2906, n40565, n1508, 
        n2907, n40564, n39181, n1409;
    wire [31:0]n1466;
    
    wire n1433, n2908, n40563, n1406, n2909, n40562, n1401, n1407, 
        n1506, n1405, n1504, n1403, n1404, n1402, n1501, n18_adj_4787, 
        n1499, n20_adj_4788, n15, n1507, n1408, n48731, n3083, 
        n40561, n3116;
    wire [31:0]n3149;
    
    wire n3084, n40560, n14, n20_adj_4789, n18_adj_4790, n1598, 
        n22_adj_4791, n1136, n51404, n1109, n34479, n1106, n1103, 
        n1108, n12_adj_4792, n1107, n1105, n1104, n1037, n51403;
    wire [31:0]n971;
    
    wire n2, n50748, n50747, n50764, n28018, n1006, n27973, n1007, 
        n1009, n25164, n1008, n8, n50769, n7, n3085, n40559, 
        n3086, n40558, n3087, n40557, n3088, n40556, n3089, n40555, 
        n3090, n40554, n3091, n40553, n3092, n40552, n3093, n40551, 
        n3094, n40550, n3095, n40549, n39180, n3096, n40548, n4, 
        n39179, n3097, n40547, n39048, n3098, n40546, n3099, n40545, 
        n3100, n40544, n3101, n40543, n3102, n40542, n39047, n3103, 
        n40541, n3104, n40540, n3105, n40539, n1400, n39664, n3106, 
        n40538, n39663, n39662, n3107, n40537, n3108, n40536, 
        n3109, n40535, n39661, n39046, n39660, n39659, n34397, 
        n48, n46, n47, n39658, n45, n39045, n39044, n39657, 
        n44, n39656, n43, n39655, n54, n49, n39163, n39162, 
        n39161, n39160, n26681, n3209, n11_adj_4801, n39159, n27_adj_4802, 
        n23_adj_4803, n39, n33_adj_4804, n13_adj_4805, n1423, n47767, 
        n47771, n47781, n47779, n47793, n25_adj_4806, n31_adj_4807, 
        n47769, n47777, n47773, n47775, n47791, n34429, n26634, 
        n5780, n47797, n47799, n49775, n47801, n47803, n47805, 
        n47807, n47809, n47811, n47813, n59, n61, n41121, n1437, 
        n49782, n44777, n51612, n51528, n50583;
    wire [4:0]color_bit_N_622;
    
    wire n51468, n49792, n51462, n50617;
    wire [3:0]state_3__N_428;
    
    wire n2689;
    wire [31:0]n2753;
    
    wire n2720, n2788, n48994, n48995, n48998, n48997, n48961, 
        n48962, n49022, n49021;
    wire [31:0]n133;
    
    wire n40390, n40389, n40388, n40387, n40386, n40385, n40384, 
        n40383, n40382, n40381, n40380, n40379, n40378, n40377, 
        n40376, n40375, n40374, n40373, n40372, n40371, n40370, 
        n40369, n40833, n40832, n40831, n40830, n40829, n40368, 
        n40828, n40827, n40826, n40825, n40824, n40823, n40822, 
        n40821, n40820, n40819, n40367, n40366, n39425, n40365, 
        n39424, n40818, n40817, n40816, n40815, n40814, n40813, 
        n39423, n40812, n40811, n40810, n40364, n40363, n40809, 
        n40808, n40807, n40806, n40805, n40362, n40804, n39422, 
        n40361, n40803, n40802, n40801, n40800, n40799, n40798, 
        n39421, n40797, n40360, n40796, n39420, n40795, n40794, 
        n40793, n39419, n40792, n40791, n40790, n40789, n40788, 
        n40787, n40786, n40785, n40784, n40783, n40782, n40781, 
        n40780, n40779, n40778, n40777, n40776, n40775, n40774, 
        n40773, n40772, n40771, n40770, n40769, n40768, n40767, 
        n40766, n40765, n40764, n40763, n39418, n40762, n40761, 
        n40760, n40759, n40758, n40757, n2621, n51408, n40756, 
        n40755, n40754, n40753, n40752, n40751, n2192, n40750, 
        n1301, n40359, n39417, n1302, n40358, n1303, n40357;
    wire [31:0]n2159;
    
    wire n40749, n1304, n40356, n40748, n40747, n40746, n1305, 
        n40355, n40745, n40744, n40743, n2707, n2806, n2705, n2804, 
        n2699, n2798, n2706, n2805, n2688, n2787, n2697, n2796, 
        n2696, n2795, n1306, n40354, n2702, n2801, n40742, n39416, 
        n40741, n2698, n2797, n40740, n2701, n2800, n2694, n2793, 
        n40739, n2700, n2799, n2692, n2791, n40738, n2693, n2792, 
        n2691, n2790, n40737, n2690, n2709, n2808, n40736, n2695, 
        n2794, n40735, n2703, n2802, n2708, n2807, n40734, n30_adj_4812, 
        n37, n2291, n40733, n2225, n36;
    wire [31:0]n2258;
    
    wire n2193, n40732, n42, n2704, n40, n2194, n40731, n2687, 
        n41, n39_adj_4813, n2195, n40730, n2809, n2196, n40729, 
        n2803, n30_adj_4814, n2197, n40728, n40_adj_4815, n26_adj_4816, 
        n2198, n40727, n38, n44_adj_4817, n2199, n40726, n42_adj_4818, 
        n2200, n40725, n2201, n40724, n1307, n40353, n2202, n40723, 
        n2203, n40722, n2204, n40721, n39415, n2205, n40720, n2206, 
        n40719, n2207, n40718, n2208, n40717, n1308, n51406, n40352, 
        n2209, n40716, n2390, n40715, n2324;
    wire [31:0]n2357;
    
    wire n2292, n40714, n2293, n40713, n1309, n2294, n40712, n2984, 
        n3017, n40351, n2985, n40350, n2295, n40711, n2296, n40710, 
        n2986, n40349, n2297, n40709, n2298, n40708, n2299, n40707, 
        n2300, n40706, n2301, n40705, n2302, n40704, n2303, n40703, 
        n2304, n40702, n2305, n40701, n2306, n40700, n2307, n40699, 
        n2308, n40698, n2309, n40697, n2489, n40696, n2423;
    wire [31:0]n2456;
    
    wire n2391, n40695, n2392, n40694, n2393, n40693, n2394, n40692, 
        n2395, n40691, n2396, n40690, n2397, n40689, n2987, n40348, 
        n2786, n43_adj_4819, n2398, n40688, n41_adj_4820, n2399, 
        n40687, n2400, n40686, n2401, n40685, n2402, n40684, n2403, 
        n40683, n2404, n40682, n2405, n40681, n2988, n40347, n2406, 
        n40680, n2989, n40346, n2990, n40345, n2407, n40679, n2991, 
        n40344, n2992, n40343, n2993, n40342, n2994, n40341, n2995, 
        n40340, n2996, n40339, n2997, n40338, n2408, n40678, n2998, 
        n40337, n2999, n40336, n3000, n40335, n3001, n40334, n3002, 
        n40333, n3003, n40332, n3004, n40331, n3005, n40330, n2409, 
        n40677, n3006, n40329, n3007, n40328, n3008, n40327, n30593, 
        n51407, n40326, n2588, n40676, n2522, n39074, n39073;
    wire [31:0]n2555;
    
    wire n2490, n40675, n2491, n40674, n2492, n40673, n2493, n40672, 
        n2494, n40671, n2495, n40670, n2496, n40669, n2497, n40668, 
        n2498, n40667, n51609, n48315, n48321, n39072, n2594, 
        n2501, n2600, n2499, n40666, n2500, n40665, n2503, n2602, 
        n2504, n2603, n2505, n2604, n2508, n2607, n2596, n2592, 
        n40664, n2502, n40663, n39071, n40662, n40661, n40660, 
        n2506, n2605, n40659, n2507, n40658, n40657, n2589, n2597, 
        n2509, n40656, n2609, n40655, n40654, n2590, n40653, n2593, 
        n2591, n40652, n2595, n2598, n2606, n39070, n2601, n2608, 
        n39069, n2599, n34, n38_adj_4821, n39068, n29_adj_4822, 
        n36_adj_4823, n44971, n7_adj_4824, n51525, n40651, n35, 
        n39_adj_4825, n41_adj_4826, n40650, n40649, n40648, n40647, 
        n39067, n40646, n40645, n40644, n40643, n40642, n40641, 
        n40640, n40639, n40638, n40637, n39066, n39209, n48313, 
        n40636, n40635, n40634, n39208, n48311, n40633, n40632, 
        n40631, n40630;
    wire [31:0]n1367;
    
    wire n1334, n40629, n40628, n40627, n14_adj_4827, n12_adj_4828, 
        n40626, n40625, n40624, n16_adj_4829, n40623, n40622, n40621, 
        n39065, n12_adj_4830, n16_adj_4831, n17_adj_4832, n40620, 
        n40619, n39207, n48309, n40618, n40617, n40616, n40615, 
        n40614, n40613, n40612, n40611, n2885, n40610, n39064, 
        n40609, n40608, n40607, n40606, n40605, n40604, n40603, 
        n39063, n40602, n40601, n40600, n40599, n40598, n40597, 
        n39206, n48307, n40596, n40595, n40594, n40593, n40592, 
        n40591, n40590, n40589, n40588, n40587, n2886, n40586, 
        n39205, n48305, n39204, n48303, n2918, n39203, n48301, 
        n39062, n51465, n39061, n39060, n39202, n48299, n51459, 
        n39201, n48297, n44847, n44118, n39200, n48295, n39199, 
        n48293, n39198, n48291, n39059, n39058, n39057, n103, 
        n39197, n48289, n16_adj_4833, n6_adj_4834, n40161, n40160, 
        n40159, n40158, n40157, n40156, n40155, n40154, n40153, 
        n39056, n39196, n48287, n39055, n39195, n48285, n39194, 
        n48283, n39193, n48281, n39192, n48279, n39054, n39191, 
        n48277, n39190, n39189, n39188, n46810, n39053, n39187, 
        n39052, n39186, n39051, n39185, n25166, n27979, n36_adj_4837, 
        n46_adj_4838, n42_adj_4839, n32_adj_4840, n22_adj_4841, n28_adj_4842, 
        n44_adj_4843, n50, n36_adj_4844, n34_adj_4845, n33_adj_4846, 
        n48_adj_4847, n49_adj_4848, n37_adj_4849, n39_adj_4850, n47_adj_4851, 
        n26_adj_4852, n34_adj_4853, n32_adj_4854, n31_adj_4855, n35_adj_4856, 
        n37_adj_4857, n32_adj_4858, n42_adj_4859, n38_adj_4860, n43_adj_4861, 
        n40_adj_4862, n46_adj_4863, n39_adj_4864, n47_adj_4865, n44_adj_4866, 
        n42_adj_4867, n43_adj_4868, n41_adj_4869, n40_adj_4870, n39_adj_4871, 
        n50_adj_4872, n45_adj_4873, n30_adj_4874, n34495, n34_adj_4875, 
        n32_adj_4876, n33_adj_4877, n31_adj_4878, n28_adj_4879, n31_adj_4880, 
        n22_adj_4881, n30_adj_4882, n34_adj_4883, n21_adj_4884;
    
    SB_DFF \neo_pixel_transmitter.t0_i0_i1  (.Q(\neo_pixel_transmitter.t0 [1]), 
           .C(CLK_c), .D(n28315));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i2  (.Q(\neo_pixel_transmitter.t0 [2]), 
           .C(CLK_c), .D(n28314));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i3  (.Q(\neo_pixel_transmitter.t0 [3]), 
           .C(CLK_c), .D(n28313));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i4  (.Q(\neo_pixel_transmitter.t0 [4]), 
           .C(CLK_c), .D(n28312));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2009_25_lut (.I0(GND_net), .I1(n2887), .I2(VCC_net), 
            .I3(n40584), .O(n2951[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i9_1_lut (.I0(\neo_pixel_transmitter.t0 [8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[8]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_DFFE \neo_pixel_transmitter.done_104  (.Q(\neo_pixel_transmitter.done ), 
            .C(CLK_c), .E(n51632), .D(\neo_pixel_transmitter.done_N_636 ));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_i1947_3_lut (.I0(n2789), .I1(n2852[28]), .I2(n2819), 
            .I3(GND_net), .O(n2888));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1947_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF \neo_pixel_transmitter.t0_i0_i5  (.Q(\neo_pixel_transmitter.t0 [5]), 
           .C(CLK_c), .D(n28311));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_inv_0_i10_1_lut (.I0(\neo_pixel_transmitter.t0 [9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[9]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \neo_pixel_transmitter.t0_i0_i6  (.Q(\neo_pixel_transmitter.t0 [6]), 
           .C(CLK_c), .D(n28310));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i7  (.Q(\neo_pixel_transmitter.t0 [7]), 
           .C(CLK_c), .D(n28309));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 i35455_4_lut (.I0(n40998), .I1(n44851), .I2(\neo_pixel_transmitter.done ), 
            .I3(\state[0] ), .O(n50261));
    defparam i35455_4_lut.LUT_INIT = 16'hcaaa;
    SB_LUT4 i53_4_lut (.I0(n49769), .I1(n34525), .I2(\state[1] ), .I3(n26525), 
            .O(n44943));
    defparam i53_4_lut.LUT_INIT = 16'hcfca;
    SB_LUT4 i52_4_lut (.I0(n44943), .I1(n50262), .I2(\state[0] ), .I3(\neo_pixel_transmitter.done ), 
            .O(n44987));
    defparam i52_4_lut.LUT_INIT = 16'h3335;
    SB_LUT4 i42_1_lut (.I0(\neo_pixel_transmitter.done ), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_642 ));
    defparam i42_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i4_3_lut (.I0(bit_ctr[23]), .I1(n1203), .I2(n1209), .I3(GND_net), 
            .O(n12));
    defparam i4_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i5_4_lut (.I0(n1208), .I1(n1205), .I2(n1207), .I3(n1204), 
            .O(n13));
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut (.I0(n13), .I1(n1206), .I2(n12), .I3(n1202), .O(n1235));
    defparam i7_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1413_3_lut (.I0(n1999), .I1(n2060[26]), .I2(n2027), 
            .I3(GND_net), .O(n2098));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1413_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1411_3_lut (.I0(n1997), .I1(n2060[28]), .I2(n2027), 
            .I3(GND_net), .O(n2096));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1411_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1412_3_lut (.I0(n1998), .I1(n2060[27]), .I2(n2027), 
            .I3(GND_net), .O(n2097));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1412_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1410_3_lut (.I0(n1996), .I1(n2060[29]), .I2(n2027), 
            .I3(GND_net), .O(n2095));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1410_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1424_3_lut (.I0(bit_ctr[15]), .I1(n2060[15]), .I2(n2027), 
            .I3(GND_net), .O(n2109));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1424_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1423_3_lut (.I0(n2009), .I1(n2060[16]), .I2(n2027), 
            .I3(GND_net), .O(n2108));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1423_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1421_3_lut (.I0(n2007), .I1(n2060[18]), .I2(n2027), 
            .I3(GND_net), .O(n2106));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1421_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1420_3_lut (.I0(n2006), .I1(n2060[19]), .I2(n2027), 
            .I3(GND_net), .O(n2105));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1420_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1422_3_lut (.I0(n2008), .I1(n2060[17]), .I2(n2027), 
            .I3(GND_net), .O(n2107));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1422_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1417_3_lut (.I0(n2003), .I1(n2060[22]), .I2(n2027), 
            .I3(GND_net), .O(n2102));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1417_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1415_3_lut (.I0(n2001), .I1(n2060[24]), .I2(n2027), 
            .I3(GND_net), .O(n2100));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1415_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1416_3_lut (.I0(n2002), .I1(n2060[23]), .I2(n2027), 
            .I3(GND_net), .O(n2101));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1416_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1414_3_lut (.I0(n2000), .I1(n2060[25]), .I2(n2027), 
            .I3(GND_net), .O(n2099));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1414_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1419_3_lut (.I0(n2005), .I1(n2060[20]), .I2(n2027), 
            .I3(GND_net), .O(n2104));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1419_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1418_3_lut (.I0(n2004), .I1(n2060[21]), .I2(n2027), 
            .I3(GND_net), .O(n2103));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1418_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1409_3_lut (.I0(n1995), .I1(n2060[30]), .I2(n2027), 
            .I3(GND_net), .O(n2094));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1409_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut (.I0(n2094), .I1(n2093), .I2(GND_net), .I3(GND_net), 
            .O(n18));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i7_2_lut (.I0(n2103), .I1(n2104), .I2(GND_net), .I3(GND_net), 
            .O(n24_adj_4769));   // verilog/neopixel.v(22[26:36])
    defparam i7_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i13_4_lut (.I0(n2107), .I1(n2105), .I2(n2106), .I3(n18), 
            .O(n30));   // verilog/neopixel.v(22[26:36])
    defparam i13_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(n2099), .I1(n2101), .I2(n2100), .I3(n2102), 
            .O(n28));   // verilog/neopixel.v(22[26:36])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(bit_ctr[14]), .I1(n24_adj_4769), .I2(n2108), 
            .I3(n2109), .O(n29));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut.LUT_INIT = 16'hfefc;
    SB_LUT4 i10_4_lut (.I0(n2095), .I1(n2097), .I2(n2096), .I3(n2098), 
            .O(n27));   // verilog/neopixel.v(22[26:36])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut (.I0(n27), .I1(n29), .I2(n28), .I3(n30), .O(n2126));   // verilog/neopixel.v(22[26:36])
    defparam i16_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i11_1_lut (.I0(\neo_pixel_transmitter.t0 [10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[10]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_DFFESR bit_ctr_i0_i1 (.Q(bit_ctr[1]), .C(CLK_c), .E(n27743), .D(n255[1]), 
            .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i2 (.Q(bit_ctr[2]), .C(CLK_c), .E(n27743), .D(n255[2]), 
            .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i3 (.Q(bit_ctr[3]), .C(CLK_c), .E(n27743), .D(n255[3]), 
            .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i4 (.Q(bit_ctr[4]), .C(CLK_c), .E(n27743), .D(n255[4]), 
            .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i5 (.Q(bit_ctr[5]), .C(CLK_c), .E(n27743), .D(n255[5]), 
            .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i6 (.Q(bit_ctr[6]), .C(CLK_c), .E(n27743), .D(n255[6]), 
            .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i7 (.Q(bit_ctr[7]), .C(CLK_c), .E(n27743), .D(n255[7]), 
            .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i8 (.Q(bit_ctr[8]), .C(CLK_c), .E(n27743), .D(n255[8]), 
            .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i9 (.Q(bit_ctr[9]), .C(CLK_c), .E(n27743), .D(n255[9]), 
            .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i10 (.Q(bit_ctr[10]), .C(CLK_c), .E(n27743), 
            .D(n255[10]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i11 (.Q(bit_ctr[11]), .C(CLK_c), .E(n27743), 
            .D(n255[11]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i12 (.Q(bit_ctr[12]), .C(CLK_c), .E(n27743), 
            .D(n255[12]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i13 (.Q(bit_ctr[13]), .C(CLK_c), .E(n27743), 
            .D(n255[13]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i14 (.Q(bit_ctr[14]), .C(CLK_c), .E(n27743), 
            .D(n255[14]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i15 (.Q(bit_ctr[15]), .C(CLK_c), .E(n27743), 
            .D(n255[15]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i16 (.Q(bit_ctr[16]), .C(CLK_c), .E(n27743), 
            .D(n255[16]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i17 (.Q(bit_ctr[17]), .C(CLK_c), .E(n27743), 
            .D(n255[17]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i18 (.Q(bit_ctr[18]), .C(CLK_c), .E(n27743), 
            .D(n255[18]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i19 (.Q(bit_ctr[19]), .C(CLK_c), .E(n27743), 
            .D(n255[19]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i20 (.Q(bit_ctr[20]), .C(CLK_c), .E(n27743), 
            .D(n255[20]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i21 (.Q(bit_ctr[21]), .C(CLK_c), .E(n27743), 
            .D(n255[21]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i22 (.Q(bit_ctr[22]), .C(CLK_c), .E(n27743), 
            .D(n255[22]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i23 (.Q(bit_ctr[23]), .C(CLK_c), .E(n27743), 
            .D(n255[23]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i24 (.Q(bit_ctr[24]), .C(CLK_c), .E(n27743), 
            .D(n255[24]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i25 (.Q(bit_ctr[25]), .C(CLK_c), .E(n27743), 
            .D(n255[25]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i26 (.Q(bit_ctr[26]), .C(CLK_c), .E(n27743), 
            .D(n255[26]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i27 (.Q(bit_ctr[27]), .C(CLK_c), .E(n27743), 
            .D(n255[27]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i28 (.Q(bit_ctr[28]), .C(CLK_c), .E(n27743), 
            .D(n255[28]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i29 (.Q(bit_ctr[29]), .C(CLK_c), .E(n27743), 
            .D(n255[29]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i30 (.Q(bit_ctr[30]), .C(CLK_c), .E(n27743), 
            .D(n255[30]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFFESR bit_ctr_i0_i31 (.Q(bit_ctr[31]), .C(CLK_c), .E(n27743), 
            .D(n255[31]), .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i8  (.Q(\neo_pixel_transmitter.t0 [8]), 
           .C(CLK_c), .D(n28308));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_2009_25 (.CI(n40584), .I0(n2887), .I1(VCC_net), 
            .CO(n40585));
    SB_LUT4 mod_5_add_2009_24_lut (.I0(GND_net), .I1(n2888), .I2(VCC_net), 
            .I3(n40583), .O(n2951[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_24 (.CI(n40583), .I0(n2888), .I1(VCC_net), 
            .CO(n40584));
    SB_LUT4 mod_5_add_2009_23_lut (.I0(GND_net), .I1(n2889), .I2(VCC_net), 
            .I3(n40582), .O(n2951[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_7_lut (.I0(GND_net), .I1(timer[5]), .I2(n1[5]), 
            .I3(n39183), .O(one_wire_N_579[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_8 (.CI(n39049), .I0(bit_ctr[6]), .I1(GND_net), .CO(n39050));
    SB_LUT4 mod_5_i1356_3_lut (.I0(bit_ctr[16]), .I1(n1961[16]), .I2(n1928), 
            .I3(GND_net), .O(n2009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1344_3_lut (.I0(n1898), .I1(n1961[28]), .I2(n1928), 
            .I3(GND_net), .O(n1997));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1352_3_lut (.I0(n1906), .I1(n1961[20]), .I2(n1928), 
            .I3(GND_net), .O(n2005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1343_3_lut (.I0(n1897), .I1(n1961[29]), .I2(n1928), 
            .I3(GND_net), .O(n1996));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1342_3_lut (.I0(n1896), .I1(n1961[30]), .I2(n1928), 
            .I3(GND_net), .O(n1995));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1342_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_2009_23 (.CI(n40582), .I0(n2889), .I1(VCC_net), 
            .CO(n40583));
    SB_LUT4 mod_5_add_2009_22_lut (.I0(GND_net), .I1(n2890), .I2(VCC_net), 
            .I3(n40581), .O(n2951[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1354_3_lut (.I0(n1908), .I1(n1961[18]), .I2(n1928), 
            .I3(GND_net), .O(n2007));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1354_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1351_3_lut (.I0(n1905), .I1(n1961[21]), .I2(n1928), 
            .I3(GND_net), .O(n2004));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1351_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1355_3_lut (.I0(n1909), .I1(n1961[17]), .I2(n1928), 
            .I3(GND_net), .O(n2008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1350_3_lut (.I0(n1904), .I1(n1961[22]), .I2(n1928), 
            .I3(GND_net), .O(n2003));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1345_3_lut (.I0(n1899), .I1(n1961[27]), .I2(n1928), 
            .I3(GND_net), .O(n1998));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1345_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1353_3_lut (.I0(n1907), .I1(n1961[19]), .I2(n1928), 
            .I3(GND_net), .O(n2006));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1349_3_lut (.I0(n1903), .I1(n1961[23]), .I2(n1928), 
            .I3(GND_net), .O(n2002));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1349_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1348_3_lut (.I0(n1902), .I1(n1961[24]), .I2(n1928), 
            .I3(GND_net), .O(n2001));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1348_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1346_3_lut (.I0(n1900), .I1(n1961[26]), .I2(n1928), 
            .I3(GND_net), .O(n1999));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1347_3_lut (.I0(n1901), .I1(n1961[25]), .I2(n1928), 
            .I3(GND_net), .O(n2000));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1347_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_2_lut (.I0(n2000), .I1(n1999), .I2(GND_net), .I3(GND_net), 
            .O(n20));   // verilog/neopixel.v(22[26:36])
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i12_4_lut_adj_1538 (.I0(n2001), .I1(n2002), .I2(n2006), .I3(n1998), 
            .O(n28_adj_4771));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1538.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut_adj_1539 (.I0(bit_ctr[15]), .I1(n20), .I2(n1997), 
            .I3(n2009), .O(n26));   // verilog/neopixel.v(22[26:36])
    defparam i10_4_lut_adj_1539.LUT_INIT = 16'hfefc;
    SB_LUT4 i11_4_lut_adj_1540 (.I0(n2003), .I1(n2008), .I2(n2004), .I3(n2007), 
            .O(n27_adj_4772));   // verilog/neopixel.v(22[26:36])
    defparam i11_4_lut_adj_1540.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(n1995), .I1(n1996), .I2(n1994), .I3(n2005), 
            .O(n25_adj_4773));   // verilog/neopixel.v(22[26:36])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25_adj_4773), .I1(n27_adj_4772), .I2(n26), 
            .I3(n28_adj_4771), .O(n2027));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1286_3_lut (.I0(n1808), .I1(n1862[19]), .I2(n1829), 
            .I3(GND_net), .O(n1907));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1287_3_lut (.I0(n1809), .I1(n1862[18]), .I2(n1829), 
            .I3(GND_net), .O(n1908));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1287_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1285_3_lut (.I0(n1807), .I1(n1862[20]), .I2(n1829), 
            .I3(GND_net), .O(n1906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1285_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1279_3_lut (.I0(n1801), .I1(n1862[26]), .I2(n1829), 
            .I3(GND_net), .O(n1900));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1279_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1277_3_lut (.I0(n1799), .I1(n1862[28]), .I2(n1829), 
            .I3(GND_net), .O(n1898));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1277_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1278_3_lut (.I0(n1800), .I1(n1862[27]), .I2(n1829), 
            .I3(GND_net), .O(n1899));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1278_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1276_3_lut (.I0(n1798), .I1(n1862[29]), .I2(n1829), 
            .I3(GND_net), .O(n1897));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1276_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1275_3_lut (.I0(n1797), .I1(n1862[30]), .I2(n1829), 
            .I3(GND_net), .O(n1896));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1275_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1283_3_lut (.I0(n1805), .I1(n1862[22]), .I2(n1829), 
            .I3(GND_net), .O(n1904));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1283_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1281_3_lut (.I0(n1803), .I1(n1862[24]), .I2(n1829), 
            .I3(GND_net), .O(n1902));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1281_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1282_3_lut (.I0(n1804), .I1(n1862[23]), .I2(n1829), 
            .I3(GND_net), .O(n1903));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1282_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1280_3_lut (.I0(n1802), .I1(n1862[25]), .I2(n1829), 
            .I3(GND_net), .O(n1901));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1288_3_lut (.I0(bit_ctr[17]), .I1(n1862[17]), .I2(n1829), 
            .I3(GND_net), .O(n1909));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1284_3_lut (.I0(n1806), .I1(n1862[21]), .I2(n1829), 
            .I3(GND_net), .O(n1905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1284_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_3_lut (.I0(bit_ctr[16]), .I1(n1905), .I2(n1909), .I3(GND_net), 
            .O(n21));   // verilog/neopixel.v(22[26:36])
    defparam i6_3_lut.LUT_INIT = 16'hecec;
    SB_CARRY sub_14_add_2_7 (.CI(n39183), .I0(timer[5]), .I1(n1[5]), .CO(n39184));
    SB_CARRY mod_5_add_2009_22 (.CI(n40581), .I0(n2890), .I1(VCC_net), 
            .CO(n40582));
    SB_LUT4 mod_5_add_2009_21_lut (.I0(GND_net), .I1(n2891), .I2(VCC_net), 
            .I3(n40580), .O(n2951[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i10_4_lut_adj_1541 (.I0(n1901), .I1(n1903), .I2(n1902), .I3(n1904), 
            .O(n25_adj_4774));   // verilog/neopixel.v(22[26:36])
    defparam i10_4_lut_adj_1541.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1542 (.I0(n1896), .I1(n1895), .I2(GND_net), .I3(GND_net), 
            .O(n16));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_adj_1542.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1543 (.I0(n1897), .I1(n1899), .I2(n1898), .I3(n1900), 
            .O(n24_adj_4775));   // verilog/neopixel.v(22[26:36])
    defparam i9_4_lut_adj_1543.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1544 (.I0(n25_adj_4774), .I1(n21), .I2(n1906), 
            .I3(n1908), .O(n28_adj_4776));   // verilog/neopixel.v(22[26:36])
    defparam i13_4_lut_adj_1544.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut (.I0(n1907), .I1(n28_adj_4776), .I2(n24_adj_4775), 
            .I3(n16), .O(n1928));   // verilog/neopixel.v(22[26:36])
    defparam i14_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2009_21 (.CI(n40580), .I0(n2891), .I1(VCC_net), 
            .CO(n40581));
    SB_LUT4 i21422_2_lut (.I0(bit_ctr[17]), .I1(n1809), .I2(GND_net), 
            .I3(GND_net), .O(n34485));
    defparam i21422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mod_5_add_2009_20_lut (.I0(GND_net), .I1(n2892), .I2(VCC_net), 
            .I3(n40579), .O(n2951[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_2_lut_adj_1545 (.I0(n1800), .I1(n1801), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4777));   // verilog/neopixel.v(22[26:36])
    defparam i4_2_lut_adj_1545.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1546 (.I0(n1803), .I1(n1804), .I2(n1808), .I3(n1807), 
            .O(n24_adj_4778));   // verilog/neopixel.v(22[26:36])
    defparam i10_4_lut_adj_1546.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(n1797), .I1(n1806), .I2(n1796), .I3(n34485), 
            .O(n22));   // verilog/neopixel.v(22[26:36])
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_add_2_6_lut (.I0(GND_net), .I1(timer[4]), .I2(n1[4]), 
            .I3(n39182), .O(one_wire_N_579[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_20 (.CI(n40579), .I0(n2892), .I1(VCC_net), 
            .CO(n40580));
    SB_CARRY sub_14_add_2_6 (.CI(n39182), .I0(timer[4]), .I1(n1[4]), .CO(n39183));
    SB_LUT4 i12_4_lut_adj_1547 (.I0(n1798), .I1(n24_adj_4778), .I2(n18_adj_4777), 
            .I3(n1799), .O(n26_adj_4780));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1547.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1548 (.I0(n1802), .I1(n26_adj_4780), .I2(n22), 
            .I3(n1805), .O(n1829));   // verilog/neopixel.v(22[26:36])
    defparam i13_4_lut_adj_1548.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2009_19_lut (.I0(GND_net), .I1(n2893), .I2(VCC_net), 
            .I3(n40578), .O(n2951[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_19 (.CI(n40578), .I0(n2893), .I1(VCC_net), 
            .CO(n40579));
    SB_LUT4 mod_5_add_2009_18_lut (.I0(GND_net), .I1(n2894), .I2(VCC_net), 
            .I3(n40577), .O(n2951[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_18_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i9  (.Q(\neo_pixel_transmitter.t0 [9]), 
           .C(CLK_c), .D(n28307));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_2009_18 (.CI(n40577), .I0(n2894), .I1(VCC_net), 
            .CO(n40578));
    SB_LUT4 i36452_1_lut (.I0(n1730), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51405));
    defparam i36452_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i1142_3_lut (.I0(n1600), .I1(n1664[29]), .I2(n1631), 
            .I3(GND_net), .O(n1699));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1142_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1145_3_lut (.I0(n1603), .I1(n1664[26]), .I2(n1631), 
            .I3(GND_net), .O(n1702));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1145_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1141_3_lut (.I0(n1599), .I1(n1664[30]), .I2(n1631), 
            .I3(GND_net), .O(n1698));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1141_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1152_3_lut (.I0(bit_ctr[19]), .I1(n1664[19]), .I2(n1631), 
            .I3(GND_net), .O(n1709));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1152_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1151_3_lut (.I0(n1609), .I1(n1664[20]), .I2(n1631), 
            .I3(GND_net), .O(n1708));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1151_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1144_3_lut (.I0(n1602), .I1(n1664[27]), .I2(n1631), 
            .I3(GND_net), .O(n1701));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1144_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1148_3_lut (.I0(n1606), .I1(n1664[23]), .I2(n1631), 
            .I3(GND_net), .O(n1705));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1148_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1147_3_lut (.I0(n1605), .I1(n1664[24]), .I2(n1631), 
            .I3(GND_net), .O(n1704));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1149_3_lut (.I0(n1607), .I1(n1664[22]), .I2(n1631), 
            .I3(GND_net), .O(n1706));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1149_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1143_3_lut (.I0(n1601), .I1(n1664[28]), .I2(n1631), 
            .I3(GND_net), .O(n1700));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1143_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_2009_17_lut (.I0(GND_net), .I1(n2895), .I2(VCC_net), 
            .I3(n40576), .O(n2951[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1150_3_lut (.I0(n1608), .I1(n1664[21]), .I2(n1631), 
            .I3(GND_net), .O(n1707));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1150_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1146_3_lut (.I0(n1604), .I1(n1664[25]), .I2(n1631), 
            .I3(GND_net), .O(n1703));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i3_2_lut (.I0(n1703), .I1(n1707), .I2(GND_net), .I3(GND_net), 
            .O(n16_adj_4781));
    defparam i3_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i9_4_lut_adj_1549 (.I0(n1700), .I1(n1706), .I2(n1704), .I3(n1705), 
            .O(n22_adj_4782));
    defparam i9_4_lut_adj_1549.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_1550 (.I0(n1701), .I1(bit_ctr[18]), .I2(n1708), 
            .I3(n1709), .O(n20_adj_4783));
    defparam i7_4_lut_adj_1550.LUT_INIT = 16'hfefa;
    SB_LUT4 i11_4_lut_adj_1551 (.I0(n1698), .I1(n22_adj_4782), .I2(n16_adj_4781), 
            .I3(n1702), .O(n24_adj_4784));
    defparam i11_4_lut_adj_1551.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1552 (.I0(n1699), .I1(n24_adj_4784), .I2(n20_adj_4783), 
            .I3(n1697), .O(n1730));
    defparam i12_4_lut_adj_1552.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2009_17 (.CI(n40576), .I0(n2895), .I1(VCC_net), 
            .CO(n40577));
    SB_LUT4 mod_5_add_2009_16_lut (.I0(GND_net), .I1(n2896), .I2(VCC_net), 
            .I3(n40575), .O(n2951[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_16 (.CI(n40575), .I0(n2896), .I1(VCC_net), 
            .CO(n40576));
    SB_LUT4 mod_5_add_2009_15_lut (.I0(GND_net), .I1(n2897), .I2(VCC_net), 
            .I3(n40574), .O(n2951[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_15 (.CI(n40574), .I0(n2897), .I1(VCC_net), 
            .CO(n40575));
    SB_LUT4 mod_5_add_2009_14_lut (.I0(GND_net), .I1(n2898), .I2(VCC_net), 
            .I3(n40573), .O(n2951[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_14 (.CI(n40573), .I0(n2898), .I1(VCC_net), 
            .CO(n40574));
    SB_DFF \neo_pixel_transmitter.t0_i0_i10  (.Q(\neo_pixel_transmitter.t0 [10]), 
           .C(CLK_c), .D(n28306));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i11  (.Q(\neo_pixel_transmitter.t0 [11]), 
           .C(CLK_c), .D(n28305));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2009_13_lut (.I0(GND_net), .I1(n2899), .I2(VCC_net), 
            .I3(n40572), .O(n2951[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_13 (.CI(n40572), .I0(n2899), .I1(VCC_net), 
            .CO(n40573));
    SB_LUT4 mod_5_add_2009_12_lut (.I0(GND_net), .I1(n2900), .I2(VCC_net), 
            .I3(n40571), .O(n2951[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_12 (.CI(n40571), .I0(n2900), .I1(VCC_net), 
            .CO(n40572));
    SB_LUT4 mod_5_add_2009_11_lut (.I0(GND_net), .I1(n2901), .I2(VCC_net), 
            .I3(n40570), .O(n2951[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_11 (.CI(n40570), .I0(n2901), .I1(VCC_net), 
            .CO(n40571));
    SB_LUT4 sub_14_inv_0_i12_1_lut (.I0(\neo_pixel_transmitter.t0 [11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[11]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_DFF \neo_pixel_transmitter.t0_i0_i12  (.Q(\neo_pixel_transmitter.t0 [12]), 
           .C(CLK_c), .D(n28304));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i13  (.Q(\neo_pixel_transmitter.t0 [13]), 
           .C(CLK_c), .D(n28303));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_i1083_3_lut (.I0(n1509), .I1(n1565[21]), .I2(n1532), 
            .I3(GND_net), .O(n1608));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1083_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1077_3_lut (.I0(n1503), .I1(n1565[27]), .I2(n1532), 
            .I3(GND_net), .O(n1602));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1077_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_2009_10_lut (.I0(GND_net), .I1(n2902), .I2(VCC_net), 
            .I3(n40569), .O(n2951[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_10 (.CI(n40569), .I0(n2902), .I1(VCC_net), 
            .CO(n40570));
    SB_LUT4 mod_5_add_2009_9_lut (.I0(GND_net), .I1(n2903), .I2(VCC_net), 
            .I3(n40568), .O(n2951[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_9 (.CI(n40568), .I0(n2903), .I1(VCC_net), 
            .CO(n40569));
    SB_LUT4 mod_5_add_2009_8_lut (.I0(GND_net), .I1(n2904), .I2(VCC_net), 
            .I3(n40567), .O(n2951[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1074_3_lut (.I0(n1500), .I1(n1565[30]), .I2(n1532), 
            .I3(GND_net), .O(n1599));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1074_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_2009_8 (.CI(n40567), .I0(n2904), .I1(VCC_net), 
            .CO(n40568));
    SB_LUT4 mod_5_add_2009_7_lut (.I0(GND_net), .I1(n2905), .I2(VCC_net), 
            .I3(n40566), .O(n2951[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_7 (.CI(n40566), .I0(n2905), .I1(VCC_net), 
            .CO(n40567));
    SB_LUT4 mod_5_i1076_3_lut (.I0(n1502), .I1(n1565[28]), .I2(n1532), 
            .I3(GND_net), .O(n1601));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1076_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1079_3_lut (.I0(n1505), .I1(n1565[25]), .I2(n1532), 
            .I3(GND_net), .O(n1604));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1079_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1084_3_lut (.I0(bit_ctr[20]), .I1(n1565[20]), .I2(n1532), 
            .I3(GND_net), .O(n1609));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1084_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF \neo_pixel_transmitter.t0_i0_i14  (.Q(\neo_pixel_transmitter.t0 [14]), 
           .C(CLK_c), .D(n28302));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2009_6_lut (.I0(GND_net), .I1(n2906), .I2(VCC_net), 
            .I3(n40565), .O(n2951[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1082_3_lut (.I0(n1508), .I1(n1565[22]), .I2(n1532), 
            .I3(GND_net), .O(n1607));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1082_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_2009_6 (.CI(n40565), .I0(n2906), .I1(VCC_net), 
            .CO(n40566));
    SB_LUT4 mod_5_add_2009_5_lut (.I0(GND_net), .I1(n2907), .I2(VCC_net), 
            .I3(n40564), .O(n2951[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_5 (.CI(n40564), .I0(n2907), .I1(VCC_net), 
            .CO(n40565));
    SB_LUT4 sub_14_add_2_5_lut (.I0(GND_net), .I1(timer[3]), .I2(n1[3]), 
            .I3(n39181), .O(one_wire_N_579[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1015_3_lut (.I0(n1409), .I1(n1466[22]), .I2(n1433), 
            .I3(GND_net), .O(n1508));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1016_3_lut (.I0(bit_ctr[21]), .I1(n1466[21]), .I2(n1433), 
            .I3(GND_net), .O(n1509));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_2009_4_lut (.I0(GND_net), .I1(n2908), .I2(VCC_net), 
            .I3(n40563), .O(n2951[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_4 (.CI(n40563), .I0(n2908), .I1(VCC_net), 
            .CO(n40564));
    SB_LUT4 mod_5_i1012_3_lut (.I0(n1406), .I1(n1466[25]), .I2(n1433), 
            .I3(GND_net), .O(n1505));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_2009_3_lut (.I0(GND_net), .I1(n2909), .I2(GND_net), 
            .I3(n40562), .O(n2951[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_3 (.CI(n40562), .I0(n2909), .I1(GND_net), 
            .CO(n40563));
    SB_LUT4 mod_5_i1007_3_lut (.I0(n1401), .I1(n1466[30]), .I2(n1433), 
            .I3(GND_net), .O(n1500));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1007_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1013_3_lut (.I0(n1407), .I1(n1466[24]), .I2(n1433), 
            .I3(GND_net), .O(n1506));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1011_3_lut (.I0(n1405), .I1(n1466[26]), .I2(n1433), 
            .I3(GND_net), .O(n1504));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1011_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1009_3_lut (.I0(n1403), .I1(n1466[28]), .I2(n1433), 
            .I3(GND_net), .O(n1502));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1010_3_lut (.I0(n1404), .I1(n1466[27]), .I2(n1433), 
            .I3(GND_net), .O(n1503));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1008_3_lut (.I0(n1402), .I1(n1466[29]), .I2(n1433), 
            .I3(GND_net), .O(n1501));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1008_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_4_lut_adj_1553 (.I0(n1501), .I1(n1503), .I2(n1502), .I3(n1504), 
            .O(n18_adj_4787));
    defparam i7_4_lut_adj_1553.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2009_2_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(VCC_net), .O(n2951[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i9_4_lut_adj_1554 (.I0(n1506), .I1(n18_adj_4787), .I2(n1500), 
            .I3(n1499), .O(n20_adj_4788));
    defparam i9_4_lut_adj_1554.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_2009_2 (.CI(VCC_net), .I0(bit_ctr[6]), .I1(GND_net), 
            .CO(n40562));
    SB_LUT4 i4_3_lut_adj_1555 (.I0(n1505), .I1(bit_ctr[20]), .I2(n1509), 
            .I3(GND_net), .O(n15));
    defparam i4_3_lut_adj_1555.LUT_INIT = 16'heaea;
    SB_LUT4 i10_4_lut_adj_1556 (.I0(n15), .I1(n20_adj_4788), .I2(n1507), 
            .I3(n1508), .O(n1532));
    defparam i10_4_lut_adj_1556.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1014_3_lut (.I0(n1408), .I1(n1466[23]), .I2(n1433), 
            .I3(GND_net), .O(n1507));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1081_3_lut (.I0(n1507), .I1(n1565[23]), .I2(n1532), 
            .I3(GND_net), .O(n1606));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1081_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_2143_29_lut (.I0(n3116), .I1(n3083), .I2(VCC_net), 
            .I3(n40561), .O(n48731)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_29_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_i1080_3_lut (.I0(n1506), .I1(n1565[24]), .I2(n1532), 
            .I3(GND_net), .O(n1605));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1080_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1078_3_lut (.I0(n1504), .I1(n1565[26]), .I2(n1532), 
            .I3(GND_net), .O(n1603));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1078_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_2143_28_lut (.I0(GND_net), .I1(n3084), .I2(VCC_net), 
            .I3(n40560), .O(n3149[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_28 (.CI(n40560), .I0(n3084), .I1(VCC_net), 
            .CO(n40561));
    SB_LUT4 mod_5_i1075_3_lut (.I0(n1501), .I1(n1565[29]), .I2(n1532), 
            .I3(GND_net), .O(n1600));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1075_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut (.I0(bit_ctr[19]), .I1(n1607), .I2(n1609), .I3(GND_net), 
            .O(n14));   // verilog/neopixel.v(22[26:36])
    defparam i2_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 i8_4_lut_adj_1557 (.I0(n1600), .I1(n1603), .I2(n1605), .I3(n1606), 
            .O(n20_adj_4789));   // verilog/neopixel.v(22[26:36])
    defparam i8_4_lut_adj_1557.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_2_lut (.I0(n1604), .I1(n1601), .I2(GND_net), .I3(GND_net), 
            .O(n18_adj_4790));   // verilog/neopixel.v(22[26:36])
    defparam i6_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i10_4_lut_adj_1558 (.I0(n1599), .I1(n20_adj_4789), .I2(n14), 
            .I3(n1598), .O(n22_adj_4791));   // verilog/neopixel.v(22[26:36])
    defparam i10_4_lut_adj_1558.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1559 (.I0(n1602), .I1(n22_adj_4791), .I2(n18_adj_4790), 
            .I3(n1608), .O(n1631));   // verilog/neopixel.v(22[26:36])
    defparam i11_4_lut_adj_1559.LUT_INIT = 16'hfffe;
    SB_LUT4 i36451_1_lut (.I0(n1136), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51404));
    defparam i36451_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21416_2_lut (.I0(bit_ctr[24]), .I1(n1109), .I2(GND_net), 
            .I3(GND_net), .O(n34479));
    defparam i21416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut_adj_1560 (.I0(n1106), .I1(n1103), .I2(n1108), .I3(n34479), 
            .O(n12_adj_4792));
    defparam i5_4_lut_adj_1560.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(n1107), .I1(n12_adj_4792), .I2(n1105), .I3(n1104), 
            .O(n1136));
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i36450_1_lut (.I0(n1037), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51403));
    defparam i36450_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i35795_2_lut (.I0(n971[28]), .I1(n2), .I2(GND_net), .I3(GND_net), 
            .O(n50748));   // verilog/neopixel.v(22[26:36])
    defparam i35795_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i35794_2_lut (.I0(n971[29]), .I1(n2), .I2(GND_net), .I3(GND_net), 
            .O(n50747));   // verilog/neopixel.v(22[26:36])
    defparam i35794_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i35811_2_lut (.I0(n971[30]), .I1(n2), .I2(GND_net), .I3(GND_net), 
            .O(n50764));   // verilog/neopixel.v(22[26:36])
    defparam i35811_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 mod_5_i673_3_lut (.I0(n28018), .I1(n971[29]), .I2(n2), .I3(GND_net), 
            .O(n1006));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i673_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i674_3_lut (.I0(n27973), .I1(n971[28]), .I2(n2), .I3(GND_net), 
            .O(n1007));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i674_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i676_3_lut (.I0(bit_ctr[26]), .I1(n971[26]), .I2(n2), 
            .I3(GND_net), .O(n1009));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i676_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 mod_5_i675_3_lut (.I0(n25164), .I1(n971[27]), .I2(n2), .I3(GND_net), 
            .O(n1008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i675_3_lut.LUT_INIT = 16'hacac;
    SB_LUT4 i2_2_lut_3_lut (.I0(n1007), .I1(n971[30]), .I2(n2), .I3(GND_net), 
            .O(n8));
    defparam i2_2_lut_3_lut.LUT_INIT = 16'haeae;
    SB_LUT4 i35816_2_lut (.I0(n971[31]), .I1(n2), .I2(GND_net), .I3(GND_net), 
            .O(n50769));   // verilog/neopixel.v(22[26:36])
    defparam i35816_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut (.I0(n1008), .I1(bit_ctr[25]), .I2(n1009), .I3(GND_net), 
            .O(n7));
    defparam i1_3_lut.LUT_INIT = 16'heaea;
    SB_LUT4 i5_4_lut_adj_1561 (.I0(n50769), .I1(n7), .I2(n1006), .I3(n8), 
            .O(n1037));
    defparam i5_4_lut_adj_1561.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_2143_27_lut (.I0(GND_net), .I1(n3085), .I2(VCC_net), 
            .I3(n40559), .O(n3149[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_27 (.CI(n40559), .I0(n3085), .I1(VCC_net), 
            .CO(n40560));
    SB_LUT4 mod_5_add_2143_26_lut (.I0(GND_net), .I1(n3086), .I2(VCC_net), 
            .I3(n40558), .O(n3149[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_26_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i15  (.Q(\neo_pixel_transmitter.t0 [15]), 
           .C(CLK_c), .D(n28301));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_2143_26 (.CI(n40558), .I0(n3086), .I1(VCC_net), 
            .CO(n40559));
    SB_LUT4 mod_5_add_2143_25_lut (.I0(GND_net), .I1(n3087), .I2(VCC_net), 
            .I3(n40557), .O(n3149[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_25 (.CI(n40557), .I0(n3087), .I1(VCC_net), 
            .CO(n40558));
    SB_LUT4 mod_5_add_2143_24_lut (.I0(GND_net), .I1(n3088), .I2(VCC_net), 
            .I3(n40556), .O(n3149[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_24 (.CI(n40556), .I0(n3088), .I1(VCC_net), 
            .CO(n40557));
    SB_LUT4 mod_5_add_2143_23_lut (.I0(GND_net), .I1(n3089), .I2(VCC_net), 
            .I3(n40555), .O(n3149[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_23 (.CI(n40555), .I0(n3089), .I1(VCC_net), 
            .CO(n40556));
    SB_LUT4 mod_5_add_2143_22_lut (.I0(GND_net), .I1(n3090), .I2(VCC_net), 
            .I3(n40554), .O(n3149[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_22 (.CI(n40554), .I0(n3090), .I1(VCC_net), 
            .CO(n40555));
    SB_LUT4 mod_5_add_2143_21_lut (.I0(GND_net), .I1(n3091), .I2(VCC_net), 
            .I3(n40553), .O(n3149[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_21 (.CI(n40553), .I0(n3091), .I1(VCC_net), 
            .CO(n40554));
    SB_LUT4 mod_5_add_2143_20_lut (.I0(GND_net), .I1(n3092), .I2(VCC_net), 
            .I3(n40552), .O(n3149[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_20 (.CI(n40552), .I0(n3092), .I1(VCC_net), 
            .CO(n40553));
    SB_LUT4 mod_5_add_2143_19_lut (.I0(GND_net), .I1(n3093), .I2(VCC_net), 
            .I3(n40551), .O(n3149[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_5 (.CI(n39181), .I0(timer[3]), .I1(n1[3]), .CO(n39182));
    SB_CARRY mod_5_add_2143_19 (.CI(n40551), .I0(n3093), .I1(VCC_net), 
            .CO(n40552));
    SB_LUT4 mod_5_add_2143_18_lut (.I0(GND_net), .I1(n3094), .I2(VCC_net), 
            .I3(n40550), .O(n3149[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_18 (.CI(n40550), .I0(n3094), .I1(VCC_net), 
            .CO(n40551));
    SB_LUT4 mod_5_add_2143_17_lut (.I0(GND_net), .I1(n3095), .I2(VCC_net), 
            .I3(n40549), .O(n3149[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_17 (.CI(n40549), .I0(n3095), .I1(VCC_net), 
            .CO(n40550));
    SB_LUT4 sub_14_add_2_4_lut (.I0(GND_net), .I1(timer[2]), .I2(n1[2]), 
            .I3(n39180), .O(one_wire_N_579[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2143_16_lut (.I0(GND_net), .I1(n3096), .I2(VCC_net), 
            .I3(n40548), .O(n3149[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_16 (.CI(n40548), .I0(n3096), .I1(VCC_net), 
            .CO(n40549));
    SB_LUT4 sub_14_inv_0_i13_1_lut (.I0(\neo_pixel_transmitter.t0 [12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[12]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY sub_14_add_2_4 (.CI(n39180), .I0(timer[2]), .I1(n1[2]), .CO(n39181));
    SB_LUT4 sub_14_add_2_3_lut (.I0(one_wire_N_579[3]), .I1(timer[1]), .I2(n1[1]), 
            .I3(n39179), .O(n4)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_3_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2143_15_lut (.I0(GND_net), .I1(n3097), .I2(VCC_net), 
            .I3(n40547), .O(n3149[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_7_lut (.I0(GND_net), .I1(bit_ctr[5]), .I2(GND_net), 
            .I3(n39048), .O(n255[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_7 (.CI(n39048), .I0(bit_ctr[5]), .I1(GND_net), .CO(n39049));
    SB_LUT4 sub_14_inv_0_i14_1_lut (.I0(\neo_pixel_transmitter.t0 [13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[13]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i15_1_lut (.I0(\neo_pixel_transmitter.t0 [14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[14]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2143_15 (.CI(n40547), .I0(n3097), .I1(VCC_net), 
            .CO(n40548));
    SB_LUT4 mod_5_add_2143_14_lut (.I0(GND_net), .I1(n3098), .I2(VCC_net), 
            .I3(n40546), .O(n3149[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_14 (.CI(n40546), .I0(n3098), .I1(VCC_net), 
            .CO(n40547));
    SB_LUT4 mod_5_add_2143_13_lut (.I0(GND_net), .I1(n3099), .I2(VCC_net), 
            .I3(n40545), .O(n3149[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_13 (.CI(n40545), .I0(n3099), .I1(VCC_net), 
            .CO(n40546));
    SB_LUT4 sub_14_inv_0_i16_1_lut (.I0(\neo_pixel_transmitter.t0 [15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[15]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i17_1_lut (.I0(\neo_pixel_transmitter.t0 [16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[16]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2143_12_lut (.I0(GND_net), .I1(n3100), .I2(VCC_net), 
            .I3(n40544), .O(n3149[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_12 (.CI(n40544), .I0(n3100), .I1(VCC_net), 
            .CO(n40545));
    SB_LUT4 mod_5_add_2143_11_lut (.I0(GND_net), .I1(n3101), .I2(VCC_net), 
            .I3(n40543), .O(n3149[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_11 (.CI(n40543), .I0(n3101), .I1(VCC_net), 
            .CO(n40544));
    SB_DFF \neo_pixel_transmitter.t0_i0_i16  (.Q(\neo_pixel_transmitter.t0 [16]), 
           .C(CLK_c), .D(n28300));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2143_10_lut (.I0(GND_net), .I1(n3102), .I2(VCC_net), 
            .I3(n40542), .O(n3149[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_3 (.CI(n39179), .I0(timer[1]), .I1(n1[1]), .CO(n39180));
    SB_CARRY sub_14_add_2_2 (.CI(VCC_net), .I0(timer[0]), .I1(n1[0]), 
            .CO(n39179));
    SB_LUT4 add_21_6_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(n39047), .O(n255[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_10 (.CI(n40542), .I0(n3102), .I1(VCC_net), 
            .CO(n40543));
    SB_DFF \neo_pixel_transmitter.t0_i0_i17  (.Q(\neo_pixel_transmitter.t0 [17]), 
           .C(CLK_c), .D(n28299));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_2143_9_lut (.I0(GND_net), .I1(n3103), .I2(VCC_net), 
            .I3(n40541), .O(n3149[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_9 (.CI(n40541), .I0(n3103), .I1(VCC_net), 
            .CO(n40542));
    SB_LUT4 mod_5_add_2143_8_lut (.I0(GND_net), .I1(n3104), .I2(VCC_net), 
            .I3(n40540), .O(n3149[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_8 (.CI(n40540), .I0(n3104), .I1(VCC_net), 
            .CO(n40541));
    SB_LUT4 mod_5_add_2143_7_lut (.I0(GND_net), .I1(n3105), .I2(VCC_net), 
            .I3(n40539), .O(n3149[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_7_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i18  (.Q(\neo_pixel_transmitter.t0 [18]), 
           .C(CLK_c), .D(n28298));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_1004_12_lut (.I0(n1433), .I1(n1400), .I2(VCC_net), 
            .I3(n39664), .O(n1499)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 sub_14_inv_0_i18_1_lut (.I0(\neo_pixel_transmitter.t0 [17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[17]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_2143_7 (.CI(n40539), .I0(n3105), .I1(VCC_net), 
            .CO(n40540));
    SB_LUT4 mod_5_add_2143_6_lut (.I0(GND_net), .I1(n3106), .I2(VCC_net), 
            .I3(n40538), .O(n3149[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_6 (.CI(n40538), .I0(n3106), .I1(VCC_net), 
            .CO(n40539));
    SB_LUT4 sub_14_inv_0_i19_1_lut (.I0(\neo_pixel_transmitter.t0 [18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[18]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1004_11_lut (.I0(GND_net), .I1(n1401), .I2(VCC_net), 
            .I3(n39663), .O(n1466[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_11 (.CI(n39663), .I0(n1401), .I1(VCC_net), 
            .CO(n39664));
    SB_LUT4 mod_5_add_1004_10_lut (.I0(GND_net), .I1(n1402), .I2(VCC_net), 
            .I3(n39662), .O(n1466[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2143_5_lut (.I0(GND_net), .I1(n3107), .I2(VCC_net), 
            .I3(n40537), .O(n3149[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_10 (.CI(n39662), .I0(n1402), .I1(VCC_net), 
            .CO(n39663));
    SB_CARRY mod_5_add_2143_5 (.CI(n40537), .I0(n3107), .I1(VCC_net), 
            .CO(n40538));
    SB_LUT4 mod_5_add_2143_4_lut (.I0(GND_net), .I1(n3108), .I2(VCC_net), 
            .I3(n40536), .O(n3149[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_4 (.CI(n40536), .I0(n3108), .I1(VCC_net), 
            .CO(n40537));
    SB_LUT4 mod_5_add_2143_3_lut (.I0(GND_net), .I1(n3109), .I2(GND_net), 
            .I3(n40535), .O(n3149[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_3 (.CI(n40535), .I0(n3109), .I1(GND_net), 
            .CO(n40536));
    SB_LUT4 mod_5_add_1004_9_lut (.I0(GND_net), .I1(n1403), .I2(VCC_net), 
            .I3(n39661), .O(n1466[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_9 (.CI(n39661), .I0(n1403), .I1(VCC_net), 
            .CO(n39662));
    SB_CARRY add_21_6 (.CI(n39047), .I0(bit_ctr[4]), .I1(GND_net), .CO(n39048));
    SB_LUT4 mod_5_add_2143_2_lut (.I0(GND_net), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(VCC_net), .O(n3149[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2143_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2143_2 (.CI(VCC_net), .I0(bit_ctr[4]), .I1(GND_net), 
            .CO(n40535));
    SB_DFF \neo_pixel_transmitter.t0_i0_i19  (.Q(\neo_pixel_transmitter.t0 [19]), 
           .C(CLK_c), .D(n28297));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_5_lut (.I0(GND_net), .I1(bit_ctr[3]), .I2(GND_net), 
            .I3(n39046), .O(n255[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1004_8_lut (.I0(GND_net), .I1(n1404), .I2(VCC_net), 
            .I3(n39660), .O(n1466[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_8 (.CI(n39660), .I0(n1404), .I1(VCC_net), 
            .CO(n39661));
    SB_LUT4 mod_5_add_1004_7_lut (.I0(GND_net), .I1(n1405), .I2(VCC_net), 
            .I3(n39659), .O(n1466[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_7 (.CI(n39659), .I0(n1405), .I1(VCC_net), 
            .CO(n39660));
    SB_LUT4 i21337_2_lut (.I0(bit_ctr[3]), .I1(bit_ctr[4]), .I2(GND_net), 
            .I3(GND_net), .O(n34397));
    defparam i21337_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20_4_lut (.I0(bit_ctr[8]), .I1(bit_ctr[18]), .I2(bit_ctr[24]), 
            .I3(bit_ctr[9]), .O(n48));
    defparam i20_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_21_5 (.CI(n39046), .I0(bit_ctr[3]), .I1(GND_net), .CO(n39047));
    SB_LUT4 i18_4_lut (.I0(bit_ctr[26]), .I1(bit_ctr[28]), .I2(bit_ctr[6]), 
            .I3(bit_ctr[19]), .O(n46));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(bit_ctr[13]), .I1(bit_ctr[20]), .I2(bit_ctr[23]), 
            .I3(bit_ctr[16]), .O(n47));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1004_6_lut (.I0(GND_net), .I1(n1406), .I2(VCC_net), 
            .I3(n39658), .O(n1466[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17_4_lut (.I0(bit_ctr[15]), .I1(bit_ctr[14]), .I2(bit_ctr[21]), 
            .I3(bit_ctr[22]), .O(n45));
    defparam i17_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF \neo_pixel_transmitter.t0_i0_i20  (.Q(\neo_pixel_transmitter.t0 [20]), 
           .C(CLK_c), .D(n28296));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i21  (.Q(\neo_pixel_transmitter.t0 [21]), 
           .C(CLK_c), .D(n28295));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i22  (.Q(\neo_pixel_transmitter.t0 [22]), 
           .C(CLK_c), .D(n28294));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_4_lut (.I0(GND_net), .I1(bit_ctr[2]), .I2(GND_net), 
            .I3(n39045), .O(n255[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_6 (.CI(n39658), .I0(n1406), .I1(VCC_net), 
            .CO(n39659));
    SB_CARRY add_21_4 (.CI(n39045), .I0(bit_ctr[2]), .I1(GND_net), .CO(n39046));
    SB_LUT4 add_21_3_lut (.I0(GND_net), .I1(bit_ctr[1]), .I2(GND_net), 
            .I3(n39044), .O(n255[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1004_5_lut (.I0(GND_net), .I1(n1407), .I2(VCC_net), 
            .I3(n39657), .O(n1466[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16_4_lut_adj_1562 (.I0(bit_ctr[11]), .I1(bit_ctr[7]), .I2(bit_ctr[17]), 
            .I3(bit_ctr[29]), .O(n44));
    defparam i16_4_lut_adj_1562.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1004_5 (.CI(n39657), .I0(n1407), .I1(VCC_net), 
            .CO(n39658));
    SB_LUT4 mod_5_add_1004_4_lut (.I0(GND_net), .I1(n1408), .I2(VCC_net), 
            .I3(n39656), .O(n1466[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_4_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i23  (.Q(\neo_pixel_transmitter.t0 [23]), 
           .C(CLK_c), .D(n28293));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i24  (.Q(\neo_pixel_transmitter.t0 [24]), 
           .C(CLK_c), .D(n28292));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i25  (.Q(\neo_pixel_transmitter.t0 [25]), 
           .C(CLK_c), .D(n28291));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i26  (.Q(\neo_pixel_transmitter.t0 [26]), 
           .C(CLK_c), .D(n28290));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i27  (.Q(\neo_pixel_transmitter.t0 [27]), 
           .C(CLK_c), .D(n28289));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY mod_5_add_1004_4 (.CI(n39656), .I0(n1408), .I1(VCC_net), 
            .CO(n39657));
    SB_LUT4 i15_4_lut_adj_1563 (.I0(bit_ctr[12]), .I1(bit_ctr[30]), .I2(n34397), 
            .I3(bit_ctr[25]), .O(n43));
    defparam i15_4_lut_adj_1563.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1004_3_lut (.I0(GND_net), .I1(n1409), .I2(GND_net), 
            .I3(n39655), .O(n1466[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_3 (.CI(n39044), .I0(bit_ctr[1]), .I1(GND_net), .CO(n39045));
    SB_CARRY mod_5_add_1004_3 (.CI(n39655), .I0(n1409), .I1(GND_net), 
            .CO(n39656));
    SB_LUT4 mod_5_add_1004_2_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(VCC_net), .O(n1466[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1004_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1004_2 (.CI(VCC_net), .I0(bit_ctr[21]), .I1(GND_net), 
            .CO(n39655));
    SB_LUT4 add_21_2_lut (.I0(GND_net), .I1(bit_ctr[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n255[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_2_lut.LUT_INIT = 16'hC33C;
    SB_DFF \neo_pixel_transmitter.t0_i0_i28  (.Q(\neo_pixel_transmitter.t0 [28]), 
           .C(CLK_c), .D(n28288));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i29  (.Q(\neo_pixel_transmitter.t0 [29]), 
           .C(CLK_c), .D(n28287));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i30  (.Q(\neo_pixel_transmitter.t0 [30]), 
           .C(CLK_c), .D(n28286));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i31  (.Q(\neo_pixel_transmitter.t0 [31]), 
           .C(CLK_c), .D(n28285));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_2 (.CI(VCC_net), .I0(bit_ctr[0]), .I1(GND_net), .CO(n39044));
    SB_LUT4 i26_4_lut (.I0(n45), .I1(n47), .I2(n46), .I3(n48), .O(n54));
    defparam i26_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 sub_14_inv_0_i20_1_lut (.I0(\neo_pixel_transmitter.t0 [19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[19]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21_4_lut (.I0(bit_ctr[27]), .I1(bit_ctr[31]), .I2(bit_ctr[10]), 
            .I3(bit_ctr[5]), .O(n49));
    defparam i21_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_669_7_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n39163), .O(n971[31])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_669_6_lut (.I0(GND_net), .I1(GND_net), .I2(VCC_net), 
            .I3(n39162), .O(n971[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i21_1_lut (.I0(\neo_pixel_transmitter.t0 [20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[20]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_669_6 (.CI(n39162), .I0(GND_net), .I1(VCC_net), 
            .CO(n39163));
    SB_LUT4 mod_5_add_669_5_lut (.I0(GND_net), .I1(n28018), .I2(VCC_net), 
            .I3(n39161), .O(n971[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_669_5 (.CI(n39161), .I0(n28018), .I1(VCC_net), 
            .CO(n39162));
    SB_LUT4 sub_14_inv_0_i22_1_lut (.I0(\neo_pixel_transmitter.t0 [21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[21]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_669_4_lut (.I0(GND_net), .I1(n27973), .I2(VCC_net), 
            .I3(n39160), .O(n971[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i23_1_lut (.I0(\neo_pixel_transmitter.t0 [22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[22]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i21462_4_lut (.I0(one_wire_N_579[8]), .I1(n26681), .I2(one_wire_N_579[10]), 
            .I3(one_wire_N_579[9]), .O(n34525));
    defparam i21462_4_lut.LUT_INIT = 16'hfcec;
    SB_LUT4 mod_5_i2172_3_lut (.I0(bit_ctr[4]), .I1(n3149[4]), .I2(n3116), 
            .I3(GND_net), .O(n3209));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2172_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_669_4 (.CI(n39160), .I0(n27973), .I1(VCC_net), 
            .CO(n39161));
    SB_LUT4 mod_5_i2171_3_lut (.I0(n3109), .I1(n3149[5]), .I2(n3116), 
            .I3(GND_net), .O(n11_adj_4801));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2171_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_669_3_lut (.I0(GND_net), .I1(n25164), .I2(GND_net), 
            .I3(n39159), .O(n971[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i2163_3_lut (.I0(n3101), .I1(n3149[13]), .I2(n3116), 
            .I3(GND_net), .O(n27_adj_4802));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2163_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2165_3_lut (.I0(n3103), .I1(n3149[11]), .I2(n3116), 
            .I3(GND_net), .O(n23_adj_4803));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2165_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_669_3 (.CI(n39159), .I0(n25164), .I1(GND_net), 
            .CO(n39160));
    SB_LUT4 mod_5_i2157_3_lut (.I0(n3095), .I1(n3149[19]), .I2(n3116), 
            .I3(GND_net), .O(n39));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2157_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2160_3_lut (.I0(n3098), .I1(n3149[16]), .I2(n3116), 
            .I3(GND_net), .O(n33_adj_4804));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2160_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2170_3_lut (.I0(n3108), .I1(n3149[6]), .I2(n3116), 
            .I3(GND_net), .O(n13_adj_4805));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2170_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_669_2_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(VCC_net), .O(n971[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_669_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i27_4_lut (.I0(n49), .I1(n54), .I2(n43), .I3(n44), .O(\state_3__N_428[1] ));
    defparam i27_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i277_2_lut (.I0(LED_c), .I1(\state_3__N_428[1] ), .I2(GND_net), 
            .I3(GND_net), .O(n1423));   // verilog/neopixel.v(40[18] 45[12])
    defparam i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(n3106), .I1(n11_adj_4801), .I2(n3149[8]), .I3(n3116), 
            .O(n47767));
    defparam i1_4_lut.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1564 (.I0(n3096), .I1(n13_adj_4805), .I2(n3149[18]), 
            .I3(n3116), .O(n47771));
    defparam i1_4_lut_adj_1564.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1565 (.I0(n3100), .I1(n33_adj_4804), .I2(n3149[14]), 
            .I3(n3116), .O(n47781));
    defparam i1_4_lut_adj_1565.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1566 (.I0(n3105), .I1(n39), .I2(n3149[9]), .I3(n3116), 
            .O(n47779));
    defparam i1_4_lut_adj_1566.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1567 (.I0(n47779), .I1(n47781), .I2(n47771), 
            .I3(n47767), .O(n47793));
    defparam i1_4_lut_adj_1567.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i2164_3_lut (.I0(n3102), .I1(n3149[12]), .I2(n3116), 
            .I3(GND_net), .O(n25_adj_4806));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2164_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2161_3_lut (.I0(n3099), .I1(n3149[15]), .I2(n3116), 
            .I3(GND_net), .O(n31_adj_4807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2161_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1568 (.I0(n3107), .I1(n27_adj_4802), .I2(n3149[7]), 
            .I3(n3116), .O(n47769));
    defparam i1_4_lut_adj_1568.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1569 (.I0(n3097), .I1(n23_adj_4803), .I2(n3149[17]), 
            .I3(n3116), .O(n47777));
    defparam i1_4_lut_adj_1569.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1570 (.I0(n3104), .I1(n31_adj_4807), .I2(n3149[10]), 
            .I3(n3116), .O(n47773));
    defparam i1_4_lut_adj_1570.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1571 (.I0(n3094), .I1(n25_adj_4806), .I2(n3149[20]), 
            .I3(n3116), .O(n47775));
    defparam i1_4_lut_adj_1571.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1572 (.I0(n47775), .I1(n47773), .I2(n47777), 
            .I3(n47769), .O(n47791));
    defparam i1_4_lut_adj_1572.LUT_INIT = 16'hfffe;
    SB_LUT4 i3799_4_lut (.I0(n34429), .I1(n1423), .I2(\state[1] ), .I3(n26634), 
            .O(n5780));
    defparam i3799_4_lut.LUT_INIT = 16'h3f35;
    SB_LUT4 i1_4_lut_adj_1573 (.I0(n3093), .I1(n47793), .I2(n3149[21]), 
            .I3(n3116), .O(n47797));
    defparam i1_4_lut_adj_1573.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1574 (.I0(n47797), .I1(n47791), .I2(bit_ctr[3]), 
            .I3(n3209), .O(n47799));
    defparam i1_4_lut_adj_1574.LUT_INIT = 16'hfeee;
    SB_LUT4 i34906_3_lut (.I0(n40998), .I1(n26634), .I2(n26525), .I3(GND_net), 
            .O(n49775));
    defparam i34906_3_lut.LUT_INIT = 16'hcdcd;
    SB_LUT4 i36443_4_lut (.I0(\state[1] ), .I1(n49775), .I2(n5780), .I3(\state[0] ), 
            .O(n27743));
    defparam i36443_4_lut.LUT_INIT = 16'h0f11;
    SB_LUT4 i1_4_lut_adj_1575 (.I0(n3092), .I1(n47799), .I2(n3149[22]), 
            .I3(n3116), .O(n47801));
    defparam i1_4_lut_adj_1575.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1576 (.I0(n3091), .I1(n47801), .I2(n3149[23]), 
            .I3(n3116), .O(n47803));
    defparam i1_4_lut_adj_1576.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1577 (.I0(n3090), .I1(n47803), .I2(n3149[24]), 
            .I3(n3116), .O(n47805));
    defparam i1_4_lut_adj_1577.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1578 (.I0(n3089), .I1(n47805), .I2(n3149[25]), 
            .I3(n3116), .O(n47807));
    defparam i1_4_lut_adj_1578.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1579 (.I0(n3088), .I1(n47807), .I2(n3149[26]), 
            .I3(n3116), .O(n47809));
    defparam i1_4_lut_adj_1579.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1580 (.I0(n3087), .I1(n47809), .I2(n3149[27]), 
            .I3(n3116), .O(n47811));
    defparam i1_4_lut_adj_1580.LUT_INIT = 16'hfcee;
    SB_LUT4 i1_4_lut_adj_1581 (.I0(n3086), .I1(n47811), .I2(n3149[28]), 
            .I3(n3116), .O(n47813));
    defparam i1_4_lut_adj_1581.LUT_INIT = 16'hfcee;
    SB_LUT4 mod_5_i2147_3_lut (.I0(n3085), .I1(n3149[29]), .I2(n3116), 
            .I3(GND_net), .O(n59));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2147_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2146_3_lut (.I0(n3084), .I1(n3149[30]), .I2(n3116), 
            .I3(GND_net), .O(n61));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2146_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1582 (.I0(n61), .I1(n48731), .I2(n59), .I3(n47813), 
            .O(n41121));
    defparam i1_4_lut_adj_1582.LUT_INIT = 16'hfffe;
    SB_LUT4 i291_2_lut (.I0(n34525), .I1(\neo_pixel_transmitter.done ), 
            .I2(GND_net), .I3(GND_net), .O(n1437));   // verilog/neopixel.v(103[9] 111[12])
    defparam i291_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i15_4_lut_adj_1583 (.I0(n34629), .I1(n49782), .I2(\state[1] ), 
            .I3(n26634), .O(n44839));   // verilog/neopixel.v(35[12] 117[6])
    defparam i15_4_lut_adj_1583.LUT_INIT = 16'h303a;
    SB_LUT4 i1_4_lut_adj_1584 (.I0(\state[1] ), .I1(n44777), .I2(n1437), 
            .I3(\state[0] ), .O(n27916));
    defparam i1_4_lut_adj_1584.LUT_INIT = 16'hee4e;
    SB_LUT4 i35630_3_lut (.I0(n51612), .I1(n51528), .I2(bit_ctr[2]), .I3(GND_net), 
            .O(n50583));
    defparam i35630_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35138_3_lut (.I0(n3209), .I1(bit_ctr[3]), .I2(n41121), .I3(GND_net), 
            .O(color_bit_N_622[4]));
    defparam i35138_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i35259_3_lut (.I0(n51468), .I1(bit_ctr[3]), .I2(n41121), .I3(GND_net), 
            .O(n49792));
    defparam i35259_3_lut.LUT_INIT = 16'h8282;
    SB_LUT4 i35664_4_lut (.I0(n50583), .I1(n51462), .I2(bit_ctr[3]), .I3(n41121), 
            .O(n50617));   // verilog/neopixel.v(22[26:36])
    defparam i35664_4_lut.LUT_INIT = 16'hacca;
    SB_LUT4 i20561_4_lut (.I0(n50617), .I1(\state_3__N_428[1] ), .I2(n49792), 
            .I3(color_bit_N_622[4]), .O(state_3__N_428[0]));   // verilog/neopixel.v(40[18] 45[12])
    defparam i20561_4_lut.LUT_INIT = 16'h3022;
    SB_CARRY mod_5_add_669_2 (.CI(VCC_net), .I0(bit_ctr[26]), .I1(GND_net), 
            .CO(n39159));
    SB_LUT4 sub_14_inv_0_i24_1_lut (.I0(\neo_pixel_transmitter.t0 [23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[23]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i1879_3_lut (.I0(n2689), .I1(n2753[29]), .I2(n2720), 
            .I3(GND_net), .O(n2788));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1879_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1946_3_lut (.I0(n2788), .I1(n2852[29]), .I2(n2819), 
            .I3(GND_net), .O(n2887));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34042_3_lut (.I0(neopxl_color[8]), .I1(neopxl_color[9]), .I2(bit_ctr[0]), 
            .I3(GND_net), .O(n48994));
    defparam i34042_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34043_3_lut (.I0(neopxl_color[10]), .I1(neopxl_color[11]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n48995));
    defparam i34043_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34046_3_lut (.I0(neopxl_color[14]), .I1(neopxl_color[15]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n48998));
    defparam i34046_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34045_3_lut (.I0(neopxl_color[12]), .I1(neopxl_color[13]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n48997));
    defparam i34045_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_inv_0_i25_1_lut (.I0(\neo_pixel_transmitter.t0 [24]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[24]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i25_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i34009_3_lut (.I0(neopxl_color[16]), .I1(neopxl_color[17]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n48961));
    defparam i34009_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34010_3_lut (.I0(neopxl_color[18]), .I1(neopxl_color[19]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n48962));
    defparam i34010_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34070_3_lut (.I0(neopxl_color[22]), .I1(neopxl_color[23]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n49022));
    defparam i34070_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34069_3_lut (.I0(neopxl_color[20]), .I1(neopxl_color[21]), 
            .I2(bit_ctr[0]), .I3(GND_net), .O(n49021));
    defparam i34069_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_inv_0_i26_1_lut (.I0(\neo_pixel_transmitter.t0 [25]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[25]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i26_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i27_1_lut (.I0(\neo_pixel_transmitter.t0 [26]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[26]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i27_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_1546_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(timer[31]), 
            .I3(n40390), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1546_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(timer[30]), 
            .I3(n40389), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_32 (.CI(n40389), .I0(GND_net), .I1(timer[30]), 
            .CO(n40390));
    SB_LUT4 timer_1546_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(timer[29]), 
            .I3(n40388), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_31 (.CI(n40388), .I0(GND_net), .I1(timer[29]), 
            .CO(n40389));
    SB_LUT4 timer_1546_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(timer[28]), 
            .I3(n40387), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_30 (.CI(n40387), .I0(GND_net), .I1(timer[28]), 
            .CO(n40388));
    SB_LUT4 timer_1546_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(timer[27]), 
            .I3(n40386), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_29 (.CI(n40386), .I0(GND_net), .I1(timer[27]), 
            .CO(n40387));
    SB_LUT4 timer_1546_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(timer[26]), 
            .I3(n40385), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_28 (.CI(n40385), .I0(GND_net), .I1(timer[26]), 
            .CO(n40386));
    SB_LUT4 timer_1546_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(timer[25]), 
            .I3(n40384), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_27 (.CI(n40384), .I0(GND_net), .I1(timer[25]), 
            .CO(n40385));
    SB_LUT4 timer_1546_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(timer[24]), 
            .I3(n40383), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_26 (.CI(n40383), .I0(GND_net), .I1(timer[24]), 
            .CO(n40384));
    SB_LUT4 timer_1546_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(timer[23]), 
            .I3(n40382), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_25 (.CI(n40382), .I0(GND_net), .I1(timer[23]), 
            .CO(n40383));
    SB_LUT4 timer_1546_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(timer[22]), 
            .I3(n40381), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_24 (.CI(n40381), .I0(GND_net), .I1(timer[22]), 
            .CO(n40382));
    SB_LUT4 timer_1546_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(timer[21]), 
            .I3(n40380), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_23 (.CI(n40380), .I0(GND_net), .I1(timer[21]), 
            .CO(n40381));
    SB_LUT4 timer_1546_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(timer[20]), 
            .I3(n40379), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i28_1_lut (.I0(\neo_pixel_transmitter.t0 [27]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[27]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i28_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY timer_1546_add_4_22 (.CI(n40379), .I0(GND_net), .I1(timer[20]), 
            .CO(n40380));
    SB_LUT4 timer_1546_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(timer[19]), 
            .I3(n40378), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_21 (.CI(n40378), .I0(GND_net), .I1(timer[19]), 
            .CO(n40379));
    SB_LUT4 timer_1546_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(timer[18]), 
            .I3(n40377), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_20 (.CI(n40377), .I0(GND_net), .I1(timer[18]), 
            .CO(n40378));
    SB_LUT4 timer_1546_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(timer[17]), 
            .I3(n40376), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_19 (.CI(n40376), .I0(GND_net), .I1(timer[17]), 
            .CO(n40377));
    SB_LUT4 timer_1546_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(timer[16]), 
            .I3(n40375), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_18 (.CI(n40375), .I0(GND_net), .I1(timer[16]), 
            .CO(n40376));
    SB_LUT4 timer_1546_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(timer[15]), 
            .I3(n40374), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_17 (.CI(n40374), .I0(GND_net), .I1(timer[15]), 
            .CO(n40375));
    SB_LUT4 timer_1546_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(timer[14]), 
            .I3(n40373), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_16 (.CI(n40373), .I0(GND_net), .I1(timer[14]), 
            .CO(n40374));
    SB_LUT4 timer_1546_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(timer[13]), 
            .I3(n40372), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_15 (.CI(n40372), .I0(GND_net), .I1(timer[13]), 
            .CO(n40373));
    SB_LUT4 timer_1546_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(timer[12]), 
            .I3(n40371), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_14 (.CI(n40371), .I0(GND_net), .I1(timer[12]), 
            .CO(n40372));
    SB_LUT4 timer_1546_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(timer[11]), 
            .I3(n40370), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_13 (.CI(n40370), .I0(GND_net), .I1(timer[11]), 
            .CO(n40371));
    SB_LUT4 timer_1546_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(timer[10]), 
            .I3(n40369), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_12 (.CI(n40369), .I0(GND_net), .I1(timer[10]), 
            .CO(n40370));
    SB_LUT4 sub_14_inv_0_i29_1_lut (.I0(\neo_pixel_transmitter.t0 [28]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[28]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i29_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_736_8_lut (.I0(n50769), .I1(n50769), .I2(n1037), 
            .I3(n40833), .O(n1103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_736_7_lut (.I0(n50764), .I1(n50764), .I2(n1037), 
            .I3(n40832), .O(n1104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_7 (.CI(n40832), .I0(n50764), .I1(n1037), .CO(n40833));
    SB_LUT4 mod_5_add_736_6_lut (.I0(n50747), .I1(n1006), .I2(n1037), 
            .I3(n40831), .O(n1105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_6 (.CI(n40831), .I0(n1006), .I1(n1037), .CO(n40832));
    SB_LUT4 mod_5_add_736_5_lut (.I0(n50748), .I1(n1007), .I2(n1037), 
            .I3(n40830), .O(n1106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_736_5 (.CI(n40830), .I0(n1007), .I1(n1037), .CO(n40831));
    SB_LUT4 mod_5_add_736_4_lut (.I0(n1008), .I1(n1008), .I2(n1037), .I3(n40829), 
            .O(n1107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 timer_1546_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(timer[9]), 
            .I3(n40368), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_11 (.CI(n40368), .I0(GND_net), .I1(timer[9]), 
            .CO(n40369));
    SB_CARRY mod_5_add_736_4 (.CI(n40829), .I0(n1008), .I1(n1037), .CO(n40830));
    SB_LUT4 mod_5_add_736_3_lut (.I0(n1009), .I1(n1009), .I2(n51403), 
            .I3(n40828), .O(n1108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_3 (.CI(n40828), .I0(n1009), .I1(n51403), .CO(n40829));
    SB_LUT4 mod_5_add_736_2_lut (.I0(bit_ctr[25]), .I1(bit_ctr[25]), .I2(n51403), 
            .I3(VCC_net), .O(n1109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_736_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_736_2 (.CI(VCC_net), .I0(bit_ctr[25]), .I1(n51403), 
            .CO(n40828));
    SB_LUT4 mod_5_add_803_9_lut (.I0(n1103), .I1(n1103), .I2(n1136), .I3(n40827), 
            .O(n1202)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_9_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_803_8_lut (.I0(n1104), .I1(n1104), .I2(n1136), .I3(n40826), 
            .O(n1203)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_8 (.CI(n40826), .I0(n1104), .I1(n1136), .CO(n40827));
    SB_LUT4 mod_5_add_803_7_lut (.I0(n1105), .I1(n1105), .I2(n1136), .I3(n40825), 
            .O(n1204)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_7 (.CI(n40825), .I0(n1105), .I1(n1136), .CO(n40826));
    SB_LUT4 mod_5_add_803_6_lut (.I0(n1106), .I1(n1106), .I2(n1136), .I3(n40824), 
            .O(n1205)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_6 (.CI(n40824), .I0(n1106), .I1(n1136), .CO(n40825));
    SB_LUT4 mod_5_add_803_5_lut (.I0(n1107), .I1(n1107), .I2(n1136), .I3(n40823), 
            .O(n1206)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_5 (.CI(n40823), .I0(n1107), .I1(n1136), .CO(n40824));
    SB_LUT4 mod_5_add_803_4_lut (.I0(n1108), .I1(n1108), .I2(n1136), .I3(n40822), 
            .O(n1207)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_803_4 (.CI(n40822), .I0(n1108), .I1(n1136), .CO(n40823));
    SB_LUT4 mod_5_add_803_3_lut (.I0(n1109), .I1(n1109), .I2(n51404), 
            .I3(n40821), .O(n1208)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_3 (.CI(n40821), .I0(n1109), .I1(n51404), .CO(n40822));
    SB_LUT4 mod_5_add_803_2_lut (.I0(bit_ctr[24]), .I1(bit_ctr[24]), .I2(n51404), 
            .I3(VCC_net), .O(n1209)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_803_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_803_2 (.CI(VCC_net), .I0(bit_ctr[24]), .I1(n51404), 
            .CO(n40821));
    SB_LUT4 mod_5_add_1138_14_lut (.I0(n1631), .I1(n1598), .I2(VCC_net), 
            .I3(n40820), .O(n1697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1138_13_lut (.I0(GND_net), .I1(n1599), .I2(VCC_net), 
            .I3(n40819), .O(n1664[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1546_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(timer[8]), 
            .I3(n40367), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_10 (.CI(n40367), .I0(GND_net), .I1(timer[8]), 
            .CO(n40368));
    SB_LUT4 timer_1546_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(timer[7]), 
            .I3(n40366), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_13_lut (.I0(n1532), .I1(n1499), .I2(VCC_net), 
            .I3(n39425), .O(n1598)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_13_lut.LUT_INIT = 16'h8228;
    SB_CARRY timer_1546_add_4_9 (.CI(n40366), .I0(GND_net), .I1(timer[7]), 
            .CO(n40367));
    SB_LUT4 timer_1546_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(timer[6]), 
            .I3(n40365), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_12_lut (.I0(GND_net), .I1(n1500), .I2(VCC_net), 
            .I3(n39424), .O(n1565[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_13 (.CI(n40819), .I0(n1599), .I1(VCC_net), 
            .CO(n40820));
    SB_CARRY mod_5_add_1071_12 (.CI(n39424), .I0(n1500), .I1(VCC_net), 
            .CO(n39425));
    SB_LUT4 mod_5_add_1138_12_lut (.I0(GND_net), .I1(n1600), .I2(VCC_net), 
            .I3(n40818), .O(n1664[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_12 (.CI(n40818), .I0(n1600), .I1(VCC_net), 
            .CO(n40819));
    SB_LUT4 mod_5_add_1138_11_lut (.I0(GND_net), .I1(n1601), .I2(VCC_net), 
            .I3(n40817), .O(n1664[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_11 (.CI(n40817), .I0(n1601), .I1(VCC_net), 
            .CO(n40818));
    SB_LUT4 mod_5_add_1138_10_lut (.I0(GND_net), .I1(n1602), .I2(VCC_net), 
            .I3(n40816), .O(n1664[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_10 (.CI(n40816), .I0(n1602), .I1(VCC_net), 
            .CO(n40817));
    SB_LUT4 mod_5_add_1138_9_lut (.I0(GND_net), .I1(n1603), .I2(VCC_net), 
            .I3(n40815), .O(n1664[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_9 (.CI(n40815), .I0(n1603), .I1(VCC_net), 
            .CO(n40816));
    SB_LUT4 mod_5_add_1138_8_lut (.I0(GND_net), .I1(n1604), .I2(VCC_net), 
            .I3(n40814), .O(n1664[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_8 (.CI(n40814), .I0(n1604), .I1(VCC_net), 
            .CO(n40815));
    SB_LUT4 mod_5_add_1138_7_lut (.I0(GND_net), .I1(n1605), .I2(VCC_net), 
            .I3(n40813), .O(n1664[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_7 (.CI(n40813), .I0(n1605), .I1(VCC_net), 
            .CO(n40814));
    SB_LUT4 mod_5_add_1071_11_lut (.I0(GND_net), .I1(n1501), .I2(VCC_net), 
            .I3(n39423), .O(n1565[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_11 (.CI(n39423), .I0(n1501), .I1(VCC_net), 
            .CO(n39424));
    SB_LUT4 mod_5_add_1138_6_lut (.I0(GND_net), .I1(n1606), .I2(VCC_net), 
            .I3(n40812), .O(n1664[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_6 (.CI(n40812), .I0(n1606), .I1(VCC_net), 
            .CO(n40813));
    SB_LUT4 mod_5_add_1138_5_lut (.I0(GND_net), .I1(n1607), .I2(VCC_net), 
            .I3(n40811), .O(n1664[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_8 (.CI(n40365), .I0(GND_net), .I1(timer[6]), 
            .CO(n40366));
    SB_CARRY mod_5_add_1138_5 (.CI(n40811), .I0(n1607), .I1(VCC_net), 
            .CO(n40812));
    SB_LUT4 mod_5_add_1138_4_lut (.I0(GND_net), .I1(n1608), .I2(VCC_net), 
            .I3(n40810), .O(n1664[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 timer_1546_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(timer[5]), 
            .I3(n40364), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_7 (.CI(n40364), .I0(GND_net), .I1(timer[5]), 
            .CO(n40365));
    SB_LUT4 timer_1546_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(timer[4]), 
            .I3(n40363), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_4 (.CI(n40810), .I0(n1608), .I1(VCC_net), 
            .CO(n40811));
    SB_CARRY timer_1546_add_4_6 (.CI(n40363), .I0(GND_net), .I1(timer[4]), 
            .CO(n40364));
    SB_LUT4 mod_5_add_1138_3_lut (.I0(GND_net), .I1(n1609), .I2(GND_net), 
            .I3(n40809), .O(n1664[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_3 (.CI(n40809), .I0(n1609), .I1(GND_net), 
            .CO(n40810));
    SB_LUT4 mod_5_add_1138_2_lut (.I0(GND_net), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(VCC_net), .O(n1664[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1138_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1138_2 (.CI(VCC_net), .I0(bit_ctr[19]), .I1(GND_net), 
            .CO(n40809));
    SB_LUT4 mod_5_add_1205_15_lut (.I0(n1697), .I1(n1697), .I2(n1730), 
            .I3(n40808), .O(n1796)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_15_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1205_14_lut (.I0(n1698), .I1(n1698), .I2(n1730), 
            .I3(n40807), .O(n1797)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_14 (.CI(n40807), .I0(n1698), .I1(n1730), .CO(n40808));
    SB_LUT4 mod_5_add_1205_13_lut (.I0(n1699), .I1(n1699), .I2(n1730), 
            .I3(n40806), .O(n1798)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_13 (.CI(n40806), .I0(n1699), .I1(n1730), .CO(n40807));
    SB_LUT4 mod_5_add_1205_12_lut (.I0(n1700), .I1(n1700), .I2(n1730), 
            .I3(n40805), .O(n1799)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_12 (.CI(n40805), .I0(n1700), .I1(n1730), .CO(n40806));
    SB_LUT4 timer_1546_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(timer[3]), 
            .I3(n40362), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1205_11_lut (.I0(n1701), .I1(n1701), .I2(n1730), 
            .I3(n40804), .O(n1800)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_11_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1071_10_lut (.I0(GND_net), .I1(n1502), .I2(VCC_net), 
            .I3(n39422), .O(n1565[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_5 (.CI(n40362), .I0(GND_net), .I1(timer[3]), 
            .CO(n40363));
    SB_CARRY mod_5_add_1205_11 (.CI(n40804), .I0(n1701), .I1(n1730), .CO(n40805));
    SB_LUT4 timer_1546_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(timer[2]), 
            .I3(n40361), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1205_10_lut (.I0(n1702), .I1(n1702), .I2(n1730), 
            .I3(n40803), .O(n1801)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_10 (.CI(n39422), .I0(n1502), .I1(VCC_net), 
            .CO(n39423));
    SB_CARRY mod_5_add_1205_10 (.CI(n40803), .I0(n1702), .I1(n1730), .CO(n40804));
    SB_LUT4 mod_5_add_1205_9_lut (.I0(n1703), .I1(n1703), .I2(n1730), 
            .I3(n40802), .O(n1802)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_9 (.CI(n40802), .I0(n1703), .I1(n1730), .CO(n40803));
    SB_LUT4 mod_5_add_1205_8_lut (.I0(n1704), .I1(n1704), .I2(n1730), 
            .I3(n40801), .O(n1803)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_8 (.CI(n40801), .I0(n1704), .I1(n1730), .CO(n40802));
    SB_LUT4 mod_5_add_1205_7_lut (.I0(n1705), .I1(n1705), .I2(n1730), 
            .I3(n40800), .O(n1804)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_7 (.CI(n40800), .I0(n1705), .I1(n1730), .CO(n40801));
    SB_LUT4 mod_5_add_1205_6_lut (.I0(n1706), .I1(n1706), .I2(n1730), 
            .I3(n40799), .O(n1805)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_6 (.CI(n40799), .I0(n1706), .I1(n1730), .CO(n40800));
    SB_LUT4 mod_5_add_1205_5_lut (.I0(n1707), .I1(n1707), .I2(n1730), 
            .I3(n40798), .O(n1806)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1205_5 (.CI(n40798), .I0(n1707), .I1(n1730), .CO(n40799));
    SB_LUT4 mod_5_add_1071_9_lut (.I0(GND_net), .I1(n1503), .I2(VCC_net), 
            .I3(n39421), .O(n1565[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY timer_1546_add_4_4 (.CI(n40361), .I0(GND_net), .I1(timer[2]), 
            .CO(n40362));
    SB_LUT4 mod_5_add_1205_4_lut (.I0(n1708), .I1(n1708), .I2(n1730), 
            .I3(n40797), .O(n1807)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_9 (.CI(n39421), .I0(n1503), .I1(VCC_net), 
            .CO(n39422));
    SB_CARRY mod_5_add_1205_4 (.CI(n40797), .I0(n1708), .I1(n1730), .CO(n40798));
    SB_LUT4 timer_1546_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(timer[1]), 
            .I3(n40360), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1205_3_lut (.I0(n1709), .I1(n1709), .I2(n51405), 
            .I3(n40796), .O(n1808)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_3 (.CI(n40796), .I0(n1709), .I1(n51405), .CO(n40797));
    SB_LUT4 mod_5_add_1071_8_lut (.I0(GND_net), .I1(n1504), .I2(VCC_net), 
            .I3(n39420), .O(n1565[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1205_2_lut (.I0(bit_ctr[18]), .I1(bit_ctr[18]), .I2(n51405), 
            .I3(VCC_net), .O(n1809)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1205_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1205_2 (.CI(VCC_net), .I0(bit_ctr[18]), .I1(n51405), 
            .CO(n40796));
    SB_LUT4 mod_5_add_1272_16_lut (.I0(n1829), .I1(n1796), .I2(VCC_net), 
            .I3(n40795), .O(n1895)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1272_15_lut (.I0(GND_net), .I1(n1797), .I2(VCC_net), 
            .I3(n40794), .O(n1862[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_8 (.CI(n39420), .I0(n1504), .I1(VCC_net), 
            .CO(n39421));
    SB_CARRY mod_5_add_1272_15 (.CI(n40794), .I0(n1797), .I1(VCC_net), 
            .CO(n40795));
    SB_LUT4 mod_5_add_1272_14_lut (.I0(GND_net), .I1(n1798), .I2(VCC_net), 
            .I3(n40793), .O(n1862[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_14 (.CI(n40793), .I0(n1798), .I1(VCC_net), 
            .CO(n40794));
    SB_LUT4 mod_5_add_1071_7_lut (.I0(GND_net), .I1(n1505), .I2(VCC_net), 
            .I3(n39419), .O(n1565[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1272_13_lut (.I0(GND_net), .I1(n1799), .I2(VCC_net), 
            .I3(n40792), .O(n1862[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_13 (.CI(n40792), .I0(n1799), .I1(VCC_net), 
            .CO(n40793));
    SB_LUT4 mod_5_add_1272_12_lut (.I0(GND_net), .I1(n1800), .I2(VCC_net), 
            .I3(n40791), .O(n1862[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_12 (.CI(n40791), .I0(n1800), .I1(VCC_net), 
            .CO(n40792));
    SB_LUT4 mod_5_add_1272_11_lut (.I0(GND_net), .I1(n1801), .I2(VCC_net), 
            .I3(n40790), .O(n1862[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_11 (.CI(n40790), .I0(n1801), .I1(VCC_net), 
            .CO(n40791));
    SB_LUT4 mod_5_add_1272_10_lut (.I0(GND_net), .I1(n1802), .I2(VCC_net), 
            .I3(n40789), .O(n1862[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_10 (.CI(n40789), .I0(n1802), .I1(VCC_net), 
            .CO(n40790));
    SB_LUT4 mod_5_add_1272_9_lut (.I0(GND_net), .I1(n1803), .I2(VCC_net), 
            .I3(n40788), .O(n1862[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_9 (.CI(n40788), .I0(n1803), .I1(VCC_net), 
            .CO(n40789));
    SB_LUT4 mod_5_add_1272_8_lut (.I0(GND_net), .I1(n1804), .I2(VCC_net), 
            .I3(n40787), .O(n1862[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_8 (.CI(n40787), .I0(n1804), .I1(VCC_net), 
            .CO(n40788));
    SB_LUT4 mod_5_add_1272_7_lut (.I0(GND_net), .I1(n1805), .I2(VCC_net), 
            .I3(n40786), .O(n1862[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_7 (.CI(n40786), .I0(n1805), .I1(VCC_net), 
            .CO(n40787));
    SB_LUT4 mod_5_add_1272_6_lut (.I0(GND_net), .I1(n1806), .I2(VCC_net), 
            .I3(n40785), .O(n1862[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_6 (.CI(n40785), .I0(n1806), .I1(VCC_net), 
            .CO(n40786));
    SB_LUT4 mod_5_add_1272_5_lut (.I0(GND_net), .I1(n1807), .I2(VCC_net), 
            .I3(n40784), .O(n1862[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_5 (.CI(n40784), .I0(n1807), .I1(VCC_net), 
            .CO(n40785));
    SB_LUT4 mod_5_add_1272_4_lut (.I0(GND_net), .I1(n1808), .I2(VCC_net), 
            .I3(n40783), .O(n1862[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_4 (.CI(n40783), .I0(n1808), .I1(VCC_net), 
            .CO(n40784));
    SB_LUT4 mod_5_add_1272_3_lut (.I0(GND_net), .I1(n1809), .I2(GND_net), 
            .I3(n40782), .O(n1862[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_3 (.CI(n40782), .I0(n1809), .I1(GND_net), 
            .CO(n40783));
    SB_LUT4 mod_5_add_1272_2_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(VCC_net), .O(n1862[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1272_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1272_2 (.CI(VCC_net), .I0(bit_ctr[17]), .I1(GND_net), 
            .CO(n40782));
    SB_LUT4 mod_5_add_1339_17_lut (.I0(n1928), .I1(n1895), .I2(VCC_net), 
            .I3(n40781), .O(n1994)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1339_16_lut (.I0(GND_net), .I1(n1896), .I2(VCC_net), 
            .I3(n40780), .O(n1961[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_16 (.CI(n40780), .I0(n1896), .I1(VCC_net), 
            .CO(n40781));
    SB_LUT4 mod_5_add_1339_15_lut (.I0(GND_net), .I1(n1897), .I2(VCC_net), 
            .I3(n40779), .O(n1961[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_15 (.CI(n40779), .I0(n1897), .I1(VCC_net), 
            .CO(n40780));
    SB_LUT4 mod_5_add_1339_14_lut (.I0(GND_net), .I1(n1898), .I2(VCC_net), 
            .I3(n40778), .O(n1961[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_14 (.CI(n40778), .I0(n1898), .I1(VCC_net), 
            .CO(n40779));
    SB_LUT4 mod_5_add_1339_13_lut (.I0(GND_net), .I1(n1899), .I2(VCC_net), 
            .I3(n40777), .O(n1961[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_13 (.CI(n40777), .I0(n1899), .I1(VCC_net), 
            .CO(n40778));
    SB_LUT4 mod_5_add_1339_12_lut (.I0(GND_net), .I1(n1900), .I2(VCC_net), 
            .I3(n40776), .O(n1961[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_12 (.CI(n40776), .I0(n1900), .I1(VCC_net), 
            .CO(n40777));
    SB_CARRY mod_5_add_1071_7 (.CI(n39419), .I0(n1505), .I1(VCC_net), 
            .CO(n39420));
    SB_CARRY timer_1546_add_4_3 (.CI(n40360), .I0(GND_net), .I1(timer[1]), 
            .CO(n40361));
    SB_LUT4 mod_5_add_1339_11_lut (.I0(GND_net), .I1(n1901), .I2(VCC_net), 
            .I3(n40775), .O(n1961[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_11 (.CI(n40775), .I0(n1901), .I1(VCC_net), 
            .CO(n40776));
    SB_LUT4 mod_5_add_1339_10_lut (.I0(GND_net), .I1(n1902), .I2(VCC_net), 
            .I3(n40774), .O(n1961[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_10 (.CI(n40774), .I0(n1902), .I1(VCC_net), 
            .CO(n40775));
    SB_LUT4 mod_5_add_1339_9_lut (.I0(GND_net), .I1(n1903), .I2(VCC_net), 
            .I3(n40773), .O(n1961[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i30_1_lut (.I0(\neo_pixel_transmitter.t0 [29]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[29]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i30_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY mod_5_add_1339_9 (.CI(n40773), .I0(n1903), .I1(VCC_net), 
            .CO(n40774));
    SB_LUT4 mod_5_add_1339_8_lut (.I0(GND_net), .I1(n1904), .I2(VCC_net), 
            .I3(n40772), .O(n1961[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_8 (.CI(n40772), .I0(n1904), .I1(VCC_net), 
            .CO(n40773));
    SB_LUT4 mod_5_add_1339_7_lut (.I0(GND_net), .I1(n1905), .I2(VCC_net), 
            .I3(n40771), .O(n1961[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_7 (.CI(n40771), .I0(n1905), .I1(VCC_net), 
            .CO(n40772));
    SB_LUT4 mod_5_add_1339_6_lut (.I0(GND_net), .I1(n1906), .I2(VCC_net), 
            .I3(n40770), .O(n1961[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_6 (.CI(n40770), .I0(n1906), .I1(VCC_net), 
            .CO(n40771));
    SB_LUT4 mod_5_add_1339_5_lut (.I0(GND_net), .I1(n1907), .I2(VCC_net), 
            .I3(n40769), .O(n1961[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_5 (.CI(n40769), .I0(n1907), .I1(VCC_net), 
            .CO(n40770));
    SB_LUT4 mod_5_add_1339_4_lut (.I0(GND_net), .I1(n1908), .I2(VCC_net), 
            .I3(n40768), .O(n1961[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_4 (.CI(n40768), .I0(n1908), .I1(VCC_net), 
            .CO(n40769));
    SB_LUT4 mod_5_add_1339_3_lut (.I0(GND_net), .I1(n1909), .I2(GND_net), 
            .I3(n40767), .O(n1961[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_3 (.CI(n40767), .I0(n1909), .I1(GND_net), 
            .CO(n40768));
    SB_LUT4 mod_5_add_1339_2_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(VCC_net), .O(n1961[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1339_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1339_2 (.CI(VCC_net), .I0(bit_ctr[16]), .I1(GND_net), 
            .CO(n40767));
    SB_LUT4 mod_5_add_1406_18_lut (.I0(n2027), .I1(n1994), .I2(VCC_net), 
            .I3(n40766), .O(n2093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_18_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1406_17_lut (.I0(GND_net), .I1(n1995), .I2(VCC_net), 
            .I3(n40765), .O(n2060[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_17 (.CI(n40765), .I0(n1995), .I1(VCC_net), 
            .CO(n40766));
    SB_LUT4 mod_5_add_1406_16_lut (.I0(GND_net), .I1(n1996), .I2(VCC_net), 
            .I3(n40764), .O(n2060[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_16 (.CI(n40764), .I0(n1996), .I1(VCC_net), 
            .CO(n40765));
    SB_LUT4 mod_5_add_1406_15_lut (.I0(GND_net), .I1(n1997), .I2(VCC_net), 
            .I3(n40763), .O(n2060[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_6_lut (.I0(GND_net), .I1(n1506), .I2(VCC_net), 
            .I3(n39418), .O(n1565[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_15 (.CI(n40763), .I0(n1997), .I1(VCC_net), 
            .CO(n40764));
    SB_LUT4 mod_5_add_1406_14_lut (.I0(GND_net), .I1(n1998), .I2(VCC_net), 
            .I3(n40762), .O(n2060[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_14 (.CI(n40762), .I0(n1998), .I1(VCC_net), 
            .CO(n40763));
    SB_LUT4 mod_5_add_1406_13_lut (.I0(GND_net), .I1(n1999), .I2(VCC_net), 
            .I3(n40761), .O(n2060[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_13 (.CI(n40761), .I0(n1999), .I1(VCC_net), 
            .CO(n40762));
    SB_LUT4 mod_5_add_1406_12_lut (.I0(GND_net), .I1(n2000), .I2(VCC_net), 
            .I3(n40760), .O(n2060[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_12 (.CI(n40760), .I0(n2000), .I1(VCC_net), 
            .CO(n40761));
    SB_LUT4 mod_5_add_1406_11_lut (.I0(GND_net), .I1(n2001), .I2(VCC_net), 
            .I3(n40759), .O(n2060[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_11 (.CI(n40759), .I0(n2001), .I1(VCC_net), 
            .CO(n40760));
    SB_LUT4 mod_5_add_1406_10_lut (.I0(GND_net), .I1(n2002), .I2(VCC_net), 
            .I3(n40758), .O(n2060[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_10 (.CI(n40758), .I0(n2002), .I1(VCC_net), 
            .CO(n40759));
    SB_LUT4 mod_5_add_1406_9_lut (.I0(GND_net), .I1(n2003), .I2(VCC_net), 
            .I3(n40757), .O(n2060[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_9 (.CI(n40757), .I0(n2003), .I1(VCC_net), 
            .CO(n40758));
    SB_LUT4 sub_14_inv_0_i31_1_lut (.I0(\neo_pixel_transmitter.t0 [30]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[30]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i31_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i36455_1_lut (.I0(n2621), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51408));
    defparam i36455_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 timer_1546_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(timer[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam timer_1546_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i32_1_lut (.I0(\neo_pixel_transmitter.t0 [31]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[31]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i32_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1406_8_lut (.I0(GND_net), .I1(n2004), .I2(VCC_net), 
            .I3(n40756), .O(n2060[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_8 (.CI(n40756), .I0(n2004), .I1(VCC_net), 
            .CO(n40757));
    SB_LUT4 mod_5_add_1406_7_lut (.I0(GND_net), .I1(n2005), .I2(VCC_net), 
            .I3(n40755), .O(n2060[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_7 (.CI(n40755), .I0(n2005), .I1(VCC_net), 
            .CO(n40756));
    SB_LUT4 mod_5_add_1406_6_lut (.I0(GND_net), .I1(n2006), .I2(VCC_net), 
            .I3(n40754), .O(n2060[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_6 (.CI(n40754), .I0(n2006), .I1(VCC_net), 
            .CO(n40755));
    SB_LUT4 mod_5_add_1406_5_lut (.I0(GND_net), .I1(n2007), .I2(VCC_net), 
            .I3(n40753), .O(n2060[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_5 (.CI(n40753), .I0(n2007), .I1(VCC_net), 
            .CO(n40754));
    SB_LUT4 mod_5_add_1406_4_lut (.I0(GND_net), .I1(n2008), .I2(VCC_net), 
            .I3(n40752), .O(n2060[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_4 (.CI(n40752), .I0(n2008), .I1(VCC_net), 
            .CO(n40753));
    SB_LUT4 mod_5_add_1406_3_lut (.I0(GND_net), .I1(n2009), .I2(GND_net), 
            .I3(n40751), .O(n2060[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_3 (.CI(n40751), .I0(n2009), .I1(GND_net), 
            .CO(n40752));
    SB_CARRY timer_1546_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(timer[0]), 
            .CO(n40360));
    SB_LUT4 mod_5_add_1406_2_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(VCC_net), .O(n2060[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1406_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1406_2 (.CI(VCC_net), .I0(bit_ctr[15]), .I1(GND_net), 
            .CO(n40751));
    SB_LUT4 mod_5_add_1473_19_lut (.I0(n2126), .I1(n2093), .I2(VCC_net), 
            .I3(n40750), .O(n2192)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_19_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_870_10_lut (.I0(n1202), .I1(n1202), .I2(n1235), 
            .I3(n40359), .O(n1301)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1071_6 (.CI(n39418), .I0(n1506), .I1(VCC_net), 
            .CO(n39419));
    SB_LUT4 mod_5_add_1071_5_lut (.I0(GND_net), .I1(n1507), .I2(VCC_net), 
            .I3(n39417), .O(n1565[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_870_9_lut (.I0(n1203), .I1(n1203), .I2(n1235), .I3(n40358), 
            .O(n1302)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_9 (.CI(n40358), .I0(n1203), .I1(n1235), .CO(n40359));
    SB_CARRY mod_5_add_1071_5 (.CI(n39417), .I0(n1507), .I1(VCC_net), 
            .CO(n39418));
    SB_LUT4 mod_5_add_870_8_lut (.I0(n1204), .I1(n1204), .I2(n1235), .I3(n40357), 
            .O(n1303)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_8_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_18_lut (.I0(GND_net), .I1(n2094), .I2(VCC_net), 
            .I3(n40749), .O(n2159[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_870_8 (.CI(n40357), .I0(n1204), .I1(n1235), .CO(n40358));
    SB_CARRY mod_5_add_1473_18 (.CI(n40749), .I0(n2094), .I1(VCC_net), 
            .CO(n40750));
    SB_LUT4 mod_5_add_870_7_lut (.I0(n1205), .I1(n1205), .I2(n1235), .I3(n40356), 
            .O(n1304)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_7 (.CI(n40356), .I0(n1205), .I1(n1235), .CO(n40357));
    SB_LUT4 mod_5_add_1473_17_lut (.I0(GND_net), .I1(n2095), .I2(VCC_net), 
            .I3(n40748), .O(n2159[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_17 (.CI(n40748), .I0(n2095), .I1(VCC_net), 
            .CO(n40749));
    SB_LUT4 mod_5_add_1473_16_lut (.I0(GND_net), .I1(n2096), .I2(VCC_net), 
            .I3(n40747), .O(n2159[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_16 (.CI(n40747), .I0(n2096), .I1(VCC_net), 
            .CO(n40748));
    SB_LUT4 mod_5_add_1473_15_lut (.I0(GND_net), .I1(n2097), .I2(VCC_net), 
            .I3(n40746), .O(n2159[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_15 (.CI(n40746), .I0(n2097), .I1(VCC_net), 
            .CO(n40747));
    SB_LUT4 mod_5_add_870_6_lut (.I0(n1206), .I1(n1206), .I2(n1235), .I3(n40355), 
            .O(n1305)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1473_14_lut (.I0(GND_net), .I1(n2098), .I2(VCC_net), 
            .I3(n40745), .O(n2159[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_14 (.CI(n40745), .I0(n2098), .I1(VCC_net), 
            .CO(n40746));
    SB_LUT4 mod_5_add_1473_13_lut (.I0(GND_net), .I1(n2099), .I2(VCC_net), 
            .I3(n40744), .O(n2159[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF timer_1546__i0 (.Q(timer[0]), .C(CLK_c), .D(n133[0]));   // verilog/neopixel.v(12[12:21])
    SB_CARRY mod_5_add_1473_13 (.CI(n40744), .I0(n2099), .I1(VCC_net), 
            .CO(n40745));
    SB_LUT4 mod_5_add_1473_12_lut (.I0(GND_net), .I1(n2100), .I2(VCC_net), 
            .I3(n40743), .O(n2159[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1897_3_lut (.I0(n2707), .I1(n2753[11]), .I2(n2720), 
            .I3(GND_net), .O(n2806));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1897_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1895_3_lut (.I0(n2705), .I1(n2753[13]), .I2(n2720), 
            .I3(GND_net), .O(n2804));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1895_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1889_3_lut (.I0(n2699), .I1(n2753[19]), .I2(n2720), 
            .I3(GND_net), .O(n2798));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1889_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1896_3_lut (.I0(n2706), .I1(n2753[12]), .I2(n2720), 
            .I3(GND_net), .O(n2805));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1896_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1878_3_lut (.I0(n2688), .I1(n2753[30]), .I2(n2720), 
            .I3(GND_net), .O(n2787));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1878_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1887_3_lut (.I0(n2697), .I1(n2753[21]), .I2(n2720), 
            .I3(GND_net), .O(n2796));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1887_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1886_3_lut (.I0(n2696), .I1(n2753[22]), .I2(n2720), 
            .I3(GND_net), .O(n2795));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1886_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_870_6 (.CI(n40355), .I0(n1206), .I1(n1235), .CO(n40356));
    SB_LUT4 mod_5_add_870_5_lut (.I0(n1207), .I1(n1207), .I2(n1235), .I3(n40354), 
            .O(n1306)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_870_5 (.CI(n40354), .I0(n1207), .I1(n1235), .CO(n40355));
    SB_CARRY mod_5_add_1473_12 (.CI(n40743), .I0(n2100), .I1(VCC_net), 
            .CO(n40744));
    SB_LUT4 mod_5_i1892_3_lut (.I0(n2702), .I1(n2753[16]), .I2(n2720), 
            .I3(GND_net), .O(n2801));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1892_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1473_11_lut (.I0(GND_net), .I1(n2101), .I2(VCC_net), 
            .I3(n40742), .O(n2159[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_4_lut (.I0(GND_net), .I1(n1508), .I2(VCC_net), 
            .I3(n39416), .O(n1565[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_11 (.CI(n40742), .I0(n2101), .I1(VCC_net), 
            .CO(n40743));
    SB_CARRY mod_5_add_1071_4 (.CI(n39416), .I0(n1508), .I1(VCC_net), 
            .CO(n39417));
    SB_LUT4 mod_5_add_1473_10_lut (.I0(GND_net), .I1(n2102), .I2(VCC_net), 
            .I3(n40741), .O(n2159[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_10 (.CI(n40741), .I0(n2102), .I1(VCC_net), 
            .CO(n40742));
    SB_LUT4 mod_5_i1888_3_lut (.I0(n2698), .I1(n2753[20]), .I2(n2720), 
            .I3(GND_net), .O(n2797));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1888_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1473_9_lut (.I0(GND_net), .I1(n2103), .I2(VCC_net), 
            .I3(n40740), .O(n2159[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1891_3_lut (.I0(n2701), .I1(n2753[17]), .I2(n2720), 
            .I3(GND_net), .O(n2800));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1891_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1473_9 (.CI(n40740), .I0(n2103), .I1(VCC_net), 
            .CO(n40741));
    SB_LUT4 mod_5_i1884_3_lut (.I0(n2694), .I1(n2753[24]), .I2(n2720), 
            .I3(GND_net), .O(n2793));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1884_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1473_8_lut (.I0(GND_net), .I1(n2104), .I2(VCC_net), 
            .I3(n40739), .O(n2159[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1890_3_lut (.I0(n2700), .I1(n2753[18]), .I2(n2720), 
            .I3(GND_net), .O(n2799));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1890_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1473_8 (.CI(n40739), .I0(n2104), .I1(VCC_net), 
            .CO(n40740));
    SB_LUT4 mod_5_i1882_3_lut (.I0(n2692), .I1(n2753[26]), .I2(n2720), 
            .I3(GND_net), .O(n2791));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1882_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1473_7_lut (.I0(GND_net), .I1(n2105), .I2(VCC_net), 
            .I3(n40738), .O(n2159[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1883_3_lut (.I0(n2693), .I1(n2753[25]), .I2(n2720), 
            .I3(GND_net), .O(n2792));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1883_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1473_7 (.CI(n40738), .I0(n2105), .I1(VCC_net), 
            .CO(n40739));
    SB_LUT4 mod_5_i1881_3_lut (.I0(n2691), .I1(n2753[27]), .I2(n2720), 
            .I3(GND_net), .O(n2790));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1881_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1473_6_lut (.I0(GND_net), .I1(n2106), .I2(VCC_net), 
            .I3(n40737), .O(n2159[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1880_3_lut (.I0(n2690), .I1(n2753[28]), .I2(n2720), 
            .I3(GND_net), .O(n2789));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1880_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1473_6 (.CI(n40737), .I0(n2106), .I1(VCC_net), 
            .CO(n40738));
    SB_LUT4 mod_5_i1899_3_lut (.I0(n2709), .I1(n2753[9]), .I2(n2720), 
            .I3(GND_net), .O(n2808));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1899_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1473_5_lut (.I0(GND_net), .I1(n2107), .I2(VCC_net), 
            .I3(n40736), .O(n2159[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1885_3_lut (.I0(n2695), .I1(n2753[23]), .I2(n2720), 
            .I3(GND_net), .O(n2794));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1885_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1473_5 (.CI(n40736), .I0(n2107), .I1(VCC_net), 
            .CO(n40737));
    SB_LUT4 mod_5_add_1473_4_lut (.I0(GND_net), .I1(n2108), .I2(VCC_net), 
            .I3(n40735), .O(n2159[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1893_3_lut (.I0(n2703), .I1(n2753[15]), .I2(n2720), 
            .I3(GND_net), .O(n2802));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1893_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1473_4 (.CI(n40735), .I0(n2108), .I1(VCC_net), 
            .CO(n40736));
    SB_LUT4 mod_5_i1898_3_lut (.I0(n2708), .I1(n2753[10]), .I2(n2720), 
            .I3(GND_net), .O(n2807));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1898_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1473_3_lut (.I0(GND_net), .I1(n2109), .I2(GND_net), 
            .I3(n40734), .O(n2159[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1473_3 (.CI(n40734), .I0(n2109), .I1(GND_net), 
            .CO(n40735));
    SB_LUT4 i7_3_lut (.I0(bit_ctr[8]), .I1(n2705), .I2(n2709), .I3(GND_net), 
            .O(n30_adj_4812));   // verilog/neopixel.v(22[26:36])
    defparam i7_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_1473_2_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(VCC_net), .O(n2159[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1473_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14_4_lut_adj_1585 (.I0(n2694), .I1(n2697), .I2(n2693), .I3(n2695), 
            .O(n37));   // verilog/neopixel.v(22[26:36])
    defparam i14_4_lut_adj_1585.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1473_2 (.CI(VCC_net), .I0(bit_ctr[14]), .I1(GND_net), 
            .CO(n40734));
    SB_LUT4 mod_5_add_1540_20_lut (.I0(n2225), .I1(n2192), .I2(VCC_net), 
            .I3(n40733), .O(n2291)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_20_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i13_4_lut_adj_1586 (.I0(n2689), .I1(n2691), .I2(n2692), .I3(n2690), 
            .O(n36));   // verilog/neopixel.v(22[26:36])
    defparam i13_4_lut_adj_1586.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_19_lut (.I0(GND_net), .I1(n2193), .I2(VCC_net), 
            .I3(n40732), .O(n2258[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i19_4_lut_adj_1587 (.I0(n37), .I1(n2698), .I2(n30_adj_4812), 
            .I3(n2696), .O(n42));   // verilog/neopixel.v(22[26:36])
    defparam i19_4_lut_adj_1587.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1540_19 (.CI(n40732), .I0(n2193), .I1(VCC_net), 
            .CO(n40733));
    SB_LUT4 i17_4_lut_adj_1588 (.I0(n2700), .I1(n2702), .I2(n2703), .I3(n2704), 
            .O(n40));   // verilog/neopixel.v(22[26:36])
    defparam i17_4_lut_adj_1588.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_18_lut (.I0(GND_net), .I1(n2194), .I2(VCC_net), 
            .I3(n40731), .O(n2258[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18_4_lut_adj_1589 (.I0(n2706), .I1(n36), .I2(n2688), .I3(n2687), 
            .O(n41));   // verilog/neopixel.v(22[26:36])
    defparam i18_4_lut_adj_1589.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1540_18 (.CI(n40731), .I0(n2194), .I1(VCC_net), 
            .CO(n40732));
    SB_LUT4 i16_4_lut_adj_1590 (.I0(n2701), .I1(n2699), .I2(n2707), .I3(n2708), 
            .O(n39_adj_4813));   // verilog/neopixel.v(22[26:36])
    defparam i16_4_lut_adj_1590.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_17_lut (.I0(GND_net), .I1(n2195), .I2(VCC_net), 
            .I3(n40730), .O(n2258[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i22_4_lut (.I0(n39_adj_4813), .I1(n41), .I2(n40), .I3(n42), 
            .O(n2720));   // verilog/neopixel.v(22[26:36])
    defparam i22_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1540_17 (.CI(n40730), .I0(n2195), .I1(VCC_net), 
            .CO(n40731));
    SB_LUT4 mod_5_i1900_3_lut (.I0(bit_ctr[8]), .I1(n2753[8]), .I2(n2720), 
            .I3(GND_net), .O(n2809));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1900_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1540_16_lut (.I0(GND_net), .I1(n2196), .I2(VCC_net), 
            .I3(n40729), .O(n2258[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1894_3_lut (.I0(n2704), .I1(n2753[14]), .I2(n2720), 
            .I3(GND_net), .O(n2803));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1894_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1540_16 (.CI(n40729), .I0(n2196), .I1(VCC_net), 
            .CO(n40730));
    SB_LUT4 i6_3_lut_adj_1591 (.I0(bit_ctr[7]), .I1(n2803), .I2(n2809), 
            .I3(GND_net), .O(n30_adj_4814));   // verilog/neopixel.v(22[26:36])
    defparam i6_3_lut_adj_1591.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_add_1540_15_lut (.I0(GND_net), .I1(n2197), .I2(VCC_net), 
            .I3(n40728), .O(n2258[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i16_4_lut_adj_1592 (.I0(n2807), .I1(n2802), .I2(n2794), .I3(n2808), 
            .O(n40_adj_4815));   // verilog/neopixel.v(22[26:36])
    defparam i16_4_lut_adj_1592.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1540_15 (.CI(n40728), .I0(n2197), .I1(VCC_net), 
            .CO(n40729));
    SB_LUT4 i2_2_lut (.I0(n2788), .I1(n2789), .I2(GND_net), .I3(GND_net), 
            .O(n26_adj_4816));   // verilog/neopixel.v(22[26:36])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_1540_14_lut (.I0(GND_net), .I1(n2198), .I2(VCC_net), 
            .I3(n40727), .O(n2258[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i14_4_lut_adj_1593 (.I0(n2790), .I1(n2792), .I2(n2791), .I3(n2799), 
            .O(n38));   // verilog/neopixel.v(22[26:36])
    defparam i14_4_lut_adj_1593.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1540_14 (.CI(n40727), .I0(n2198), .I1(VCC_net), 
            .CO(n40728));
    SB_LUT4 i20_4_lut_adj_1594 (.I0(n2793), .I1(n40_adj_4815), .I2(n30_adj_4814), 
            .I3(n2800), .O(n44_adj_4817));   // verilog/neopixel.v(22[26:36])
    defparam i20_4_lut_adj_1594.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1540_13_lut (.I0(GND_net), .I1(n2199), .I2(VCC_net), 
            .I3(n40726), .O(n2258[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i18_4_lut_adj_1595 (.I0(n2797), .I1(n2801), .I2(n2795), .I3(n2796), 
            .O(n42_adj_4818));   // verilog/neopixel.v(22[26:36])
    defparam i18_4_lut_adj_1595.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1540_13 (.CI(n40726), .I0(n2199), .I1(VCC_net), 
            .CO(n40727));
    SB_LUT4 mod_5_add_1540_12_lut (.I0(GND_net), .I1(n2200), .I2(VCC_net), 
            .I3(n40725), .O(n2258[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_12 (.CI(n40725), .I0(n2200), .I1(VCC_net), 
            .CO(n40726));
    SB_LUT4 mod_5_add_1540_11_lut (.I0(GND_net), .I1(n2201), .I2(VCC_net), 
            .I3(n40724), .O(n2258[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_11 (.CI(n40724), .I0(n2201), .I1(VCC_net), 
            .CO(n40725));
    SB_LUT4 mod_5_add_870_4_lut (.I0(n1208), .I1(n1208), .I2(n1235), .I3(n40353), 
            .O(n1307)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_4_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1540_10_lut (.I0(GND_net), .I1(n2202), .I2(VCC_net), 
            .I3(n40723), .O(n2258[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_10 (.CI(n40723), .I0(n2202), .I1(VCC_net), 
            .CO(n40724));
    SB_LUT4 mod_5_add_1540_9_lut (.I0(GND_net), .I1(n2203), .I2(VCC_net), 
            .I3(n40722), .O(n2258[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_9 (.CI(n40722), .I0(n2203), .I1(VCC_net), 
            .CO(n40723));
    SB_LUT4 mod_5_add_1540_8_lut (.I0(GND_net), .I1(n2204), .I2(VCC_net), 
            .I3(n40721), .O(n2258[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1071_3_lut (.I0(GND_net), .I1(n1509), .I2(GND_net), 
            .I3(n39415), .O(n1565[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_8 (.CI(n40721), .I0(n2204), .I1(VCC_net), 
            .CO(n40722));
    SB_LUT4 mod_5_add_1540_7_lut (.I0(GND_net), .I1(n2205), .I2(VCC_net), 
            .I3(n40720), .O(n2258[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_7 (.CI(n40720), .I0(n2205), .I1(VCC_net), 
            .CO(n40721));
    SB_LUT4 mod_5_add_1540_6_lut (.I0(GND_net), .I1(n2206), .I2(VCC_net), 
            .I3(n40719), .O(n2258[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_6 (.CI(n40719), .I0(n2206), .I1(VCC_net), 
            .CO(n40720));
    SB_LUT4 mod_5_add_1540_5_lut (.I0(GND_net), .I1(n2207), .I2(VCC_net), 
            .I3(n40718), .O(n2258[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_3 (.CI(n39415), .I0(n1509), .I1(GND_net), 
            .CO(n39416));
    SB_CARRY mod_5_add_1540_5 (.CI(n40718), .I0(n2207), .I1(VCC_net), 
            .CO(n40719));
    SB_LUT4 mod_5_add_1540_4_lut (.I0(GND_net), .I1(n2208), .I2(VCC_net), 
            .I3(n40717), .O(n2258[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_4 (.CI(n40717), .I0(n2208), .I1(VCC_net), 
            .CO(n40718));
    SB_CARRY mod_5_add_870_4 (.CI(n40353), .I0(n1208), .I1(n1235), .CO(n40354));
    SB_LUT4 mod_5_add_1071_2_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(VCC_net), .O(n1565[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1071_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1071_2 (.CI(VCC_net), .I0(bit_ctr[20]), .I1(GND_net), 
            .CO(n39415));
    SB_LUT4 mod_5_add_870_3_lut (.I0(n1209), .I1(n1209), .I2(n51406), 
            .I3(n40352), .O(n1308)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 mod_5_add_1540_3_lut (.I0(GND_net), .I1(n2209), .I2(GND_net), 
            .I3(n40716), .O(n2258[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_3 (.CI(n40716), .I0(n2209), .I1(GND_net), 
            .CO(n40717));
    SB_LUT4 mod_5_add_1540_2_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(VCC_net), .O(n2258[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1540_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1540_2 (.CI(VCC_net), .I0(bit_ctr[13]), .I1(GND_net), 
            .CO(n40716));
    SB_LUT4 mod_5_add_1607_21_lut (.I0(n2324), .I1(n2291), .I2(VCC_net), 
            .I3(n40715), .O(n2390)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_21_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1607_20_lut (.I0(GND_net), .I1(n2292), .I2(VCC_net), 
            .I3(n40714), .O(n2357[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_20 (.CI(n40714), .I0(n2292), .I1(VCC_net), 
            .CO(n40715));
    SB_LUT4 mod_5_add_1607_19_lut (.I0(GND_net), .I1(n2293), .I2(VCC_net), 
            .I3(n40713), .O(n2357[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_870_3 (.CI(n40352), .I0(n1209), .I1(n51406), .CO(n40353));
    SB_LUT4 mod_5_add_870_2_lut (.I0(bit_ctr[23]), .I1(bit_ctr[23]), .I2(n51406), 
            .I3(VCC_net), .O(n1309)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_870_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1607_19 (.CI(n40713), .I0(n2293), .I1(VCC_net), 
            .CO(n40714));
    SB_LUT4 mod_5_add_1607_18_lut (.I0(GND_net), .I1(n2294), .I2(VCC_net), 
            .I3(n40712), .O(n2357[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_870_2 (.CI(VCC_net), .I0(bit_ctr[23]), .I1(n51406), 
            .CO(n40352));
    SB_LUT4 mod_5_add_2076_28_lut (.I0(n2984), .I1(n2984), .I2(n3017), 
            .I3(n40351), .O(n3083)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_28_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_2076_27_lut (.I0(n2985), .I1(n2985), .I2(n3017), 
            .I3(n40350), .O(n3084)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_27_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1607_18 (.CI(n40712), .I0(n2294), .I1(VCC_net), 
            .CO(n40713));
    SB_LUT4 mod_5_add_1607_17_lut (.I0(GND_net), .I1(n2295), .I2(VCC_net), 
            .I3(n40711), .O(n2357[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_17 (.CI(n40711), .I0(n2295), .I1(VCC_net), 
            .CO(n40712));
    SB_LUT4 mod_5_add_1607_16_lut (.I0(GND_net), .I1(n2296), .I2(VCC_net), 
            .I3(n40710), .O(n2357[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_16 (.CI(n40710), .I0(n2296), .I1(VCC_net), 
            .CO(n40711));
    SB_CARRY mod_5_add_2076_27 (.CI(n40350), .I0(n2985), .I1(n3017), .CO(n40351));
    SB_LUT4 mod_5_add_2076_26_lut (.I0(n2986), .I1(n2986), .I2(n3017), 
            .I3(n40349), .O(n3085)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_26_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1607_15_lut (.I0(GND_net), .I1(n2297), .I2(VCC_net), 
            .I3(n40709), .O(n2357[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_15 (.CI(n40709), .I0(n2297), .I1(VCC_net), 
            .CO(n40710));
    SB_LUT4 mod_5_add_1607_14_lut (.I0(GND_net), .I1(n2298), .I2(VCC_net), 
            .I3(n40708), .O(n2357[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_14 (.CI(n40708), .I0(n2298), .I1(VCC_net), 
            .CO(n40709));
    SB_LUT4 mod_5_add_1607_13_lut (.I0(GND_net), .I1(n2299), .I2(VCC_net), 
            .I3(n40707), .O(n2357[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_13 (.CI(n40707), .I0(n2299), .I1(VCC_net), 
            .CO(n40708));
    SB_LUT4 mod_5_add_1607_12_lut (.I0(GND_net), .I1(n2300), .I2(VCC_net), 
            .I3(n40706), .O(n2357[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_12 (.CI(n40706), .I0(n2300), .I1(VCC_net), 
            .CO(n40707));
    SB_LUT4 mod_5_add_1607_11_lut (.I0(GND_net), .I1(n2301), .I2(VCC_net), 
            .I3(n40705), .O(n2357[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_11 (.CI(n40705), .I0(n2301), .I1(VCC_net), 
            .CO(n40706));
    SB_LUT4 mod_5_add_1607_10_lut (.I0(GND_net), .I1(n2302), .I2(VCC_net), 
            .I3(n40704), .O(n2357[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_10 (.CI(n40704), .I0(n2302), .I1(VCC_net), 
            .CO(n40705));
    SB_LUT4 mod_5_add_1607_9_lut (.I0(GND_net), .I1(n2303), .I2(VCC_net), 
            .I3(n40703), .O(n2357[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_9 (.CI(n40703), .I0(n2303), .I1(VCC_net), 
            .CO(n40704));
    SB_LUT4 mod_5_add_1607_8_lut (.I0(GND_net), .I1(n2304), .I2(VCC_net), 
            .I3(n40702), .O(n2357[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_8 (.CI(n40702), .I0(n2304), .I1(VCC_net), 
            .CO(n40703));
    SB_LUT4 mod_5_add_1607_7_lut (.I0(GND_net), .I1(n2305), .I2(VCC_net), 
            .I3(n40701), .O(n2357[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_7 (.CI(n40701), .I0(n2305), .I1(VCC_net), 
            .CO(n40702));
    SB_LUT4 mod_5_add_1607_6_lut (.I0(GND_net), .I1(n2306), .I2(VCC_net), 
            .I3(n40700), .O(n2357[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_6 (.CI(n40700), .I0(n2306), .I1(VCC_net), 
            .CO(n40701));
    SB_LUT4 mod_5_add_1607_5_lut (.I0(GND_net), .I1(n2307), .I2(VCC_net), 
            .I3(n40699), .O(n2357[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_5 (.CI(n40699), .I0(n2307), .I1(VCC_net), 
            .CO(n40700));
    SB_LUT4 mod_5_add_1607_4_lut (.I0(GND_net), .I1(n2308), .I2(VCC_net), 
            .I3(n40698), .O(n2357[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_4 (.CI(n40698), .I0(n2308), .I1(VCC_net), 
            .CO(n40699));
    SB_LUT4 mod_5_add_1607_3_lut (.I0(GND_net), .I1(n2309), .I2(GND_net), 
            .I3(n40697), .O(n2357[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_3 (.CI(n40697), .I0(n2309), .I1(GND_net), 
            .CO(n40698));
    SB_LUT4 mod_5_add_1607_2_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(VCC_net), .O(n2357[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1607_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1607_2 (.CI(VCC_net), .I0(bit_ctr[12]), .I1(GND_net), 
            .CO(n40697));
    SB_LUT4 mod_5_add_1674_22_lut (.I0(n2423), .I1(n2390), .I2(VCC_net), 
            .I3(n40696), .O(n2489)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_22_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1674_21_lut (.I0(GND_net), .I1(n2391), .I2(VCC_net), 
            .I3(n40695), .O(n2456[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_21 (.CI(n40695), .I0(n2391), .I1(VCC_net), 
            .CO(n40696));
    SB_LUT4 mod_5_add_1674_20_lut (.I0(GND_net), .I1(n2392), .I2(VCC_net), 
            .I3(n40694), .O(n2456[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_20 (.CI(n40694), .I0(n2392), .I1(VCC_net), 
            .CO(n40695));
    SB_LUT4 mod_5_add_1674_19_lut (.I0(GND_net), .I1(n2393), .I2(VCC_net), 
            .I3(n40693), .O(n2456[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_19 (.CI(n40693), .I0(n2393), .I1(VCC_net), 
            .CO(n40694));
    SB_LUT4 mod_5_add_1674_18_lut (.I0(GND_net), .I1(n2394), .I2(VCC_net), 
            .I3(n40692), .O(n2456[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_18 (.CI(n40692), .I0(n2394), .I1(VCC_net), 
            .CO(n40693));
    SB_LUT4 mod_5_add_1674_17_lut (.I0(GND_net), .I1(n2395), .I2(VCC_net), 
            .I3(n40691), .O(n2456[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_17 (.CI(n40691), .I0(n2395), .I1(VCC_net), 
            .CO(n40692));
    SB_LUT4 mod_5_add_1674_16_lut (.I0(GND_net), .I1(n2396), .I2(VCC_net), 
            .I3(n40690), .O(n2456[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_16 (.CI(n40690), .I0(n2396), .I1(VCC_net), 
            .CO(n40691));
    SB_CARRY mod_5_add_2076_26 (.CI(n40349), .I0(n2986), .I1(n3017), .CO(n40350));
    SB_LUT4 mod_5_add_1674_15_lut (.I0(GND_net), .I1(n2397), .I2(VCC_net), 
            .I3(n40689), .O(n2456[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2076_25_lut (.I0(n2987), .I1(n2987), .I2(n3017), 
            .I3(n40348), .O(n3086)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_25_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_15 (.CI(n40689), .I0(n2397), .I1(VCC_net), 
            .CO(n40690));
    SB_LUT4 i19_4_lut_adj_1596 (.I0(n2787), .I1(n38), .I2(n26_adj_4816), 
            .I3(n2786), .O(n43_adj_4819));   // verilog/neopixel.v(22[26:36])
    defparam i19_4_lut_adj_1596.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1674_14_lut (.I0(GND_net), .I1(n2398), .I2(VCC_net), 
            .I3(n40688), .O(n2456[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i17_4_lut_adj_1597 (.I0(n2805), .I1(n2798), .I2(n2804), .I3(n2806), 
            .O(n41_adj_4820));   // verilog/neopixel.v(22[26:36])
    defparam i17_4_lut_adj_1597.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1674_14 (.CI(n40688), .I0(n2398), .I1(VCC_net), 
            .CO(n40689));
    SB_LUT4 mod_5_add_1674_13_lut (.I0(GND_net), .I1(n2399), .I2(VCC_net), 
            .I3(n40687), .O(n2456[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_13 (.CI(n40687), .I0(n2399), .I1(VCC_net), 
            .CO(n40688));
    SB_LUT4 mod_5_add_1674_12_lut (.I0(GND_net), .I1(n2400), .I2(VCC_net), 
            .I3(n40686), .O(n2456[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_12 (.CI(n40686), .I0(n2400), .I1(VCC_net), 
            .CO(n40687));
    SB_LUT4 mod_5_add_1674_11_lut (.I0(GND_net), .I1(n2401), .I2(VCC_net), 
            .I3(n40685), .O(n2456[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_11 (.CI(n40685), .I0(n2401), .I1(VCC_net), 
            .CO(n40686));
    SB_LUT4 mod_5_add_1674_10_lut (.I0(GND_net), .I1(n2402), .I2(VCC_net), 
            .I3(n40684), .O(n2456[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_10 (.CI(n40684), .I0(n2402), .I1(VCC_net), 
            .CO(n40685));
    SB_LUT4 mod_5_add_1674_9_lut (.I0(GND_net), .I1(n2403), .I2(VCC_net), 
            .I3(n40683), .O(n2456[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_9 (.CI(n40683), .I0(n2403), .I1(VCC_net), 
            .CO(n40684));
    SB_CARRY mod_5_add_2076_25 (.CI(n40348), .I0(n2987), .I1(n3017), .CO(n40349));
    SB_LUT4 mod_5_add_1674_8_lut (.I0(GND_net), .I1(n2404), .I2(VCC_net), 
            .I3(n40682), .O(n2456[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_8 (.CI(n40682), .I0(n2404), .I1(VCC_net), 
            .CO(n40683));
    SB_LUT4 mod_5_add_1674_7_lut (.I0(GND_net), .I1(n2405), .I2(VCC_net), 
            .I3(n40681), .O(n2456[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1674_7 (.CI(n40681), .I0(n2405), .I1(VCC_net), 
            .CO(n40682));
    SB_LUT4 mod_5_add_2076_24_lut (.I0(n2988), .I1(n2988), .I2(n3017), 
            .I3(n40347), .O(n3087)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1674_6_lut (.I0(GND_net), .I1(n2406), .I2(VCC_net), 
            .I3(n40680), .O(n2456[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_24 (.CI(n40347), .I0(n2988), .I1(n3017), .CO(n40348));
    SB_LUT4 mod_5_add_2076_23_lut (.I0(n2989), .I1(n2989), .I2(n3017), 
            .I3(n40346), .O(n3088)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_23 (.CI(n40346), .I0(n2989), .I1(n3017), .CO(n40347));
    SB_LUT4 mod_5_add_2076_22_lut (.I0(n2990), .I1(n2990), .I2(n3017), 
            .I3(n40345), .O(n3089)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_22 (.CI(n40345), .I0(n2990), .I1(n3017), .CO(n40346));
    SB_CARRY mod_5_add_1674_6 (.CI(n40680), .I0(n2406), .I1(VCC_net), 
            .CO(n40681));
    SB_LUT4 mod_5_add_1674_5_lut (.I0(GND_net), .I1(n2407), .I2(VCC_net), 
            .I3(n40679), .O(n2456[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2076_21_lut (.I0(n2991), .I1(n2991), .I2(n3017), 
            .I3(n40344), .O(n3090)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_21_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_21 (.CI(n40344), .I0(n2991), .I1(n3017), .CO(n40345));
    SB_LUT4 mod_5_add_2076_20_lut (.I0(n2992), .I1(n2992), .I2(n3017), 
            .I3(n40343), .O(n3091)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_20_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_20 (.CI(n40343), .I0(n2992), .I1(n3017), .CO(n40344));
    SB_LUT4 mod_5_add_2076_19_lut (.I0(n2993), .I1(n2993), .I2(n3017), 
            .I3(n40342), .O(n3092)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_19 (.CI(n40342), .I0(n2993), .I1(n3017), .CO(n40343));
    SB_LUT4 mod_5_add_2076_18_lut (.I0(n2994), .I1(n2994), .I2(n3017), 
            .I3(n40341), .O(n3093)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_18 (.CI(n40341), .I0(n2994), .I1(n3017), .CO(n40342));
    SB_CARRY mod_5_add_1674_5 (.CI(n40679), .I0(n2407), .I1(VCC_net), 
            .CO(n40680));
    SB_LUT4 mod_5_add_2076_17_lut (.I0(n2995), .I1(n2995), .I2(n3017), 
            .I3(n40340), .O(n3094)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_17 (.CI(n40340), .I0(n2995), .I1(n3017), .CO(n40341));
    SB_LUT4 mod_5_add_2076_16_lut (.I0(n2996), .I1(n2996), .I2(n3017), 
            .I3(n40339), .O(n3095)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_16 (.CI(n40339), .I0(n2996), .I1(n3017), .CO(n40340));
    SB_LUT4 mod_5_add_2076_15_lut (.I0(n2997), .I1(n2997), .I2(n3017), 
            .I3(n40338), .O(n3096)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_15 (.CI(n40338), .I0(n2997), .I1(n3017), .CO(n40339));
    SB_LUT4 mod_5_add_1674_4_lut (.I0(GND_net), .I1(n2408), .I2(VCC_net), 
            .I3(n40678), .O(n2456[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2076_14_lut (.I0(n2998), .I1(n2998), .I2(n3017), 
            .I3(n40337), .O(n3097)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_14 (.CI(n40337), .I0(n2998), .I1(n3017), .CO(n40338));
    SB_LUT4 mod_5_add_2076_13_lut (.I0(n2999), .I1(n2999), .I2(n3017), 
            .I3(n40336), .O(n3098)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_13 (.CI(n40336), .I0(n2999), .I1(n3017), .CO(n40337));
    SB_LUT4 mod_5_add_2076_12_lut (.I0(n3000), .I1(n3000), .I2(n3017), 
            .I3(n40335), .O(n3099)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_12 (.CI(n40335), .I0(n3000), .I1(n3017), .CO(n40336));
    SB_LUT4 mod_5_add_2076_11_lut (.I0(n3001), .I1(n3001), .I2(n3017), 
            .I3(n40334), .O(n3100)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_11 (.CI(n40334), .I0(n3001), .I1(n3017), .CO(n40335));
    SB_LUT4 mod_5_add_2076_10_lut (.I0(n3002), .I1(n3002), .I2(n3017), 
            .I3(n40333), .O(n3101)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_10 (.CI(n40333), .I0(n3002), .I1(n3017), .CO(n40334));
    SB_LUT4 mod_5_add_2076_9_lut (.I0(n3003), .I1(n3003), .I2(n3017), 
            .I3(n40332), .O(n3102)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_9 (.CI(n40332), .I0(n3003), .I1(n3017), .CO(n40333));
    SB_LUT4 mod_5_add_2076_8_lut (.I0(n3004), .I1(n3004), .I2(n3017), 
            .I3(n40331), .O(n3103)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_8 (.CI(n40331), .I0(n3004), .I1(n3017), .CO(n40332));
    SB_LUT4 mod_5_add_2076_7_lut (.I0(n3005), .I1(n3005), .I2(n3017), 
            .I3(n40330), .O(n3104)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1674_4 (.CI(n40678), .I0(n2408), .I1(VCC_net), 
            .CO(n40679));
    SB_LUT4 mod_5_add_1674_3_lut (.I0(GND_net), .I1(n2409), .I2(GND_net), 
            .I3(n40677), .O(n2456[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2076_7 (.CI(n40330), .I0(n3005), .I1(n3017), .CO(n40331));
    SB_CARRY mod_5_add_1674_3 (.CI(n40677), .I0(n2409), .I1(GND_net), 
            .CO(n40678));
    SB_LUT4 mod_5_add_2076_6_lut (.I0(n3006), .I1(n3006), .I2(n3017), 
            .I3(n40329), .O(n3105)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_6_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_6 (.CI(n40329), .I0(n3006), .I1(n3017), .CO(n40330));
    SB_LUT4 mod_5_add_1674_2_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(VCC_net), .O(n2456[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1674_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_2076_5_lut (.I0(n3007), .I1(n3007), .I2(n3017), 
            .I3(n40328), .O(n3106)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_5 (.CI(n40328), .I0(n3007), .I1(n3017), .CO(n40329));
    SB_LUT4 mod_5_add_2076_4_lut (.I0(n3008), .I1(n3008), .I2(n3017), 
            .I3(n40327), .O(n3107)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_2076_4 (.CI(n40327), .I0(n3008), .I1(n3017), .CO(n40328));
    SB_CARRY mod_5_add_1674_2 (.CI(VCC_net), .I0(bit_ctr[11]), .I1(GND_net), 
            .CO(n40677));
    SB_LUT4 mod_5_add_2076_3_lut (.I0(n30593), .I1(n30593), .I2(n51407), 
            .I3(n40326), .O(n3108)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_3_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_3 (.CI(n40326), .I0(n30593), .I1(n51407), 
            .CO(n40327));
    SB_LUT4 mod_5_add_2076_2_lut (.I0(bit_ctr[5]), .I1(bit_ctr[5]), .I2(n51407), 
            .I3(VCC_net), .O(n3109)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2076_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_2076_2 (.CI(VCC_net), .I0(bit_ctr[5]), .I1(n51407), 
            .CO(n40326));
    SB_LUT4 mod_5_add_1741_23_lut (.I0(n2522), .I1(n2489), .I2(VCC_net), 
            .I3(n40676), .O(n2588)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_23_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_33_lut (.I0(GND_net), .I1(bit_ctr[31]), .I2(GND_net), 
            .I3(n39074), .O(n255[31])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_32_lut (.I0(GND_net), .I1(bit_ctr[30]), .I2(GND_net), 
            .I3(n39073), .O(n255[30])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_32_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_22_lut (.I0(GND_net), .I1(n2490), .I2(VCC_net), 
            .I3(n40675), .O(n2555[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_22 (.CI(n40675), .I0(n2490), .I1(VCC_net), 
            .CO(n40676));
    SB_LUT4 mod_5_add_1741_21_lut (.I0(GND_net), .I1(n2491), .I2(VCC_net), 
            .I3(n40674), .O(n2555[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_21 (.CI(n40674), .I0(n2491), .I1(VCC_net), 
            .CO(n40675));
    SB_LUT4 mod_5_add_1741_20_lut (.I0(GND_net), .I1(n2492), .I2(VCC_net), 
            .I3(n40673), .O(n2555[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_20 (.CI(n40673), .I0(n2492), .I1(VCC_net), 
            .CO(n40674));
    SB_LUT4 mod_5_add_1741_19_lut (.I0(GND_net), .I1(n2493), .I2(VCC_net), 
            .I3(n40672), .O(n2555[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_19 (.CI(n40672), .I0(n2493), .I1(VCC_net), 
            .CO(n40673));
    SB_LUT4 mod_5_add_1741_18_lut (.I0(GND_net), .I1(n2494), .I2(VCC_net), 
            .I3(n40671), .O(n2555[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_18 (.CI(n40671), .I0(n2494), .I1(VCC_net), 
            .CO(n40672));
    SB_LUT4 mod_5_add_1741_17_lut (.I0(GND_net), .I1(n2495), .I2(VCC_net), 
            .I3(n40670), .O(n2555[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_17 (.CI(n40670), .I0(n2495), .I1(VCC_net), 
            .CO(n40671));
    SB_LUT4 mod_5_add_1741_16_lut (.I0(GND_net), .I1(n2496), .I2(VCC_net), 
            .I3(n40669), .O(n2555[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_32 (.CI(n39073), .I0(bit_ctr[30]), .I1(GND_net), .CO(n39074));
    SB_CARRY mod_5_add_1741_16 (.CI(n40669), .I0(n2496), .I1(VCC_net), 
            .CO(n40670));
    SB_LUT4 mod_5_add_1741_15_lut (.I0(GND_net), .I1(n2497), .I2(VCC_net), 
            .I3(n40668), .O(n2555[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_15 (.CI(n40668), .I0(n2497), .I1(VCC_net), 
            .CO(n40669));
    SB_LUT4 mod_5_add_1741_14_lut (.I0(GND_net), .I1(n2498), .I2(VCC_net), 
            .I3(n40667), .O(n2555[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_14 (.CI(n40667), .I0(n2498), .I1(VCC_net), 
            .CO(n40668));
    SB_LUT4 bit_ctr_0__bdd_4_lut (.I0(bit_ctr[0]), .I1(neopxl_color[2]), 
            .I2(neopxl_color[3]), .I3(bit_ctr[1]), .O(n51609));
    defparam bit_ctr_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n51609_bdd_4_lut (.I0(n51609), .I1(neopxl_color[1]), .I2(neopxl_color[0]), 
            .I3(bit_ctr[1]), .O(n51612));
    defparam n51609_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i29934_4_lut (.I0(n26525), .I1(n40998), .I2(n44851), .I3(\state[0] ), 
            .O(n34629));   // verilog/neopixel.v(36[4] 116[11])
    defparam i29934_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 equal_418_i8_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(start), 
            .I2(GND_net), .I3(GND_net), .O(n26634));
    defparam equal_418_i8_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i2_2_lut_adj_1598 (.I0(one_wire_N_579[2]), .I1(n4), .I2(GND_net), 
            .I3(GND_net), .O(n40998));
    defparam i2_2_lut_adj_1598.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_1599 (.I0(one_wire_N_579[2]), .I1(one_wire_N_579[3]), 
            .I2(GND_net), .I3(GND_net), .O(n44851));
    defparam i1_2_lut_adj_1599.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1600 (.I0(one_wire_N_579[5]), .I1(one_wire_N_579[4]), 
            .I2(GND_net), .I3(GND_net), .O(n48315));   // verilog/neopixel.v(104[14:39])
    defparam i1_2_lut_adj_1600.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1601 (.I0(one_wire_N_579[8]), .I1(one_wire_N_579[7]), 
            .I2(one_wire_N_579[6]), .I3(n48315), .O(n48321));   // verilog/neopixel.v(104[14:39])
    defparam i1_4_lut_adj_1601.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_31_lut (.I0(GND_net), .I1(bit_ctr[29]), .I2(GND_net), 
            .I3(n39072), .O(n255[29])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_31_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1749_3_lut (.I0(n2495), .I1(n2555[25]), .I2(n2522), 
            .I3(GND_net), .O(n2594));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1749_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_21_31 (.CI(n39072), .I0(bit_ctr[29]), .I1(GND_net), .CO(n39073));
    SB_LUT4 mod_5_i1755_3_lut (.I0(n2501), .I1(n2555[19]), .I2(n2522), 
            .I3(GND_net), .O(n2600));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1755_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1741_13_lut (.I0(GND_net), .I1(n2499), .I2(VCC_net), 
            .I3(n40666), .O(n2555[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_13 (.CI(n40666), .I0(n2499), .I1(VCC_net), 
            .CO(n40667));
    SB_LUT4 mod_5_add_1741_12_lut (.I0(GND_net), .I1(n2500), .I2(VCC_net), 
            .I3(n40665), .O(n2555[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_12 (.CI(n40665), .I0(n2500), .I1(VCC_net), 
            .CO(n40666));
    SB_LUT4 mod_5_i1757_3_lut (.I0(n2503), .I1(n2555[17]), .I2(n2522), 
            .I3(GND_net), .O(n2602));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1757_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1758_3_lut (.I0(n2504), .I1(n2555[16]), .I2(n2522), 
            .I3(GND_net), .O(n2603));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1758_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1759_3_lut (.I0(n2505), .I1(n2555[15]), .I2(n2522), 
            .I3(GND_net), .O(n2604));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1759_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1762_3_lut (.I0(n2508), .I1(n2555[12]), .I2(n2522), 
            .I3(GND_net), .O(n2607));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1762_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1751_3_lut (.I0(n2497), .I1(n2555[23]), .I2(n2522), 
            .I3(GND_net), .O(n2596));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1751_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1747_3_lut (.I0(n2493), .I1(n2555[27]), .I2(n2522), 
            .I3(GND_net), .O(n2592));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1747_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1741_11_lut (.I0(GND_net), .I1(n2501), .I2(VCC_net), 
            .I3(n40664), .O(n2555[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_11 (.CI(n40664), .I0(n2501), .I1(VCC_net), 
            .CO(n40665));
    SB_LUT4 mod_5_add_1741_10_lut (.I0(GND_net), .I1(n2502), .I2(VCC_net), 
            .I3(n40663), .O(n2555[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_10 (.CI(n40663), .I0(n2502), .I1(VCC_net), 
            .CO(n40664));
    SB_LUT4 add_21_30_lut (.I0(GND_net), .I1(bit_ctr[28]), .I2(GND_net), 
            .I3(n39071), .O(n255[28])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_30_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1741_9_lut (.I0(GND_net), .I1(n2503), .I2(VCC_net), 
            .I3(n40662), .O(n2555[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_9 (.CI(n40662), .I0(n2503), .I1(VCC_net), 
            .CO(n40663));
    SB_LUT4 mod_5_add_1741_8_lut (.I0(GND_net), .I1(n2504), .I2(VCC_net), 
            .I3(n40661), .O(n2555[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_8 (.CI(n40661), .I0(n2504), .I1(VCC_net), 
            .CO(n40662));
    SB_LUT4 mod_5_add_1741_7_lut (.I0(GND_net), .I1(n2505), .I2(VCC_net), 
            .I3(n40660), .O(n2555[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i1760_3_lut (.I0(n2506), .I1(n2555[14]), .I2(n2522), 
            .I3(GND_net), .O(n2605));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1760_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1741_7 (.CI(n40660), .I0(n2505), .I1(VCC_net), 
            .CO(n40661));
    SB_LUT4 mod_5_add_1741_6_lut (.I0(GND_net), .I1(n2506), .I2(VCC_net), 
            .I3(n40659), .O(n2555[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_6 (.CI(n40659), .I0(n2506), .I1(VCC_net), 
            .CO(n40660));
    SB_LUT4 mod_5_add_1741_5_lut (.I0(GND_net), .I1(n2507), .I2(VCC_net), 
            .I3(n40658), .O(n2555[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_5 (.CI(n40658), .I0(n2507), .I1(VCC_net), 
            .CO(n40659));
    SB_CARRY add_21_30 (.CI(n39071), .I0(bit_ctr[28]), .I1(GND_net), .CO(n39072));
    SB_LUT4 mod_5_add_1741_4_lut (.I0(GND_net), .I1(n2508), .I2(VCC_net), 
            .I3(n40657), .O(n2555[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_4 (.CI(n40657), .I0(n2508), .I1(VCC_net), 
            .CO(n40658));
    SB_LUT4 mod_5_i1744_3_lut (.I0(n2490), .I1(n2555[30]), .I2(n2522), 
            .I3(GND_net), .O(n2589));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1744_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1752_3_lut (.I0(n2498), .I1(n2555[22]), .I2(n2522), 
            .I3(GND_net), .O(n2597));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1752_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1741_3_lut (.I0(GND_net), .I1(n2509), .I2(GND_net), 
            .I3(n40656), .O(n2555[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_3 (.CI(n40656), .I0(n2509), .I1(GND_net), 
            .CO(n40657));
    SB_LUT4 mod_5_i1764_3_lut (.I0(bit_ctr[10]), .I1(n2555[10]), .I2(n2522), 
            .I3(GND_net), .O(n2609));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1764_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1741_2_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(VCC_net), .O(n2555[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1741_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1741_2 (.CI(VCC_net), .I0(bit_ctr[10]), .I1(GND_net), 
            .CO(n40656));
    SB_LUT4 mod_5_add_1808_24_lut (.I0(n2588), .I1(n2588), .I2(n2621), 
            .I3(n40655), .O(n2687)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_24_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_add_1808_23_lut (.I0(n2589), .I1(n2589), .I2(n2621), 
            .I3(n40654), .O(n2688)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_23_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_23 (.CI(n40654), .I0(n2589), .I1(n2621), .CO(n40655));
    SB_LUT4 mod_5_i1745_3_lut (.I0(n2491), .I1(n2555[29]), .I2(n2522), 
            .I3(GND_net), .O(n2590));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1745_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1808_22_lut (.I0(n2590), .I1(n2590), .I2(n2621), 
            .I3(n40653), .O(n2689)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_22_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_22 (.CI(n40653), .I0(n2590), .I1(n2621), .CO(n40654));
    SB_LUT4 mod_5_i1748_3_lut (.I0(n2494), .I1(n2555[26]), .I2(n2522), 
            .I3(GND_net), .O(n2593));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1748_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1808_21_lut (.I0(n2591), .I1(n2591), .I2(n2621), 
            .I3(n40652), .O(n2690)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_21_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 mod_5_i1750_3_lut (.I0(n2496), .I1(n2555[24]), .I2(n2522), 
            .I3(GND_net), .O(n2595));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1750_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1753_3_lut (.I0(n2499), .I1(n2555[21]), .I2(n2522), 
            .I3(GND_net), .O(n2598));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1753_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1761_3_lut (.I0(n2507), .I1(n2555[13]), .I2(n2522), 
            .I3(GND_net), .O(n2606));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1761_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1808_21 (.CI(n40652), .I0(n2591), .I1(n2621), .CO(n40653));
    SB_LUT4 add_21_29_lut (.I0(GND_net), .I1(bit_ctr[27]), .I2(GND_net), 
            .I3(n39070), .O(n255[27])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_29 (.CI(n39070), .I0(bit_ctr[27]), .I1(GND_net), .CO(n39071));
    SB_LUT4 mod_5_i1756_3_lut (.I0(n2502), .I1(n2555[18]), .I2(n2522), 
            .I3(GND_net), .O(n2601));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1756_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1746_3_lut (.I0(n2492), .I1(n2555[28]), .I2(n2522), 
            .I3(GND_net), .O(n2591));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1746_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1763_3_lut (.I0(n2509), .I1(n2555[11]), .I2(n2522), 
            .I3(GND_net), .O(n2608));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1763_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1602 (.I0(one_wire_N_579[10]), .I1(n26681), .I2(one_wire_N_579[9]), 
            .I3(n48321), .O(n26525));   // verilog/neopixel.v(104[14:39])
    defparam i1_4_lut_adj_1602.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_28_lut (.I0(GND_net), .I1(bit_ctr[26]), .I2(GND_net), 
            .I3(n39069), .O(n255[26])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_28 (.CI(n39069), .I0(bit_ctr[26]), .I1(GND_net), .CO(n39070));
    SB_LUT4 mod_5_i1754_3_lut (.I0(n2500), .I1(n2555[20]), .I2(n2522), 
            .I3(GND_net), .O(n2599));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1754_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i12_4_lut_adj_1603 (.I0(n2599), .I1(n2608), .I2(n2591), .I3(n2601), 
            .O(n34));
    defparam i12_4_lut_adj_1603.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1604 (.I0(n2606), .I1(n2598), .I2(n2595), .I3(n2593), 
            .O(n38_adj_4821));
    defparam i16_4_lut_adj_1604.LUT_INIT = 16'hfffe;
    SB_LUT4 add_21_27_lut (.I0(GND_net), .I1(bit_ctr[25]), .I2(GND_net), 
            .I3(n39068), .O(n255[25])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_27_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i7_3_lut_adj_1605 (.I0(n2590), .I1(bit_ctr[9]), .I2(n2609), 
            .I3(GND_net), .O(n29_adj_4822));
    defparam i7_3_lut_adj_1605.LUT_INIT = 16'heaea;
    SB_LUT4 i14_4_lut_adj_1606 (.I0(n2597), .I1(n2588), .I2(n2589), .I3(n2605), 
            .O(n36_adj_4823));
    defparam i14_4_lut_adj_1606.LUT_INIT = 16'hfffe;
    SB_LUT4 i30081_4_lut (.I0(n26525), .I1(n44851), .I2(n40998), .I3(\state[0] ), 
            .O(n44971));
    defparam i30081_4_lut.LUT_INIT = 16'hfaee;
    SB_LUT4 i20_4_lut_adj_1607 (.I0(\neo_pixel_transmitter.done ), .I1(\state[1] ), 
            .I2(start), .I3(n44971), .O(n7_adj_4824));
    defparam i20_4_lut_adj_1607.LUT_INIT = 16'hcecf;
    SB_LUT4 i1_4_lut_adj_1608 (.I0(n26634), .I1(n7_adj_4824), .I2(n34629), 
            .I3(\state[1] ), .O(n43085));
    defparam i1_4_lut_adj_1608.LUT_INIT = 16'hcc8c;
    SB_LUT4 bit_ctr_0__bdd_4_lut_36620 (.I0(bit_ctr[0]), .I1(neopxl_color[6]), 
            .I2(neopxl_color[7]), .I3(bit_ctr[1]), .O(n51525));
    defparam bit_ctr_0__bdd_4_lut_36620.LUT_INIT = 16'he4aa;
    SB_LUT4 n51525_bdd_4_lut (.I0(n51525), .I1(neopxl_color[5]), .I2(neopxl_color[4]), 
            .I3(bit_ctr[1]), .O(n51528));
    defparam n51525_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 mod_5_add_1808_20_lut (.I0(n2592), .I1(n2592), .I2(n2621), 
            .I3(n40651), .O(n2691)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_20_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 i13_4_lut_adj_1609 (.I0(n2592), .I1(n2596), .I2(n2607), .I3(n2604), 
            .O(n35));
    defparam i13_4_lut_adj_1609.LUT_INIT = 16'hfffe;
    SB_CARRY mod_5_add_1808_20 (.CI(n40651), .I0(n2592), .I1(n2621), .CO(n40652));
    SB_LUT4 i17_3_lut (.I0(n2603), .I1(n34), .I2(n2602), .I3(GND_net), 
            .O(n39_adj_4825));
    defparam i17_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i19_4_lut_adj_1610 (.I0(n29_adj_4822), .I1(n38_adj_4821), .I2(n2600), 
            .I3(n2594), .O(n41_adj_4826));
    defparam i19_4_lut_adj_1610.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1611 (.I0(n41_adj_4826), .I1(n39_adj_4825), .I2(n35), 
            .I3(n36_adj_4823), .O(n2621));
    defparam i21_4_lut_adj_1611.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_add_1808_19_lut (.I0(n2593), .I1(n2593), .I2(n2621), 
            .I3(n40650), .O(n2692)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_19_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_19 (.CI(n40650), .I0(n2593), .I1(n2621), .CO(n40651));
    SB_LUT4 mod_5_add_1808_18_lut (.I0(n2594), .I1(n2594), .I2(n2621), 
            .I3(n40649), .O(n2693)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_18_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_18 (.CI(n40649), .I0(n2594), .I1(n2621), .CO(n40650));
    SB_LUT4 mod_5_add_1808_17_lut (.I0(n2595), .I1(n2595), .I2(n2621), 
            .I3(n40648), .O(n2694)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_17_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_17 (.CI(n40648), .I0(n2595), .I1(n2621), .CO(n40649));
    SB_LUT4 mod_5_add_1808_16_lut (.I0(n2596), .I1(n2596), .I2(n2621), 
            .I3(n40647), .O(n2695)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_16_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY add_21_27 (.CI(n39068), .I0(bit_ctr[25]), .I1(GND_net), .CO(n39069));
    SB_CARRY mod_5_add_1808_16 (.CI(n40647), .I0(n2596), .I1(n2621), .CO(n40648));
    SB_LUT4 add_21_26_lut (.I0(GND_net), .I1(bit_ctr[24]), .I2(GND_net), 
            .I3(n39067), .O(n255[24])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1808_15_lut (.I0(n2597), .I1(n2597), .I2(n2621), 
            .I3(n40646), .O(n2696)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_15_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_15 (.CI(n40646), .I0(n2597), .I1(n2621), .CO(n40647));
    SB_LUT4 mod_5_add_1808_14_lut (.I0(n2598), .I1(n2598), .I2(n2621), 
            .I3(n40645), .O(n2697)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_14_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_14 (.CI(n40645), .I0(n2598), .I1(n2621), .CO(n40646));
    SB_LUT4 mod_5_add_1808_13_lut (.I0(n2599), .I1(n2599), .I2(n2621), 
            .I3(n40644), .O(n2698)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_13_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_13 (.CI(n40644), .I0(n2599), .I1(n2621), .CO(n40645));
    SB_LUT4 mod_5_add_1808_12_lut (.I0(n2600), .I1(n2600), .I2(n2621), 
            .I3(n40643), .O(n2699)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_12_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_12 (.CI(n40643), .I0(n2600), .I1(n2621), .CO(n40644));
    SB_LUT4 mod_5_add_1808_11_lut (.I0(n2601), .I1(n2601), .I2(n2621), 
            .I3(n40642), .O(n2700)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_11_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_11 (.CI(n40642), .I0(n2601), .I1(n2621), .CO(n40643));
    SB_LUT4 mod_5_add_1808_10_lut (.I0(n2602), .I1(n2602), .I2(n2621), 
            .I3(n40641), .O(n2701)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_10_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_10 (.CI(n40641), .I0(n2602), .I1(n2621), .CO(n40642));
    SB_LUT4 mod_5_add_1808_9_lut (.I0(n2603), .I1(n2603), .I2(n2621), 
            .I3(n40640), .O(n2702)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_9_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_9 (.CI(n40640), .I0(n2603), .I1(n2621), .CO(n40641));
    SB_CARRY add_21_26 (.CI(n39067), .I0(bit_ctr[24]), .I1(GND_net), .CO(n39068));
    SB_LUT4 mod_5_add_1808_8_lut (.I0(n2604), .I1(n2604), .I2(n2621), 
            .I3(n40639), .O(n2703)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_8_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_8 (.CI(n40639), .I0(n2604), .I1(n2621), .CO(n40640));
    SB_LUT4 mod_5_add_1808_7_lut (.I0(n2605), .I1(n2605), .I2(n2621), 
            .I3(n40638), .O(n2704)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_7_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_7 (.CI(n40638), .I0(n2605), .I1(n2621), .CO(n40639));
    SB_LUT4 mod_5_add_1808_6_lut (.I0(n2606), .I1(n2606), .I2(n2621), 
            .I3(n40637), .O(n2705)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_6_lut.LUT_INIT = 16'hCA3A;
    SB_LUT4 add_21_25_lut (.I0(GND_net), .I1(bit_ctr[23]), .I2(GND_net), 
            .I3(n39066), .O(n255[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1808_6 (.CI(n40637), .I0(n2606), .I1(n2621), .CO(n40638));
    SB_LUT4 sub_14_add_2_33_lut (.I0(n48313), .I1(timer[31]), .I2(n1[31]), 
            .I3(n39209), .O(n26681)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_33_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 mod_5_add_1808_5_lut (.I0(n2607), .I1(n2607), .I2(n2621), 
            .I3(n40636), .O(n2706)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_5_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_5 (.CI(n40636), .I0(n2607), .I1(n2621), .CO(n40637));
    SB_LUT4 mod_5_add_1808_4_lut (.I0(n2608), .I1(n2608), .I2(n2621), 
            .I3(n40635), .O(n2707)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_4_lut.LUT_INIT = 16'hCA3A;
    SB_CARRY mod_5_add_1808_4 (.CI(n40635), .I0(n2608), .I1(n2621), .CO(n40636));
    SB_LUT4 mod_5_add_1808_3_lut (.I0(n2609), .I1(n2609), .I2(n51408), 
            .I3(n40634), .O(n2708)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_3_lut.LUT_INIT = 16'hA3AC;
    SB_LUT4 sub_14_add_2_32_lut (.I0(n48311), .I1(timer[30]), .I2(n1[30]), 
            .I3(n39208), .O(n48313)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_32_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1808_3 (.CI(n40634), .I0(n2609), .I1(n51408), .CO(n40635));
    SB_LUT4 mod_5_add_1808_2_lut (.I0(bit_ctr[9]), .I1(bit_ctr[9]), .I2(n51408), 
            .I3(VCC_net), .O(n2709)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1808_2_lut.LUT_INIT = 16'hA3AC;
    SB_CARRY mod_5_add_1808_2 (.CI(VCC_net), .I0(bit_ctr[9]), .I1(n51408), 
            .CO(n40634));
    SB_LUT4 mod_5_add_1875_25_lut (.I0(n2720), .I1(n2687), .I2(VCC_net), 
            .I3(n40633), .O(n2786)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_25_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_1875_24_lut (.I0(GND_net), .I1(n2688), .I2(VCC_net), 
            .I3(n40632), .O(n2753[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_24 (.CI(n40632), .I0(n2688), .I1(VCC_net), 
            .CO(n40633));
    SB_LUT4 mod_5_add_1875_23_lut (.I0(GND_net), .I1(n2689), .I2(VCC_net), 
            .I3(n40631), .O(n2753[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_23 (.CI(n40631), .I0(n2689), .I1(VCC_net), 
            .CO(n40632));
    SB_LUT4 mod_5_add_1875_22_lut (.I0(GND_net), .I1(n2690), .I2(VCC_net), 
            .I3(n40630), .O(n2753[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_22 (.CI(n40630), .I0(n2690), .I1(VCC_net), 
            .CO(n40631));
    SB_LUT4 mod_5_i946_3_lut (.I0(n1308), .I1(n1367[24]), .I2(n1334), 
            .I3(GND_net), .O(n1407));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i946_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i945_3_lut (.I0(n1307), .I1(n1367[25]), .I2(n1334), 
            .I3(GND_net), .O(n1406));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i944_3_lut (.I0(n1306), .I1(n1367[26]), .I2(n1334), 
            .I3(GND_net), .O(n1405));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i944_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i941_3_lut (.I0(n1303), .I1(n1367[29]), .I2(n1334), 
            .I3(GND_net), .O(n1402));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i941_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1875_21_lut (.I0(GND_net), .I1(n2691), .I2(VCC_net), 
            .I3(n40629), .O(n2753[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_21 (.CI(n40629), .I0(n2691), .I1(VCC_net), 
            .CO(n40630));
    SB_LUT4 mod_5_i948_3_lut (.I0(bit_ctr[22]), .I1(n1367[22]), .I2(n1334), 
            .I3(GND_net), .O(n1409));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_add_1875_20_lut (.I0(GND_net), .I1(n2692), .I2(VCC_net), 
            .I3(n40628), .O(n2753[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i942_3_lut (.I0(n1304), .I1(n1367[28]), .I2(n1334), 
            .I3(GND_net), .O(n1403));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i942_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1875_20 (.CI(n40628), .I0(n2692), .I1(VCC_net), 
            .CO(n40629));
    SB_LUT4 mod_5_add_1875_19_lut (.I0(GND_net), .I1(n2693), .I2(VCC_net), 
            .I3(n40627), .O(n2753[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i943_3_lut (.I0(n1305), .I1(n1367[27]), .I2(n1334), 
            .I3(GND_net), .O(n1404));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i943_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1875_19 (.CI(n40627), .I0(n2693), .I1(VCC_net), 
            .CO(n40628));
    SB_LUT4 i5_3_lut (.I0(n1307), .I1(n1302), .I2(n1301), .I3(GND_net), 
            .O(n14_adj_4827));   // verilog/neopixel.v(22[26:36])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_2_lut_adj_1612 (.I0(n1305), .I1(n1306), .I2(GND_net), .I3(GND_net), 
            .O(n12_adj_4828));   // verilog/neopixel.v(22[26:36])
    defparam i3_2_lut_adj_1612.LUT_INIT = 16'heeee;
    SB_LUT4 mod_5_add_1875_18_lut (.I0(GND_net), .I1(n2694), .I2(VCC_net), 
            .I3(n40626), .O(n2753[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_25 (.CI(n39066), .I0(bit_ctr[23]), .I1(GND_net), .CO(n39067));
    SB_CARRY mod_5_add_1875_18 (.CI(n40626), .I0(n2694), .I1(VCC_net), 
            .CO(n40627));
    SB_LUT4 mod_5_add_1875_17_lut (.I0(GND_net), .I1(n2695), .I2(VCC_net), 
            .I3(n40625), .O(n2753[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_17 (.CI(n40625), .I0(n2695), .I1(VCC_net), 
            .CO(n40626));
    SB_LUT4 mod_5_add_1875_16_lut (.I0(GND_net), .I1(n2696), .I2(VCC_net), 
            .I3(n40624), .O(n2753[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_16 (.CI(n40624), .I0(n2696), .I1(VCC_net), 
            .CO(n40625));
    SB_LUT4 i7_4_lut_adj_1613 (.I0(bit_ctr[22]), .I1(n14_adj_4827), .I2(n1308), 
            .I3(n1309), .O(n16_adj_4829));   // verilog/neopixel.v(22[26:36])
    defparam i7_4_lut_adj_1613.LUT_INIT = 16'hfefc;
    SB_LUT4 mod_5_add_1875_15_lut (.I0(GND_net), .I1(n2697), .I2(VCC_net), 
            .I3(n40623), .O(n2753[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_15 (.CI(n40623), .I0(n2697), .I1(VCC_net), 
            .CO(n40624));
    SB_LUT4 mod_5_add_1875_14_lut (.I0(GND_net), .I1(n2698), .I2(VCC_net), 
            .I3(n40622), .O(n2753[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i8_4_lut_adj_1614 (.I0(n1303), .I1(n16_adj_4829), .I2(n12_adj_4828), 
            .I3(n1304), .O(n1334));   // verilog/neopixel.v(22[26:36])
    defparam i8_4_lut_adj_1614.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i940_3_lut (.I0(n1302), .I1(n1367[30]), .I2(n1334), 
            .I3(GND_net), .O(n1401));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i940_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1875_14 (.CI(n40622), .I0(n2698), .I1(VCC_net), 
            .CO(n40623));
    SB_LUT4 mod_5_add_1875_13_lut (.I0(GND_net), .I1(n2699), .I2(VCC_net), 
            .I3(n40621), .O(n2753[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_24_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(n39065), .O(n255[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i947_3_lut (.I0(n1309), .I1(n1367[23]), .I2(n1334), 
            .I3(GND_net), .O(n1408));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i947_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY mod_5_add_1875_13 (.CI(n40621), .I0(n2699), .I1(VCC_net), 
            .CO(n40622));
    SB_LUT4 i2_2_lut_adj_1615 (.I0(n1408), .I1(n1401), .I2(GND_net), .I3(GND_net), 
            .O(n12_adj_4830));   // verilog/neopixel.v(22[26:36])
    defparam i2_2_lut_adj_1615.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_1616 (.I0(bit_ctr[21]), .I1(n12_adj_4830), .I2(n1400), 
            .I3(n1409), .O(n16_adj_4831));   // verilog/neopixel.v(22[26:36])
    defparam i6_4_lut_adj_1616.LUT_INIT = 16'hfefc;
    SB_LUT4 i7_4_lut_adj_1617 (.I0(n1402), .I1(n1405), .I2(n1406), .I3(n1407), 
            .O(n17_adj_4832));   // verilog/neopixel.v(22[26:36])
    defparam i7_4_lut_adj_1617.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1618 (.I0(n17_adj_4832), .I1(n1404), .I2(n16_adj_4831), 
            .I3(n1403), .O(n1433));   // verilog/neopixel.v(22[26:36])
    defparam i9_4_lut_adj_1618.LUT_INIT = 16'hfffe;
    SB_CARRY sub_14_add_2_32 (.CI(n39208), .I0(timer[30]), .I1(n1[30]), 
            .CO(n39209));
    SB_LUT4 mod_5_add_1875_12_lut (.I0(GND_net), .I1(n2700), .I2(VCC_net), 
            .I3(n40620), .O(n2753[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_12 (.CI(n40620), .I0(n2700), .I1(VCC_net), 
            .CO(n40621));
    SB_LUT4 mod_5_add_1875_11_lut (.I0(GND_net), .I1(n2701), .I2(VCC_net), 
            .I3(n40619), .O(n2753[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_31_lut (.I0(n48309), .I1(timer[29]), .I2(n1[29]), 
            .I3(n39207), .O(n48311)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_31_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1875_11 (.CI(n40619), .I0(n2701), .I1(VCC_net), 
            .CO(n40620));
    SB_LUT4 mod_5_add_1875_10_lut (.I0(GND_net), .I1(n2702), .I2(VCC_net), 
            .I3(n40618), .O(n2753[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_10 (.CI(n40618), .I0(n2702), .I1(VCC_net), 
            .CO(n40619));
    SB_LUT4 mod_5_add_1875_9_lut (.I0(GND_net), .I1(n2703), .I2(VCC_net), 
            .I3(n40617), .O(n2753[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_9 (.CI(n40617), .I0(n2703), .I1(VCC_net), 
            .CO(n40618));
    SB_LUT4 mod_5_add_1875_8_lut (.I0(GND_net), .I1(n2704), .I2(VCC_net), 
            .I3(n40616), .O(n2753[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_8 (.CI(n40616), .I0(n2704), .I1(VCC_net), 
            .CO(n40617));
    SB_LUT4 mod_5_add_1875_7_lut (.I0(GND_net), .I1(n2705), .I2(VCC_net), 
            .I3(n40615), .O(n2753[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_7 (.CI(n40615), .I0(n2705), .I1(VCC_net), 
            .CO(n40616));
    SB_LUT4 mod_5_add_1875_6_lut (.I0(GND_net), .I1(n2706), .I2(VCC_net), 
            .I3(n40614), .O(n2753[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_6 (.CI(n40614), .I0(n2706), .I1(VCC_net), 
            .CO(n40615));
    SB_LUT4 mod_5_add_1875_5_lut (.I0(GND_net), .I1(n2707), .I2(VCC_net), 
            .I3(n40613), .O(n2753[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_5 (.CI(n40613), .I0(n2707), .I1(VCC_net), 
            .CO(n40614));
    SB_CARRY add_21_24 (.CI(n39065), .I0(bit_ctr[22]), .I1(GND_net), .CO(n39066));
    SB_LUT4 mod_5_add_1875_4_lut (.I0(GND_net), .I1(n2708), .I2(VCC_net), 
            .I3(n40612), .O(n2753[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_4 (.CI(n40612), .I0(n2708), .I1(VCC_net), 
            .CO(n40613));
    SB_LUT4 mod_5_add_1875_3_lut (.I0(GND_net), .I1(n2709), .I2(GND_net), 
            .I3(n40611), .O(n2753[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1875_3 (.CI(n40611), .I0(n2709), .I1(GND_net), 
            .CO(n40612));
    SB_LUT4 mod_5_add_1875_2_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(VCC_net), .O(n2753[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1875_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_31 (.CI(n39207), .I0(timer[29]), .I1(n1[29]), 
            .CO(n39208));
    SB_CARRY mod_5_add_1875_2 (.CI(VCC_net), .I0(bit_ctr[8]), .I1(GND_net), 
            .CO(n40611));
    SB_LUT4 mod_5_add_1942_26_lut (.I0(n2819), .I1(n2786), .I2(VCC_net), 
            .I3(n40610), .O(n2885)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_26_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_21_23_lut (.I0(GND_net), .I1(bit_ctr[21]), .I2(GND_net), 
            .I3(n39064), .O(n255[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_add_1942_25_lut (.I0(GND_net), .I1(n2787), .I2(VCC_net), 
            .I3(n40609), .O(n2852[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_23 (.CI(n39064), .I0(bit_ctr[21]), .I1(GND_net), .CO(n39065));
    SB_CARRY mod_5_add_1942_25 (.CI(n40609), .I0(n2787), .I1(VCC_net), 
            .CO(n40610));
    SB_LUT4 mod_5_add_1942_24_lut (.I0(GND_net), .I1(n2788), .I2(VCC_net), 
            .I3(n40608), .O(n2852[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_24 (.CI(n40608), .I0(n2788), .I1(VCC_net), 
            .CO(n40609));
    SB_LUT4 mod_5_add_1942_23_lut (.I0(GND_net), .I1(n2789), .I2(VCC_net), 
            .I3(n40607), .O(n2852[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_23 (.CI(n40607), .I0(n2789), .I1(VCC_net), 
            .CO(n40608));
    SB_LUT4 mod_5_add_1942_22_lut (.I0(GND_net), .I1(n2790), .I2(VCC_net), 
            .I3(n40606), .O(n2852[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_22 (.CI(n40606), .I0(n2790), .I1(VCC_net), 
            .CO(n40607));
    SB_LUT4 mod_5_add_1942_21_lut (.I0(GND_net), .I1(n2791), .I2(VCC_net), 
            .I3(n40605), .O(n2852[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_21 (.CI(n40605), .I0(n2791), .I1(VCC_net), 
            .CO(n40606));
    SB_LUT4 sub_14_inv_0_i1_1_lut (.I0(\neo_pixel_transmitter.t0 [0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[0]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_1942_20_lut (.I0(GND_net), .I1(n2792), .I2(VCC_net), 
            .I3(n40604), .O(n2852[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_20 (.CI(n40604), .I0(n2792), .I1(VCC_net), 
            .CO(n40605));
    SB_LUT4 mod_5_add_1942_19_lut (.I0(GND_net), .I1(n2793), .I2(VCC_net), 
            .I3(n40603), .O(n2852[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_22_lut (.I0(GND_net), .I1(bit_ctr[20]), .I2(GND_net), 
            .I3(n39063), .O(n255[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_19 (.CI(n40603), .I0(n2793), .I1(VCC_net), 
            .CO(n40604));
    SB_LUT4 mod_5_add_1942_18_lut (.I0(GND_net), .I1(n2794), .I2(VCC_net), 
            .I3(n40602), .O(n2852[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_18 (.CI(n40602), .I0(n2794), .I1(VCC_net), 
            .CO(n40603));
    SB_LUT4 mod_5_add_1942_17_lut (.I0(GND_net), .I1(n2795), .I2(VCC_net), 
            .I3(n40601), .O(n2852[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_17 (.CI(n40601), .I0(n2795), .I1(VCC_net), 
            .CO(n40602));
    SB_LUT4 mod_5_add_1942_16_lut (.I0(GND_net), .I1(n2796), .I2(VCC_net), 
            .I3(n40600), .O(n2852[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_16 (.CI(n40600), .I0(n2796), .I1(VCC_net), 
            .CO(n40601));
    SB_LUT4 mod_5_add_1942_15_lut (.I0(GND_net), .I1(n2797), .I2(VCC_net), 
            .I3(n40599), .O(n2852[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_15 (.CI(n40599), .I0(n2797), .I1(VCC_net), 
            .CO(n40600));
    SB_LUT4 mod_5_add_1942_14_lut (.I0(GND_net), .I1(n2798), .I2(VCC_net), 
            .I3(n40598), .O(n2852[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_14 (.CI(n40598), .I0(n2798), .I1(VCC_net), 
            .CO(n40599));
    SB_LUT4 mod_5_add_1942_13_lut (.I0(GND_net), .I1(n2799), .I2(VCC_net), 
            .I3(n40597), .O(n2852[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_30_lut (.I0(n48307), .I1(timer[28]), .I2(n1[28]), 
            .I3(n39206), .O(n48309)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_30_lut.LUT_INIT = 16'hebbe;
    SB_CARRY mod_5_add_1942_13 (.CI(n40597), .I0(n2799), .I1(VCC_net), 
            .CO(n40598));
    SB_LUT4 mod_5_add_1942_12_lut (.I0(GND_net), .I1(n2800), .I2(VCC_net), 
            .I3(n40596), .O(n2852[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_12 (.CI(n40596), .I0(n2800), .I1(VCC_net), 
            .CO(n40597));
    SB_LUT4 mod_5_add_1942_11_lut (.I0(GND_net), .I1(n2801), .I2(VCC_net), 
            .I3(n40595), .O(n2852[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_11 (.CI(n40595), .I0(n2801), .I1(VCC_net), 
            .CO(n40596));
    SB_LUT4 mod_5_add_1942_10_lut (.I0(GND_net), .I1(n2802), .I2(VCC_net), 
            .I3(n40594), .O(n2852[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_10 (.CI(n40594), .I0(n2802), .I1(VCC_net), 
            .CO(n40595));
    SB_LUT4 mod_5_add_1942_9_lut (.I0(GND_net), .I1(n2803), .I2(VCC_net), 
            .I3(n40593), .O(n2852[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_9 (.CI(n40593), .I0(n2803), .I1(VCC_net), 
            .CO(n40594));
    SB_LUT4 mod_5_add_1942_8_lut (.I0(GND_net), .I1(n2804), .I2(VCC_net), 
            .I3(n40592), .O(n2852[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_8 (.CI(n40592), .I0(n2804), .I1(VCC_net), 
            .CO(n40593));
    SB_LUT4 mod_5_add_1942_7_lut (.I0(GND_net), .I1(n2805), .I2(VCC_net), 
            .I3(n40591), .O(n2852[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_7 (.CI(n40591), .I0(n2805), .I1(VCC_net), 
            .CO(n40592));
    SB_LUT4 mod_5_add_1942_6_lut (.I0(GND_net), .I1(n2806), .I2(VCC_net), 
            .I3(n40590), .O(n2852[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_6 (.CI(n40590), .I0(n2806), .I1(VCC_net), 
            .CO(n40591));
    SB_LUT4 mod_5_add_1942_5_lut (.I0(GND_net), .I1(n2807), .I2(VCC_net), 
            .I3(n40589), .O(n2852[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_5 (.CI(n40589), .I0(n2807), .I1(VCC_net), 
            .CO(n40590));
    SB_LUT4 mod_5_add_1942_4_lut (.I0(GND_net), .I1(n2808), .I2(VCC_net), 
            .I3(n40588), .O(n2852[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_4 (.CI(n40588), .I0(n2808), .I1(VCC_net), 
            .CO(n40589));
    SB_LUT4 mod_5_add_1942_3_lut (.I0(GND_net), .I1(n2809), .I2(GND_net), 
            .I3(n40587), .O(n2852[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_1942_3 (.CI(n40587), .I0(n2809), .I1(GND_net), 
            .CO(n40588));
    SB_LUT4 mod_5_add_1942_2_lut (.I0(GND_net), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(VCC_net), .O(n2852[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_1942_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_2009_26 (.CI(n40585), .I0(n2886), .I1(VCC_net), 
            .CO(n40586));
    SB_CARRY sub_14_add_2_30 (.CI(n39206), .I0(timer[28]), .I1(n1[28]), 
            .CO(n39207));
    SB_LUT4 sub_14_add_2_29_lut (.I0(n48305), .I1(timer[27]), .I2(n1[27]), 
            .I3(n39205), .O(n48307)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_29_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_22 (.CI(n39063), .I0(bit_ctr[20]), .I1(GND_net), .CO(n39064));
    SB_CARRY mod_5_add_1942_2 (.CI(VCC_net), .I0(bit_ctr[7]), .I1(GND_net), 
            .CO(n40587));
    SB_CARRY sub_14_add_2_29 (.CI(n39205), .I0(timer[27]), .I1(n1[27]), 
            .CO(n39206));
    SB_LUT4 sub_14_add_2_28_lut (.I0(n48303), .I1(timer[26]), .I2(n1[26]), 
            .I3(n39204), .O(n48305)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_28_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_28 (.CI(n39204), .I0(timer[26]), .I1(n1[26]), 
            .CO(n39205));
    SB_LUT4 sub_14_inv_0_i2_1_lut (.I0(\neo_pixel_transmitter.t0 [1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[1]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_add_2009_27_lut (.I0(n2918), .I1(n2885), .I2(VCC_net), 
            .I3(n40586), .O(n2984)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_2009_26_lut (.I0(GND_net), .I1(n2886), .I2(VCC_net), 
            .I3(n40585), .O(n2951[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_2009_26_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_27_lut (.I0(n48301), .I1(timer[25]), .I2(n1[25]), 
            .I3(n39203), .O(n48303)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_27_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 add_21_21_lut (.I0(GND_net), .I1(bit_ctr[19]), .I2(GND_net), 
            .I3(n39062), .O(n255[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_inv_0_i3_1_lut (.I0(\neo_pixel_transmitter.t0 [2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[2]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_21_21 (.CI(n39062), .I0(bit_ctr[19]), .I1(GND_net), .CO(n39063));
    SB_CARRY sub_14_add_2_27 (.CI(n39203), .I0(timer[25]), .I1(n1[25]), 
            .CO(n39204));
    SB_LUT4 bit_ctr_1__bdd_4_lut (.I0(bit_ctr[1]), .I1(n49021), .I2(n49022), 
            .I3(bit_ctr[2]), .O(n51465));
    defparam bit_ctr_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n51465_bdd_4_lut (.I0(n51465), .I1(n48962), .I2(n48961), .I3(bit_ctr[2]), 
            .O(n51468));
    defparam n51465_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 add_21_20_lut (.I0(GND_net), .I1(bit_ctr[18]), .I2(GND_net), 
            .I3(n39061), .O(n255[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_20 (.CI(n39061), .I0(bit_ctr[18]), .I1(GND_net), .CO(n39062));
    SB_LUT4 add_21_19_lut (.I0(GND_net), .I1(bit_ctr[17]), .I2(GND_net), 
            .I3(n39060), .O(n255[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_26_lut (.I0(n48299), .I1(timer[24]), .I2(n1[24]), 
            .I3(n39202), .O(n48301)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_26_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 bit_ctr_1__bdd_4_lut_36503 (.I0(bit_ctr[1]), .I1(n48997), .I2(n48998), 
            .I3(bit_ctr[2]), .O(n51459));
    defparam bit_ctr_1__bdd_4_lut_36503.LUT_INIT = 16'he4aa;
    SB_LUT4 n51459_bdd_4_lut (.I0(n51459), .I1(n48995), .I2(n48994), .I3(bit_ctr[2]), 
            .O(n51462));
    defparam n51459_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_CARRY sub_14_add_2_26 (.CI(n39202), .I0(timer[24]), .I1(n1[24]), 
            .CO(n39203));
    SB_LUT4 sub_14_add_2_25_lut (.I0(n48297), .I1(timer[23]), .I2(n1[23]), 
            .I3(n39201), .O(n48299)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_25_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_25 (.CI(n39201), .I0(timer[23]), .I1(n1[23]), 
            .CO(n39202));
    SB_LUT4 i29962_2_lut (.I0(start), .I1(\state[1] ), .I2(GND_net), .I3(GND_net), 
            .O(n44847));
    defparam i29962_2_lut.LUT_INIT = 16'heeee;
    SB_DFFESS state_i0 (.Q(\state[0] ), .C(CLK_c), .E(n27916), .D(state_3__N_428[0]), 
            .S(n44839));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF timer_1546__i1 (.Q(timer[1]), .C(CLK_c), .D(n133[1]));   // verilog/neopixel.v(12[12:21])
    SB_LUT4 i35722_2_lut (.I0(\neo_pixel_transmitter.done ), .I1(\state[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n44118));
    defparam i35722_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 sub_14_add_2_24_lut (.I0(n48295), .I1(timer[22]), .I2(n1[22]), 
            .I3(n39200), .O(n48297)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_24_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_24 (.CI(n39200), .I0(timer[22]), .I1(n1[22]), 
            .CO(n39201));
    SB_LUT4 sub_14_add_2_23_lut (.I0(n48293), .I1(timer[21]), .I2(n1[21]), 
            .I3(n39199), .O(n48295)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_23_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_23 (.CI(n39199), .I0(timer[21]), .I1(n1[21]), 
            .CO(n39200));
    SB_CARRY add_21_19 (.CI(n39060), .I0(bit_ctr[17]), .I1(GND_net), .CO(n39061));
    SB_LUT4 sub_14_add_2_22_lut (.I0(n48291), .I1(timer[20]), .I2(n1[20]), 
            .I3(n39198), .O(n48293)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_22_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_22 (.CI(n39198), .I0(timer[20]), .I1(n1[20]), 
            .CO(n39199));
    SB_LUT4 add_21_18_lut (.I0(GND_net), .I1(bit_ctr[16]), .I2(GND_net), 
            .I3(n39059), .O(n255[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_18 (.CI(n39059), .I0(bit_ctr[16]), .I1(GND_net), .CO(n39060));
    SB_LUT4 add_21_17_lut (.I0(GND_net), .I1(bit_ctr[15]), .I2(GND_net), 
            .I3(n39058), .O(n255[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_17 (.CI(n39058), .I0(bit_ctr[15]), .I1(GND_net), .CO(n39059));
    SB_LUT4 add_21_16_lut (.I0(GND_net), .I1(bit_ctr[14]), .I2(GND_net), 
            .I3(n39057), .O(n255[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut_adj_1619 (.I0(one_wire_N_579[2]), .I1(n44118), .I2(one_wire_N_579[3]), 
            .I3(n4), .O(n103));
    defparam i1_4_lut_adj_1619.LUT_INIT = 16'h45cd;
    SB_LUT4 sub_14_add_2_21_lut (.I0(n48289), .I1(timer[19]), .I2(n1[19]), 
            .I3(n39197), .O(n48291)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_21_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_21 (.CI(n39197), .I0(timer[19]), .I1(n1[19]), 
            .CO(n39198));
    SB_LUT4 i6_4_lut_adj_1620 (.I0(one_wire_N_579[7]), .I1(one_wire_N_579[9]), 
            .I2(n44847), .I3(n103), .O(n16_adj_4833));
    defparam i6_4_lut_adj_1620.LUT_INIT = 16'h0100;
    SB_LUT4 i1_4_lut_adj_1621 (.I0(one_wire_N_579[8]), .I1(one_wire_N_579[4]), 
            .I2(n16_adj_4833), .I3(n26681), .O(n6_adj_4834));
    defparam i1_4_lut_adj_1621.LUT_INIT = 16'hffef;
    SB_LUT4 i4_4_lut (.I0(one_wire_N_579[10]), .I1(one_wire_N_579[6]), .I2(one_wire_N_579[5]), 
            .I3(n6_adj_4834), .O(n51632));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_747_Mux_0_i3_3_lut (.I0(start), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[1] ), .I3(GND_net), .O(\neo_pixel_transmitter.done_N_636 ));   // verilog/neopixel.v(36[4] 116[11])
    defparam mux_747_Mux_0_i3_3_lut.LUT_INIT = 16'hc1c1;
    SB_LUT4 mod_5_add_937_11_lut (.I0(n1334), .I1(n1301), .I2(VCC_net), 
            .I3(n40161), .O(n1400)) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_11_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mod_5_add_937_10_lut (.I0(GND_net), .I1(n1302), .I2(VCC_net), 
            .I3(n40160), .O(n1367[30])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_10 (.CI(n40160), .I0(n1302), .I1(VCC_net), 
            .CO(n40161));
    SB_LUT4 mod_5_add_937_9_lut (.I0(GND_net), .I1(n1303), .I2(VCC_net), 
            .I3(n40159), .O(n1367[29])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_9 (.CI(n40159), .I0(n1303), .I1(VCC_net), .CO(n40160));
    SB_LUT4 mod_5_add_937_8_lut (.I0(GND_net), .I1(n1304), .I2(VCC_net), 
            .I3(n40158), .O(n1367[28])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_8 (.CI(n40158), .I0(n1304), .I1(VCC_net), .CO(n40159));
    SB_LUT4 mod_5_add_937_7_lut (.I0(GND_net), .I1(n1305), .I2(VCC_net), 
            .I3(n40157), .O(n1367[27])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_7 (.CI(n40157), .I0(n1305), .I1(VCC_net), .CO(n40158));
    SB_LUT4 mod_5_add_937_6_lut (.I0(GND_net), .I1(n1306), .I2(VCC_net), 
            .I3(n40156), .O(n1367[26])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_6 (.CI(n40156), .I0(n1306), .I1(VCC_net), .CO(n40157));
    SB_LUT4 mod_5_add_937_5_lut (.I0(GND_net), .I1(n1307), .I2(VCC_net), 
            .I3(n40155), .O(n1367[25])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_5 (.CI(n40155), .I0(n1307), .I1(VCC_net), .CO(n40156));
    SB_LUT4 mod_5_add_937_4_lut (.I0(GND_net), .I1(n1308), .I2(VCC_net), 
            .I3(n40154), .O(n1367[24])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_4 (.CI(n40154), .I0(n1308), .I1(VCC_net), .CO(n40155));
    SB_LUT4 mod_5_add_937_3_lut (.I0(GND_net), .I1(n1309), .I2(GND_net), 
            .I3(n40153), .O(n1367[23])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_3 (.CI(n40153), .I0(n1309), .I1(GND_net), .CO(n40154));
    SB_DFFE start_103 (.Q(start), .C(CLK_c), .E(VCC_net), .D(n42985));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 mod_5_add_937_2_lut (.I0(GND_net), .I1(bit_ctr[22]), .I2(GND_net), 
            .I3(VCC_net), .O(n1367[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mod_5_add_937_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_16 (.CI(n39057), .I0(bit_ctr[14]), .I1(GND_net), .CO(n39058));
    SB_LUT4 add_21_15_lut (.I0(GND_net), .I1(bit_ctr[13]), .I2(GND_net), 
            .I3(n39056), .O(n255[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mod_5_add_937_2 (.CI(VCC_net), .I0(bit_ctr[22]), .I1(GND_net), 
            .CO(n40153));
    SB_LUT4 sub_14_add_2_20_lut (.I0(n48287), .I1(timer[18]), .I2(n1[18]), 
            .I3(n39196), .O(n48289)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_20_lut.LUT_INIT = 16'hebbe;
    SB_CARRY add_21_15 (.CI(n39056), .I0(bit_ctr[13]), .I1(GND_net), .CO(n39057));
    SB_CARRY sub_14_add_2_20 (.CI(n39196), .I0(timer[18]), .I1(n1[18]), 
            .CO(n39197));
    SB_LUT4 add_21_14_lut (.I0(GND_net), .I1(bit_ctr[12]), .I2(GND_net), 
            .I3(n39055), .O(n255[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_14 (.CI(n39055), .I0(bit_ctr[12]), .I1(GND_net), .CO(n39056));
    SB_LUT4 sub_14_add_2_19_lut (.I0(n48285), .I1(timer[17]), .I2(n1[17]), 
            .I3(n39195), .O(n48287)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_19_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_19 (.CI(n39195), .I0(timer[17]), .I1(n1[17]), 
            .CO(n39196));
    SB_DFFESR bit_ctr_i0_i0 (.Q(bit_ctr[0]), .C(CLK_c), .E(n27743), .D(n255[0]), 
            .R(n28088));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 sub_14_add_2_18_lut (.I0(n48283), .I1(timer[16]), .I2(n1[16]), 
            .I3(n39194), .O(n48285)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_18_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_18 (.CI(n39194), .I0(timer[16]), .I1(n1[16]), 
            .CO(n39195));
    SB_LUT4 sub_14_add_2_17_lut (.I0(n48281), .I1(timer[15]), .I2(n1[15]), 
            .I3(n39193), .O(n48283)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_17_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_17 (.CI(n39193), .I0(timer[15]), .I1(n1[15]), 
            .CO(n39194));
    SB_LUT4 sub_14_add_2_16_lut (.I0(n48279), .I1(timer[14]), .I2(n1[14]), 
            .I3(n39192), .O(n48281)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_16_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_16 (.CI(n39192), .I0(timer[14]), .I1(n1[14]), 
            .CO(n39193));
    SB_LUT4 add_21_13_lut (.I0(GND_net), .I1(bit_ctr[11]), .I2(GND_net), 
            .I3(n39054), .O(n255[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_15_lut (.I0(n48277), .I1(timer[13]), .I2(n1[13]), 
            .I3(n39191), .O(n48279)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_15_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_15 (.CI(n39191), .I0(timer[13]), .I1(n1[13]), 
            .CO(n39192));
    SB_LUT4 sub_14_add_2_14_lut (.I0(one_wire_N_579[11]), .I1(timer[12]), 
            .I2(n1[12]), .I3(n39190), .O(n48277)) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_14_lut.LUT_INIT = 16'hebbe;
    SB_CARRY sub_14_add_2_14 (.CI(n39190), .I0(timer[12]), .I1(n1[12]), 
            .CO(n39191));
    SB_DFF timer_1546__i2 (.Q(timer[2]), .C(CLK_c), .D(n133[2]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i3 (.Q(timer[3]), .C(CLK_c), .D(n133[3]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i4 (.Q(timer[4]), .C(CLK_c), .D(n133[4]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i5 (.Q(timer[5]), .C(CLK_c), .D(n133[5]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i6 (.Q(timer[6]), .C(CLK_c), .D(n133[6]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i7 (.Q(timer[7]), .C(CLK_c), .D(n133[7]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i8 (.Q(timer[8]), .C(CLK_c), .D(n133[8]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i9 (.Q(timer[9]), .C(CLK_c), .D(n133[9]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i10 (.Q(timer[10]), .C(CLK_c), .D(n133[10]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i11 (.Q(timer[11]), .C(CLK_c), .D(n133[11]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i12 (.Q(timer[12]), .C(CLK_c), .D(n133[12]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i13 (.Q(timer[13]), .C(CLK_c), .D(n133[13]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i14 (.Q(timer[14]), .C(CLK_c), .D(n133[14]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i15 (.Q(timer[15]), .C(CLK_c), .D(n133[15]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i16 (.Q(timer[16]), .C(CLK_c), .D(n133[16]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i17 (.Q(timer[17]), .C(CLK_c), .D(n133[17]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i18 (.Q(timer[18]), .C(CLK_c), .D(n133[18]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i19 (.Q(timer[19]), .C(CLK_c), .D(n133[19]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i20 (.Q(timer[20]), .C(CLK_c), .D(n133[20]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i21 (.Q(timer[21]), .C(CLK_c), .D(n133[21]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i22 (.Q(timer[22]), .C(CLK_c), .D(n133[22]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i23 (.Q(timer[23]), .C(CLK_c), .D(n133[23]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i24 (.Q(timer[24]), .C(CLK_c), .D(n133[24]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i25 (.Q(timer[25]), .C(CLK_c), .D(n133[25]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i26 (.Q(timer[26]), .C(CLK_c), .D(n133[26]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i27 (.Q(timer[27]), .C(CLK_c), .D(n133[27]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i28 (.Q(timer[28]), .C(CLK_c), .D(n133[28]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i29 (.Q(timer[29]), .C(CLK_c), .D(n133[29]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i30 (.Q(timer[30]), .C(CLK_c), .D(n133[30]));   // verilog/neopixel.v(12[12:21])
    SB_DFF timer_1546__i31 (.Q(timer[31]), .C(CLK_c), .D(n133[31]));   // verilog/neopixel.v(12[12:21])
    SB_DFFE state_i1 (.Q(\state[1] ), .C(CLK_c), .E(VCC_net), .D(n28194));   // verilog/neopixel.v(35[12] 117[6])
    SB_DFF \neo_pixel_transmitter.t0_i0_i0  (.Q(\neo_pixel_transmitter.t0 [0]), 
           .C(CLK_c), .D(n28188));   // verilog/neopixel.v(35[12] 117[6])
    SB_CARRY add_21_13 (.CI(n39054), .I0(bit_ctr[11]), .I1(GND_net), .CO(n39055));
    SB_LUT4 sub_14_add_2_13_lut (.I0(GND_net), .I1(timer[11]), .I2(n1[11]), 
            .I3(n39189), .O(one_wire_N_579[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_13 (.CI(n39189), .I0(timer[11]), .I1(n1[11]), 
            .CO(n39190));
    SB_LUT4 sub_14_add_2_12_lut (.I0(GND_net), .I1(timer[10]), .I2(n1[10]), 
            .I3(n39188), .O(one_wire_N_579[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR one_wire_108 (.Q(NEOPXL_c), .C(CLK_c), .E(n44987), .D(\neo_pixel_transmitter.done_N_642 ), 
            .R(n46810));   // verilog/neopixel.v(35[12] 117[6])
    SB_LUT4 add_21_12_lut (.I0(GND_net), .I1(bit_ctr[10]), .I2(GND_net), 
            .I3(n39053), .O(n255[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_12 (.CI(n39188), .I0(timer[10]), .I1(n1[10]), 
            .CO(n39189));
    SB_LUT4 sub_14_add_2_11_lut (.I0(GND_net), .I1(timer[9]), .I2(n1[9]), 
            .I3(n39187), .O(one_wire_N_579[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_11 (.CI(n39187), .I0(timer[9]), .I1(n1[9]), 
            .CO(n39188));
    SB_CARRY add_21_12 (.CI(n39053), .I0(bit_ctr[10]), .I1(GND_net), .CO(n39054));
    SB_LUT4 add_21_11_lut (.I0(GND_net), .I1(bit_ctr[9]), .I2(GND_net), 
            .I3(n39052), .O(n255[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_14_add_2_10_lut (.I0(GND_net), .I1(timer[8]), .I2(n1[8]), 
            .I3(n39186), .O(one_wire_N_579[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_11 (.CI(n39052), .I0(bit_ctr[9]), .I1(GND_net), .CO(n39053));
    SB_LUT4 add_21_10_lut (.I0(GND_net), .I1(bit_ctr[8]), .I2(GND_net), 
            .I3(n39051), .O(n255[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_10 (.CI(n39186), .I0(timer[8]), .I1(n1[8]), 
            .CO(n39187));
    SB_LUT4 sub_14_add_2_9_lut (.I0(GND_net), .I1(timer[7]), .I2(n1[7]), 
            .I3(n39185), .O(one_wire_N_579[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_14_add_2_9 (.CI(n39185), .I0(timer[7]), .I1(n1[7]), .CO(n39186));
    SB_CARRY add_21_10 (.CI(n39051), .I0(bit_ctr[8]), .I1(GND_net), .CO(n39052));
    SB_LUT4 sub_14_add_2_8_lut (.I0(GND_net), .I1(timer[6]), .I2(n1[6]), 
            .I3(n39184), .O(one_wire_N_579[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_14_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_21_9_lut (.I0(GND_net), .I1(bit_ctr[7]), .I2(GND_net), 
            .I3(n39050), .O(n255[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_21_9 (.CI(n39050), .I0(bit_ctr[7]), .I1(GND_net), .CO(n39051));
    SB_CARRY sub_14_add_2_8 (.CI(n39184), .I0(timer[6]), .I1(n1[6]), .CO(n39185));
    SB_LUT4 add_21_8_lut (.I0(GND_net), .I1(bit_ctr[6]), .I2(GND_net), 
            .I3(n39049), .O(n255[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_21_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mod_5_i606_3_lut_3_lut_4_lut_3_lut (.I0(bit_ctr[27]), .I1(n25166), 
            .I2(n27979), .I3(GND_net), .O(n28018));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i606_3_lut_3_lut_4_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 i35145_3_lut_4_lut_3_lut (.I0(bit_ctr[27]), .I1(n25166), .I2(n27979), 
            .I3(GND_net), .O(n27973));   // verilog/neopixel.v(22[26:36])
    defparam i35145_3_lut_4_lut_3_lut.LUT_INIT = 16'h1919;
    SB_LUT4 i1_2_lut_3_lut_3_lut (.I0(bit_ctr[27]), .I1(n25166), .I2(n27979), 
            .I3(GND_net), .O(n25164));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_3_lut_3_lut.LUT_INIT = 16'h8585;
    SB_LUT4 i1_4_lut_4_lut (.I0(bit_ctr[26]), .I1(n25164), .I2(n28018), 
            .I3(n27973), .O(n2));   // verilog/neopixel.v(22[26:36])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'h0007;
    SB_LUT4 i1_2_lut_3_lut (.I0(n34629), .I1(\neo_pixel_transmitter.done ), 
            .I2(start), .I3(GND_net), .O(n44777));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 i35017_2_lut_3_lut (.I0(n34525), .I1(\neo_pixel_transmitter.done ), 
            .I2(\state[0] ), .I3(GND_net), .O(n49782));   // verilog/neopixel.v(35[12] 117[6])
    defparam i35017_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i2_2_lut_3_lut_adj_1622 (.I0(n26525), .I1(one_wire_N_579[2]), 
            .I2(one_wire_N_579[3]), .I3(GND_net), .O(n34429));
    defparam i2_2_lut_3_lut_adj_1622.LUT_INIT = 16'hfefe;
    SB_LUT4 mod_5_i1689_3_lut (.I0(n2403), .I1(n2456[18]), .I2(n2423), 
            .I3(GND_net), .O(n2502));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1689_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1688_3_lut (.I0(n2402), .I1(n2456[19]), .I2(n2423), 
            .I3(GND_net), .O(n2501));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1688_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1690_3_lut (.I0(n2404), .I1(n2456[17]), .I2(n2423), 
            .I3(GND_net), .O(n2503));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1690_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1695_3_lut (.I0(n2409), .I1(n2456[12]), .I2(n2423), 
            .I3(GND_net), .O(n2508));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1687_3_lut (.I0(n2401), .I1(n2456[20]), .I2(n2423), 
            .I3(GND_net), .O(n2500));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(LED_c), 
            .I3(\state_3__N_428[1] ), .O(n28088));   // verilog/neopixel.v(35[12] 117[6])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i17555_3_lut_4_lut (.I0(bit_ctr[29]), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[28]), .O(n27979));   // verilog/neopixel.v(18[12:19])
    defparam i17555_3_lut_4_lut.LUT_INIT = 16'hdb6d;
    SB_LUT4 mod_5_i1686_3_lut (.I0(n2400), .I1(n2456[21]), .I2(n2423), 
            .I3(GND_net), .O(n2499));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1686_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17557_3_lut_4_lut (.I0(bit_ctr[29]), .I1(bit_ctr[30]), .I2(bit_ctr[31]), 
            .I3(bit_ctr[28]), .O(n25166));   // verilog/neopixel.v(18[12:19])
    defparam i17557_3_lut_4_lut.LUT_INIT = 16'hb6db;
    SB_LUT4 mod_5_i1691_3_lut (.I0(n2405), .I1(n2456[16]), .I2(n2423), 
            .I3(GND_net), .O(n2504));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1694_3_lut (.I0(n2408), .I1(n2456[13]), .I2(n2423), 
            .I3(GND_net), .O(n2507));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1694_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1692_3_lut (.I0(n2406), .I1(n2456[15]), .I2(n2423), 
            .I3(GND_net), .O(n2505));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1692_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1681_3_lut (.I0(n2395), .I1(n2456[26]), .I2(n2423), 
            .I3(GND_net), .O(n2494));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1681_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1679_3_lut (.I0(n2393), .I1(n2456[28]), .I2(n2423), 
            .I3(GND_net), .O(n2492));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1679_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1680_3_lut (.I0(n2394), .I1(n2456[27]), .I2(n2423), 
            .I3(GND_net), .O(n2493));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1680_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1678_3_lut (.I0(n2392), .I1(n2456[29]), .I2(n2423), 
            .I3(GND_net), .O(n2491));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1678_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1685_3_lut (.I0(n2399), .I1(n2456[22]), .I2(n2423), 
            .I3(GND_net), .O(n2498));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1683_3_lut (.I0(n2397), .I1(n2456[24]), .I2(n2423), 
            .I3(GND_net), .O(n2496));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1683_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1684_3_lut (.I0(n2398), .I1(n2456[23]), .I2(n2423), 
            .I3(GND_net), .O(n2497));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1684_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1682_3_lut (.I0(n2396), .I1(n2456[25]), .I2(n2423), 
            .I3(GND_net), .O(n2495));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1682_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1677_3_lut (.I0(n2391), .I1(n2456[30]), .I2(n2423), 
            .I3(GND_net), .O(n2490));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1677_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1696_3_lut (.I0(bit_ctr[11]), .I1(n2456[11]), .I2(n2423), 
            .I3(GND_net), .O(n2509));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1696_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i9_3_lut (.I0(bit_ctr[4]), .I1(n3103), .I2(n3109), .I3(GND_net), 
            .O(n36_adj_4837));   // verilog/neopixel.v(22[26:36])
    defparam i9_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 mod_5_i1693_3_lut (.I0(n2407), .I1(n2456[14]), .I2(n2423), 
            .I3(GND_net), .O(n2506));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1693_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i19_4_lut_adj_1623 (.I0(n3105), .I1(n3099), .I2(n3108), .I3(n3107), 
            .O(n46_adj_4838));   // verilog/neopixel.v(22[26:36])
    defparam i19_4_lut_adj_1623.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1624 (.I0(n3085), .I1(n3087), .I2(n3086), .I3(n3088), 
            .O(n42_adj_4839));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1624.LUT_INIT = 16'hfffe;
    SB_LUT4 i5_2_lut (.I0(n3091), .I1(n3092), .I2(GND_net), .I3(GND_net), 
            .O(n32_adj_4840));   // verilog/neopixel.v(22[26:36])
    defparam i5_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1625 (.I0(n2490), .I1(n2489), .I2(GND_net), .I3(GND_net), 
            .O(n22_adj_4841));   // verilog/neopixel.v(22[26:36])
    defparam i1_2_lut_adj_1625.LUT_INIT = 16'heeee;
    SB_LUT4 i7_3_lut_adj_1626 (.I0(bit_ctr[10]), .I1(n2506), .I2(n2509), 
            .I3(GND_net), .O(n28_adj_4842));   // verilog/neopixel.v(22[26:36])
    defparam i7_3_lut_adj_1626.LUT_INIT = 16'hecec;
    SB_LUT4 i17_4_lut_adj_1627 (.I0(n3093), .I1(n3095), .I2(n3094), .I3(n3097), 
            .O(n44_adj_4843));   // verilog/neopixel.v(22[26:36])
    defparam i17_4_lut_adj_1627.LUT_INIT = 16'hfffe;
    SB_LUT4 i23_4_lut (.I0(n3096), .I1(n46_adj_4838), .I2(n36_adj_4837), 
            .I3(n3101), .O(n50));   // verilog/neopixel.v(22[26:36])
    defparam i23_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1628 (.I0(n2508), .I1(n2503), .I2(n2501), .I3(n2502), 
            .O(n36_adj_4844));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1628.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1629 (.I0(n2495), .I1(n2497), .I2(n2496), .I3(n2498), 
            .O(n34_adj_4845));   // verilog/neopixel.v(22[26:36])
    defparam i13_4_lut_adj_1629.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1630 (.I0(n2491), .I1(n2493), .I2(n2492), .I3(n2494), 
            .O(n33_adj_4846));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1630.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1631 (.I0(n3104), .I1(n42_adj_4839), .I2(n3084), 
            .I3(n3083), .O(n48_adj_4847));   // verilog/neopixel.v(22[26:36])
    defparam i21_4_lut_adj_1631.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1632 (.I0(n3089), .I1(n44_adj_4843), .I2(n32_adj_4840), 
            .I3(n3090), .O(n49_adj_4848));   // verilog/neopixel.v(22[26:36])
    defparam i22_4_lut_adj_1632.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1633 (.I0(n2505), .I1(n2507), .I2(n2504), .I3(n22_adj_4841), 
            .O(n37_adj_4849));   // verilog/neopixel.v(22[26:36])
    defparam i16_4_lut_adj_1633.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1634 (.I0(n2499), .I1(n36_adj_4844), .I2(n28_adj_4842), 
            .I3(n2500), .O(n39_adj_4850));   // verilog/neopixel.v(22[26:36])
    defparam i18_4_lut_adj_1634.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1635 (.I0(n3098), .I1(n3102), .I2(n3106), .I3(n3100), 
            .O(n47_adj_4851));   // verilog/neopixel.v(22[26:36])
    defparam i20_4_lut_adj_1635.LUT_INIT = 16'hfffe;
    SB_LUT4 i26_4_lut_adj_1636 (.I0(n47_adj_4851), .I1(n49_adj_4848), .I2(n48_adj_4847), 
            .I3(n50), .O(n3116));   // verilog/neopixel.v(22[26:36])
    defparam i26_4_lut_adj_1636.LUT_INIT = 16'hfffe;
    SB_LUT4 i20_4_lut_adj_1637 (.I0(n39_adj_4850), .I1(n37_adj_4849), .I2(n33_adj_4846), 
            .I3(n34_adj_4845), .O(n2522));   // verilog/neopixel.v(22[26:36])
    defparam i20_4_lut_adj_1637.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1968_3_lut (.I0(bit_ctr[7]), .I1(n2852[7]), .I2(n2819), 
            .I3(GND_net), .O(n2909));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1968_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1967_3_lut (.I0(n2809), .I1(n2852[8]), .I2(n2819), 
            .I3(GND_net), .O(n2908));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1967_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_inv_0_i4_1_lut (.I0(\neo_pixel_transmitter.t0 [3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[3]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i1966_3_lut (.I0(n2808), .I1(n2852[9]), .I2(n2819), 
            .I3(GND_net), .O(n2907));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1966_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1965_3_lut (.I0(n2807), .I1(n2852[10]), .I2(n2819), 
            .I3(GND_net), .O(n2906));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1965_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1964_3_lut (.I0(n2806), .I1(n2852[11]), .I2(n2819), 
            .I3(GND_net), .O(n2905));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1963_3_lut (.I0(n2805), .I1(n2852[12]), .I2(n2819), 
            .I3(GND_net), .O(n2904));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1963_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1962_3_lut (.I0(n2804), .I1(n2852[13]), .I2(n2819), 
            .I3(GND_net), .O(n2903));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1961_3_lut (.I0(n2803), .I1(n2852[14]), .I2(n2819), 
            .I3(GND_net), .O(n2902));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i36454_1_lut (.I0(n3017), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51407));
    defparam i36454_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i1960_3_lut (.I0(n2802), .I1(n2852[15]), .I2(n2819), 
            .I3(GND_net), .O(n2901));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1960_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1959_3_lut (.I0(n2801), .I1(n2852[16]), .I2(n2819), 
            .I3(GND_net), .O(n2900));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1959_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1958_3_lut (.I0(n2800), .I1(n2852[17]), .I2(n2819), 
            .I3(GND_net), .O(n2899));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1958_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1957_3_lut (.I0(n2799), .I1(n2852[18]), .I2(n2819), 
            .I3(GND_net), .O(n2898));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1957_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1956_3_lut (.I0(n2798), .I1(n2852[19]), .I2(n2819), 
            .I3(GND_net), .O(n2897));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1956_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1955_3_lut (.I0(n2797), .I1(n2852[20]), .I2(n2819), 
            .I3(GND_net), .O(n2896));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1955_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1954_3_lut (.I0(n2796), .I1(n2852[21]), .I2(n2819), 
            .I3(GND_net), .O(n2895));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1954_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1953_3_lut (.I0(n2795), .I1(n2852[22]), .I2(n2819), 
            .I3(GND_net), .O(n2894));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1953_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1952_3_lut (.I0(n2794), .I1(n2852[23]), .I2(n2819), 
            .I3(GND_net), .O(n2893));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1952_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_inv_0_i5_1_lut (.I0(\neo_pixel_transmitter.t0 [4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[4]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i1951_3_lut (.I0(n2793), .I1(n2852[24]), .I2(n2819), 
            .I3(GND_net), .O(n2892));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1951_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1950_3_lut (.I0(n2792), .I1(n2852[25]), .I2(n2819), 
            .I3(GND_net), .O(n2891));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1950_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1949_3_lut (.I0(n2791), .I1(n2852[26]), .I2(n2819), 
            .I3(GND_net), .O(n2890));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1949_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 sub_14_inv_0_i6_1_lut (.I0(\neo_pixel_transmitter.t0 [5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[5]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mod_5_i1948_3_lut (.I0(n2790), .I1(n2852[27]), .I2(n2819), 
            .I3(GND_net), .O(n2889));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1948_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1619_3_lut (.I0(n2301), .I1(n2357[21]), .I2(n2324), 
            .I3(GND_net), .O(n2400));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1619_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1616_3_lut (.I0(n2298), .I1(n2357[24]), .I2(n2324), 
            .I3(GND_net), .O(n2397));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1616_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1624_3_lut (.I0(n2306), .I1(n2357[16]), .I2(n2324), 
            .I3(GND_net), .O(n2405));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1624_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1617_3_lut (.I0(n2299), .I1(n2357[23]), .I2(n2324), 
            .I3(GND_net), .O(n2398));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1617_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1625_3_lut (.I0(n2307), .I1(n2357[15]), .I2(n2324), 
            .I3(GND_net), .O(n2406));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1625_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1622_3_lut (.I0(n2304), .I1(n2357[18]), .I2(n2324), 
            .I3(GND_net), .O(n2403));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1622_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1612_3_lut (.I0(n2294), .I1(n2357[28]), .I2(n2324), 
            .I3(GND_net), .O(n2393));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1612_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1611_3_lut (.I0(n2293), .I1(n2357[29]), .I2(n2324), 
            .I3(GND_net), .O(n2392));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1611_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1610_3_lut (.I0(n2292), .I1(n2357[30]), .I2(n2324), 
            .I3(GND_net), .O(n2391));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1610_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1626_3_lut (.I0(n2308), .I1(n2357[14]), .I2(n2324), 
            .I3(GND_net), .O(n2407));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1626_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1627_3_lut (.I0(n2309), .I1(n2357[13]), .I2(n2324), 
            .I3(GND_net), .O(n2408));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1627_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1614_3_lut (.I0(n2296), .I1(n2357[26]), .I2(n2324), 
            .I3(GND_net), .O(n2395));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1614_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1613_3_lut (.I0(n2295), .I1(n2357[27]), .I2(n2324), 
            .I3(GND_net), .O(n2394));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1613_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1615_3_lut (.I0(n2297), .I1(n2357[25]), .I2(n2324), 
            .I3(GND_net), .O(n2396));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1615_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1623_3_lut (.I0(n2305), .I1(n2357[17]), .I2(n2324), 
            .I3(GND_net), .O(n2404));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1623_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1618_3_lut (.I0(n2300), .I1(n2357[22]), .I2(n2324), 
            .I3(GND_net), .O(n2399));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1618_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1620_3_lut (.I0(n2302), .I1(n2357[20]), .I2(n2324), 
            .I3(GND_net), .O(n2401));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1620_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1628_3_lut (.I0(bit_ctr[12]), .I1(n2357[12]), .I2(n2324), 
            .I3(GND_net), .O(n2409));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1628_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1621_3_lut (.I0(n2303), .I1(n2357[19]), .I2(n2324), 
            .I3(GND_net), .O(n2402));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1621_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i6_3_lut_adj_1638 (.I0(n2402), .I1(bit_ctr[11]), .I2(n2409), 
            .I3(GND_net), .O(n26_adj_4852));   // verilog/neopixel.v(22[26:36])
    defparam i6_3_lut_adj_1638.LUT_INIT = 16'heaea;
    SB_LUT4 i14_4_lut_adj_1639 (.I0(n2401), .I1(n2399), .I2(n2404), .I3(n2396), 
            .O(n34_adj_4853));   // verilog/neopixel.v(22[26:36])
    defparam i14_4_lut_adj_1639.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1640 (.I0(n2394), .I1(n2395), .I2(n2408), .I3(n2407), 
            .O(n32_adj_4854));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1640.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut_adj_1641 (.I0(n2391), .I1(n2392), .I2(n2390), .I3(n2393), 
            .O(n31_adj_4855));   // verilog/neopixel.v(22[26:36])
    defparam i11_4_lut_adj_1641.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1642 (.I0(n2403), .I1(n2406), .I2(n2398), .I3(n2405), 
            .O(n35_adj_4856));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1642.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1643 (.I0(n2397), .I1(n34_adj_4853), .I2(n26_adj_4852), 
            .I3(n2400), .O(n37_adj_4857));   // verilog/neopixel.v(22[26:36])
    defparam i17_4_lut_adj_1643.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1644 (.I0(n37_adj_4857), .I1(n35_adj_4856), .I2(n31_adj_4855), 
            .I3(n32_adj_4854), .O(n2423));   // verilog/neopixel.v(22[26:36])
    defparam i19_4_lut_adj_1644.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i2033_3_lut (.I0(n2907), .I1(n2951[9]), .I2(n2918), 
            .I3(GND_net), .O(n3006));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2015_3_lut (.I0(n2889), .I1(n2951[27]), .I2(n2918), 
            .I3(GND_net), .O(n2988));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2018_3_lut (.I0(n2892), .I1(n2951[24]), .I2(n2918), 
            .I3(GND_net), .O(n2991));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2018_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2013_3_lut (.I0(n2887), .I1(n2951[29]), .I2(n2918), 
            .I3(GND_net), .O(n2986));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2013_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i17538_3_lut (.I0(bit_ctr[6]), .I1(n2951[6]), .I2(n2918), 
            .I3(GND_net), .O(n30593));
    defparam i17538_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2030_3_lut (.I0(n2904), .I1(n2951[12]), .I2(n2918), 
            .I3(GND_net), .O(n3003));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2024_3_lut (.I0(n2898), .I1(n2951[18]), .I2(n2918), 
            .I3(GND_net), .O(n2997));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2029_3_lut (.I0(n2903), .I1(n2951[13]), .I2(n2918), 
            .I3(GND_net), .O(n3002));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2029_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2012_3_lut (.I0(n2886), .I1(n2951[30]), .I2(n2918), 
            .I3(GND_net), .O(n2985));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2012_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2023_3_lut (.I0(n2897), .I1(n2951[19]), .I2(n2918), 
            .I3(GND_net), .O(n2996));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2023_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2031_3_lut (.I0(n2905), .I1(n2951[11]), .I2(n2918), 
            .I3(GND_net), .O(n3004));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2020_3_lut (.I0(n2894), .I1(n2951[22]), .I2(n2918), 
            .I3(GND_net), .O(n2993));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2020_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2022_3_lut (.I0(n2896), .I1(n2951[20]), .I2(n2918), 
            .I3(GND_net), .O(n2995));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2017_3_lut (.I0(n2891), .I1(n2951[25]), .I2(n2918), 
            .I3(GND_net), .O(n2990));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2017_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2016_3_lut (.I0(n2890), .I1(n2951[26]), .I2(n2918), 
            .I3(GND_net), .O(n2989));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2021_3_lut (.I0(n2895), .I1(n2951[21]), .I2(n2918), 
            .I3(GND_net), .O(n2994));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2014_3_lut (.I0(n2888), .I1(n2951[28]), .I2(n2918), 
            .I3(GND_net), .O(n2987));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2014_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2027_3_lut (.I0(n2901), .I1(n2951[15]), .I2(n2918), 
            .I3(GND_net), .O(n3000));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2019_3_lut (.I0(n2893), .I1(n2951[23]), .I2(n2918), 
            .I3(GND_net), .O(n2992));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2035_3_lut (.I0(n2909), .I1(n2951[7]), .I2(n2918), 
            .I3(GND_net), .O(n3008));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2035_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2034_3_lut (.I0(n2908), .I1(n2951[8]), .I2(n2918), 
            .I3(GND_net), .O(n3007));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2026_3_lut (.I0(n2900), .I1(n2951[16]), .I2(n2918), 
            .I3(GND_net), .O(n2999));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2026_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1945_3_lut (.I0(n2787), .I1(n2852[30]), .I2(n2819), 
            .I3(GND_net), .O(n2886));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1945_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i7_3_lut_adj_1645 (.I0(bit_ctr[6]), .I1(n2897), .I2(n2909), 
            .I3(GND_net), .O(n32_adj_4858));   // verilog/neopixel.v(22[26:36])
    defparam i7_3_lut_adj_1645.LUT_INIT = 16'hecec;
    SB_LUT4 i17_4_lut_adj_1646 (.I0(n2906), .I1(n2901), .I2(n2899), .I3(n2905), 
            .O(n42_adj_4859));   // verilog/neopixel.v(22[26:36])
    defparam i17_4_lut_adj_1646.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut (.I0(n2903), .I1(n2886), .I2(n2885), .I3(GND_net), 
            .O(n38_adj_4860));   // verilog/neopixel.v(22[26:36])
    defparam i13_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i18_4_lut_adj_1647 (.I0(n2904), .I1(n2900), .I2(n2907), .I3(n2898), 
            .O(n43_adj_4861));   // verilog/neopixel.v(22[26:36])
    defparam i18_4_lut_adj_1647.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1648 (.I0(n2891), .I1(n2893), .I2(n2892), .I3(n2894), 
            .O(n40_adj_4862));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1648.LUT_INIT = 16'hfffe;
    SB_LUT4 i21_4_lut_adj_1649 (.I0(n2895), .I1(n42_adj_4859), .I2(n32_adj_4858), 
            .I3(n2896), .O(n46_adj_4863));   // verilog/neopixel.v(22[26:36])
    defparam i21_4_lut_adj_1649.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1650 (.I0(n2887), .I1(n2889), .I2(n2888), .I3(n2890), 
            .O(n39_adj_4864));   // verilog/neopixel.v(22[26:36])
    defparam i14_4_lut_adj_1650.LUT_INIT = 16'hfffe;
    SB_LUT4 i22_4_lut_adj_1651 (.I0(n43_adj_4861), .I1(n2902), .I2(n38_adj_4860), 
            .I3(n2908), .O(n47_adj_4865));   // verilog/neopixel.v(22[26:36])
    defparam i22_4_lut_adj_1651.LUT_INIT = 16'hfffe;
    SB_LUT4 i24_4_lut (.I0(n47_adj_4865), .I1(n39_adj_4864), .I2(n46_adj_4863), 
            .I3(n40_adj_4862), .O(n2918));   // verilog/neopixel.v(22[26:36])
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i2028_3_lut (.I0(n2902), .I1(n2951[14]), .I2(n2918), 
            .I3(GND_net), .O(n3001));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2032_3_lut (.I0(n2906), .I1(n2951[10]), .I2(n2918), 
            .I3(GND_net), .O(n3005));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2032_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i2025_3_lut (.I0(n2899), .I1(n2951[17]), .I2(n2918), 
            .I3(GND_net), .O(n2998));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i2025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i18_4_lut_adj_1652 (.I0(n2984), .I1(n2998), .I2(n3005), .I3(n3001), 
            .O(n44_adj_4866));
    defparam i18_4_lut_adj_1652.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1653 (.I0(n2999), .I1(n3007), .I2(n3008), .I3(n2992), 
            .O(n42_adj_4867));
    defparam i16_4_lut_adj_1653.LUT_INIT = 16'hfffe;
    SB_LUT4 i17_4_lut_adj_1654 (.I0(n2990), .I1(n2995), .I2(n2993), .I3(n3004), 
            .O(n43_adj_4868));
    defparam i17_4_lut_adj_1654.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1655 (.I0(n3000), .I1(n2987), .I2(n2994), .I3(n2989), 
            .O(n41_adj_4869));
    defparam i15_4_lut_adj_1655.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1656 (.I0(n2996), .I1(n2985), .I2(n3002), .I3(n2997), 
            .O(n40_adj_4870));
    defparam i14_4_lut_adj_1656.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_3_lut_adj_1657 (.I0(n3003), .I1(bit_ctr[5]), .I2(n30593), 
            .I3(GND_net), .O(n39_adj_4871));
    defparam i13_3_lut_adj_1657.LUT_INIT = 16'heaea;
    SB_LUT4 i24_4_lut_adj_1658 (.I0(n41_adj_4869), .I1(n43_adj_4868), .I2(n42_adj_4867), 
            .I3(n44_adj_4866), .O(n50_adj_4872));
    defparam i24_4_lut_adj_1658.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut_adj_1659 (.I0(n2986), .I1(n2991), .I2(n2988), .I3(n3006), 
            .O(n45_adj_4873));
    defparam i19_4_lut_adj_1659.LUT_INIT = 16'hfffe;
    SB_LUT4 i25_4_lut (.I0(n45_adj_4873), .I1(n50_adj_4872), .I2(n39_adj_4871), 
            .I3(n40_adj_4870), .O(n3017));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1549_3_lut (.I0(n2199), .I1(n2258[24]), .I2(n2225), 
            .I3(GND_net), .O(n2298));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1549_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1547_3_lut (.I0(n2197), .I1(n2258[26]), .I2(n2225), 
            .I3(GND_net), .O(n2296));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1547_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1551_3_lut (.I0(n2201), .I1(n2258[22]), .I2(n2225), 
            .I3(GND_net), .O(n2300));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1551_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1550_3_lut (.I0(n2200), .I1(n2258[23]), .I2(n2225), 
            .I3(GND_net), .O(n2299));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1550_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1556_3_lut (.I0(n2206), .I1(n2258[17]), .I2(n2225), 
            .I3(GND_net), .O(n2305));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1556_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1554_3_lut (.I0(n2204), .I1(n2258[19]), .I2(n2225), 
            .I3(GND_net), .O(n2303));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1554_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1559_3_lut (.I0(n2209), .I1(n2258[14]), .I2(n2225), 
            .I3(GND_net), .O(n2308));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1559_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1558_3_lut (.I0(n2208), .I1(n2258[15]), .I2(n2225), 
            .I3(GND_net), .O(n2307));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1558_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1553_3_lut (.I0(n2203), .I1(n2258[20]), .I2(n2225), 
            .I3(GND_net), .O(n2302));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1553_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1557_3_lut (.I0(n2207), .I1(n2258[16]), .I2(n2225), 
            .I3(GND_net), .O(n2306));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1557_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1552_3_lut (.I0(n2202), .I1(n2258[21]), .I2(n2225), 
            .I3(GND_net), .O(n2301));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1552_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1543_3_lut (.I0(n2193), .I1(n2258[30]), .I2(n2225), 
            .I3(GND_net), .O(n2292));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1555_3_lut (.I0(n2205), .I1(n2258[18]), .I2(n2225), 
            .I3(GND_net), .O(n2304));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1555_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1546_3_lut (.I0(n2196), .I1(n2258[27]), .I2(n2225), 
            .I3(GND_net), .O(n2295));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1546_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1548_3_lut (.I0(n2198), .I1(n2258[25]), .I2(n2225), 
            .I3(GND_net), .O(n2297));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1544_3_lut (.I0(n2194), .I1(n2258[29]), .I2(n2225), 
            .I3(GND_net), .O(n2293));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1544_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1545_3_lut (.I0(n2195), .I1(n2258[28]), .I2(n2225), 
            .I3(GND_net), .O(n2294));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1545_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1560_3_lut (.I0(bit_ctr[13]), .I1(n2258[13]), .I2(n2225), 
            .I3(GND_net), .O(n2309));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1560_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i11_4_lut_adj_1660 (.I0(n2294), .I1(n2293), .I2(n2297), .I3(n2295), 
            .O(n30_adj_4874));   // verilog/neopixel.v(22[26:36])
    defparam i11_4_lut_adj_1660.LUT_INIT = 16'hfffe;
    SB_LUT4 i21432_2_lut (.I0(bit_ctr[12]), .I1(n2309), .I2(GND_net), 
            .I3(GND_net), .O(n34495));
    defparam i21432_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i15_4_lut_adj_1661 (.I0(n2304), .I1(n30_adj_4874), .I2(n2292), 
            .I3(n2291), .O(n34_adj_4875));   // verilog/neopixel.v(22[26:36])
    defparam i15_4_lut_adj_1661.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1662 (.I0(n2301), .I1(n2306), .I2(n34495), .I3(n2302), 
            .O(n32_adj_4876));   // verilog/neopixel.v(22[26:36])
    defparam i13_4_lut_adj_1662.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_1663 (.I0(n2307), .I1(n2308), .I2(n2303), .I3(n2305), 
            .O(n33_adj_4877));   // verilog/neopixel.v(22[26:36])
    defparam i14_4_lut_adj_1663.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut_adj_1664 (.I0(n2299), .I1(n2300), .I2(n2296), .I3(n2298), 
            .O(n31_adj_4878));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1664.LUT_INIT = 16'hfffe;
    SB_LUT4 i18_4_lut_adj_1665 (.I0(n31_adj_4878), .I1(n33_adj_4877), .I2(n32_adj_4876), 
            .I3(n34_adj_4875), .O(n2324));   // verilog/neopixel.v(22[26:36])
    defparam i18_4_lut_adj_1665.LUT_INIT = 16'hfffe;
    SB_LUT4 i36453_1_lut (.I0(n1235), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51406));
    defparam i36453_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i23_4_lut_adj_1666 (.I0(n41_adj_4820), .I1(n43_adj_4819), .I2(n42_adj_4818), 
            .I3(n44_adj_4817), .O(n2819));   // verilog/neopixel.v(22[26:36])
    defparam i23_4_lut_adj_1666.LUT_INIT = 16'hfffe;
    SB_LUT4 mod_5_i1479_3_lut (.I0(n2097), .I1(n2159[27]), .I2(n2126), 
            .I3(GND_net), .O(n2196));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1479_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1481_3_lut (.I0(n2099), .I1(n2159[25]), .I2(n2126), 
            .I3(GND_net), .O(n2198));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1481_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1488_3_lut (.I0(n2106), .I1(n2159[18]), .I2(n2126), 
            .I3(GND_net), .O(n2205));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1488_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1485_3_lut (.I0(n2103), .I1(n2159[21]), .I2(n2126), 
            .I3(GND_net), .O(n2202));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1485_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1484_3_lut (.I0(n2102), .I1(n2159[22]), .I2(n2126), 
            .I3(GND_net), .O(n2201));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1484_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1482_3_lut (.I0(n2100), .I1(n2159[24]), .I2(n2126), 
            .I3(GND_net), .O(n2199));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1482_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1486_3_lut (.I0(n2104), .I1(n2159[20]), .I2(n2126), 
            .I3(GND_net), .O(n2203));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1486_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1490_3_lut (.I0(n2108), .I1(n2159[16]), .I2(n2126), 
            .I3(GND_net), .O(n2207));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1490_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1492_3_lut (.I0(bit_ctr[14]), .I1(n2159[14]), .I2(n2126), 
            .I3(GND_net), .O(n2209));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1492_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1489_3_lut (.I0(n2107), .I1(n2159[17]), .I2(n2126), 
            .I3(GND_net), .O(n2206));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1489_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1483_3_lut (.I0(n2101), .I1(n2159[23]), .I2(n2126), 
            .I3(GND_net), .O(n2200));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1483_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1491_3_lut (.I0(n2109), .I1(n2159[15]), .I2(n2126), 
            .I3(GND_net), .O(n2208));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1491_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1480_3_lut (.I0(n2098), .I1(n2159[26]), .I2(n2126), 
            .I3(GND_net), .O(n2197));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1480_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1487_3_lut (.I0(n2105), .I1(n2159[19]), .I2(n2126), 
            .I3(GND_net), .O(n2204));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1487_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1478_3_lut (.I0(n2096), .I1(n2159[28]), .I2(n2126), 
            .I3(GND_net), .O(n2195));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1478_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1477_3_lut (.I0(n2095), .I1(n2159[29]), .I2(n2126), 
            .I3(GND_net), .O(n2194));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1477_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mod_5_i1476_3_lut (.I0(n2094), .I1(n2159[30]), .I2(n2126), 
            .I3(GND_net), .O(n2193));   // verilog/neopixel.v(22[26:36])
    defparam mod_5_i1476_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i10_4_lut_adj_1667 (.I0(n2193), .I1(n2194), .I2(n2192), .I3(n2195), 
            .O(n28_adj_4879));   // verilog/neopixel.v(22[26:36])
    defparam i10_4_lut_adj_1667.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_4_lut_adj_1668 (.I0(n2204), .I1(n2197), .I2(n2208), .I3(n2200), 
            .O(n31_adj_4880));   // verilog/neopixel.v(22[26:36])
    defparam i13_4_lut_adj_1668.LUT_INIT = 16'hfffe;
    SB_LUT4 i4_3_lut_adj_1669 (.I0(bit_ctr[13]), .I1(n2206), .I2(n2209), 
            .I3(GND_net), .O(n22_adj_4881));   // verilog/neopixel.v(22[26:36])
    defparam i4_3_lut_adj_1669.LUT_INIT = 16'hecec;
    SB_LUT4 i12_4_lut_adj_1670 (.I0(n2207), .I1(n2203), .I2(n2199), .I3(n2201), 
            .O(n30_adj_4882));   // verilog/neopixel.v(22[26:36])
    defparam i12_4_lut_adj_1670.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_1671 (.I0(n31_adj_4880), .I1(n2202), .I2(n28_adj_4879), 
            .I3(n2205), .O(n34_adj_4883));   // verilog/neopixel.v(22[26:36])
    defparam i16_4_lut_adj_1671.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_2_lut_adj_1672 (.I0(n2198), .I1(n2196), .I2(GND_net), .I3(GND_net), 
            .O(n21_adj_4884));   // verilog/neopixel.v(22[26:36])
    defparam i3_2_lut_adj_1672.LUT_INIT = 16'heeee;
    SB_LUT4 i17_4_lut_adj_1673 (.I0(n21_adj_4884), .I1(n34_adj_4883), .I2(n30_adj_4882), 
            .I3(n22_adj_4881), .O(n2225));   // verilog/neopixel.v(22[26:36])
    defparam i17_4_lut_adj_1673.LUT_INIT = 16'hfffe;
    SB_LUT4 i35309_3_lut_4_lut (.I0(n26525), .I1(n50261), .I2(start), 
            .I3(\state[1] ), .O(n50262));
    defparam i35309_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i34962_2_lut_3_lut (.I0(one_wire_N_579[2]), .I1(one_wire_N_579[3]), 
            .I2(start), .I3(GND_net), .O(n49769));
    defparam i34962_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i3_4_lut_4_lut (.I0(n34525), .I1(\state[1] ), .I2(\state[0] ), 
            .I3(\neo_pixel_transmitter.done ), .O(n46810));
    defparam i3_4_lut_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 sub_14_inv_0_i7_1_lut (.I0(\neo_pixel_transmitter.t0 [6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[6]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 sub_14_inv_0_i8_1_lut (.I0(\neo_pixel_transmitter.t0 [7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1[7]));   // verilog/neopixel.v(53[15:25])
    defparam sub_14_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1,500000)_U0 
//

module \quadrature_decoder(1,500000)_U0  (b_prev, GND_net, a_new, direction_N_3807, 
            ENCODER0_B_N_keep, n1188, ENCODER0_A_N_keep, encoder0_position, 
            VCC_net, n28241, n1152) /* synthesis lattice_noprune=1 */ ;
    output b_prev;
    input GND_net;
    output [1:0]a_new;
    output direction_N_3807;
    input ENCODER0_B_N_keep;
    input n1188;
    input ENCODER0_A_N_keep;
    output [31:0]encoder0_position;
    input VCC_net;
    input n28241;
    output n1152;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(41[9:14])
    
    wire direction_N_3810, debounce_cnt, a_prev;
    wire [1:0]a_new_c;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [31:0]n133;
    
    wire direction_N_3806, n40498, n40497, n40496, n40495, n40494, 
        n40493, n40492, n40491, n40490, n40489, n40488, n40487, 
        n40486, n40485, n40484, n40483, n40482, a_prev_N_3813, n40481, 
        n40480, n40479, n40478, n40477, n40476, n40475, n40474, 
        n40473, n40472, n40471, n40470, n40469, n40468, n28243, 
        n28242;
    
    SB_LUT4 b_prev_I_0_65_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3810));   // vhdl/quadrature_decoder.vhd(80[37:56])
    defparam b_prev_I_0_65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(direction_N_3810), 
            .I3(a_new[1]), .O(direction_N_3807));   // vhdl/quadrature_decoder.vhd(79[10] 80[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1188), .D(ENCODER0_B_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i0 (.Q(a_new_c[0]), .C(n1188), .D(ENCODER0_A_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 position_1553_add_4_33_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[31]), .I3(n40498), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_1553_add_4_32_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[30]), .I3(n40497), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_32 (.CI(n40497), .I0(direction_N_3806), 
            .I1(encoder0_position[30]), .CO(n40498));
    SB_LUT4 position_1553_add_4_31_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[29]), .I3(n40496), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_31 (.CI(n40496), .I0(direction_N_3806), 
            .I1(encoder0_position[29]), .CO(n40497));
    SB_LUT4 position_1553_add_4_30_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[28]), .I3(n40495), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_30 (.CI(n40495), .I0(direction_N_3806), 
            .I1(encoder0_position[28]), .CO(n40496));
    SB_LUT4 position_1553_add_4_29_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[27]), .I3(n40494), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_29 (.CI(n40494), .I0(direction_N_3806), 
            .I1(encoder0_position[27]), .CO(n40495));
    SB_LUT4 position_1553_add_4_28_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[26]), .I3(n40493), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_28 (.CI(n40493), .I0(direction_N_3806), 
            .I1(encoder0_position[26]), .CO(n40494));
    SB_LUT4 position_1553_add_4_27_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[25]), .I3(n40492), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_27 (.CI(n40492), .I0(direction_N_3806), 
            .I1(encoder0_position[25]), .CO(n40493));
    SB_LUT4 position_1553_add_4_26_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[24]), .I3(n40491), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_26 (.CI(n40491), .I0(direction_N_3806), 
            .I1(encoder0_position[24]), .CO(n40492));
    SB_LUT4 position_1553_add_4_25_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[23]), .I3(n40490), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_25 (.CI(n40490), .I0(direction_N_3806), 
            .I1(encoder0_position[23]), .CO(n40491));
    SB_LUT4 position_1553_add_4_24_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[22]), .I3(n40489), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_24 (.CI(n40489), .I0(direction_N_3806), 
            .I1(encoder0_position[22]), .CO(n40490));
    SB_LUT4 position_1553_add_4_23_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[21]), .I3(n40488), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_23 (.CI(n40488), .I0(direction_N_3806), 
            .I1(encoder0_position[21]), .CO(n40489));
    SB_LUT4 position_1553_add_4_22_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[20]), .I3(n40487), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_22 (.CI(n40487), .I0(direction_N_3806), 
            .I1(encoder0_position[20]), .CO(n40488));
    SB_LUT4 position_1553_add_4_21_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[19]), .I3(n40486), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_21 (.CI(n40486), .I0(direction_N_3806), 
            .I1(encoder0_position[19]), .CO(n40487));
    SB_LUT4 position_1553_add_4_20_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[18]), .I3(n40485), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_20 (.CI(n40485), .I0(direction_N_3806), 
            .I1(encoder0_position[18]), .CO(n40486));
    SB_LUT4 position_1553_add_4_19_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[17]), .I3(n40484), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_19 (.CI(n40484), .I0(direction_N_3806), 
            .I1(encoder0_position[17]), .CO(n40485));
    SB_LUT4 position_1553_add_4_18_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[16]), .I3(n40483), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_18 (.CI(n40483), .I0(direction_N_3806), 
            .I1(encoder0_position[16]), .CO(n40484));
    SB_LUT4 position_1553_add_4_17_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[15]), .I3(n40482), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_17 (.CI(n40482), .I0(direction_N_3806), 
            .I1(encoder0_position[15]), .CO(n40483));
    SB_DFF debounce_cnt_50 (.Q(debounce_cnt), .C(n1188), .D(a_prev_N_3813));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 position_1553_add_4_16_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[14]), .I3(n40481), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_16 (.CI(n40481), .I0(direction_N_3806), 
            .I1(encoder0_position[14]), .CO(n40482));
    SB_LUT4 position_1553_add_4_15_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[13]), .I3(n40480), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_15 (.CI(n40480), .I0(direction_N_3806), 
            .I1(encoder0_position[13]), .CO(n40481));
    SB_LUT4 position_1553_add_4_14_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[12]), .I3(n40479), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_14 (.CI(n40479), .I0(direction_N_3806), 
            .I1(encoder0_position[12]), .CO(n40480));
    SB_LUT4 position_1553_add_4_13_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[11]), .I3(n40478), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_13 (.CI(n40478), .I0(direction_N_3806), 
            .I1(encoder0_position[11]), .CO(n40479));
    SB_LUT4 position_1553_add_4_12_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[10]), .I3(n40477), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_12 (.CI(n40477), .I0(direction_N_3806), 
            .I1(encoder0_position[10]), .CO(n40478));
    SB_LUT4 position_1553_add_4_11_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[9]), .I3(n40476), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_11 (.CI(n40476), .I0(direction_N_3806), 
            .I1(encoder0_position[9]), .CO(n40477));
    SB_LUT4 position_1553_add_4_10_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[8]), .I3(n40475), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_10 (.CI(n40475), .I0(direction_N_3806), 
            .I1(encoder0_position[8]), .CO(n40476));
    SB_LUT4 position_1553_add_4_9_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[7]), .I3(n40474), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_9 (.CI(n40474), .I0(direction_N_3806), 
            .I1(encoder0_position[7]), .CO(n40475));
    SB_LUT4 position_1553_add_4_8_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[6]), .I3(n40473), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_8 (.CI(n40473), .I0(direction_N_3806), 
            .I1(encoder0_position[6]), .CO(n40474));
    SB_LUT4 position_1553_add_4_7_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[5]), .I3(n40472), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_7 (.CI(n40472), .I0(direction_N_3806), 
            .I1(encoder0_position[5]), .CO(n40473));
    SB_LUT4 position_1553_add_4_6_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[4]), .I3(n40471), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_6 (.CI(n40471), .I0(direction_N_3806), 
            .I1(encoder0_position[4]), .CO(n40472));
    SB_LUT4 position_1553_add_4_5_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[3]), .I3(n40470), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_5 (.CI(n40470), .I0(direction_N_3806), 
            .I1(encoder0_position[3]), .CO(n40471));
    SB_LUT4 position_1553_add_4_4_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[2]), .I3(n40469), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_4 (.CI(n40469), .I0(direction_N_3806), 
            .I1(encoder0_position[2]), .CO(n40470));
    SB_LUT4 position_1553_add_4_3_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder0_position[1]), .I3(n40468), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_3 (.CI(n40468), .I0(direction_N_3806), 
            .I1(encoder0_position[1]), .CO(n40469));
    SB_LUT4 position_1553_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder0_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1553_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1553_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder0_position[0]), 
            .CO(n40468));
    SB_DFF a_new_i1 (.Q(a_new[1]), .C(n1188), .D(a_new_c[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1188), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_prev_51 (.Q(a_prev), .C(n1188), .D(n28243));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_prev_52 (.Q(b_prev), .C(n1188), .D(n28242));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF direction_57 (.Q(n1152), .C(n1188), .D(n28241));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 i35760_4_lut (.I0(a_new_c[0]), .I1(b_new[0]), .I2(a_new[1]), 
            .I3(b_new[1]), .O(a_prev_N_3813));   // vhdl/quadrature_decoder.vhd(57[8:58])
    defparam i35760_4_lut.LUT_INIT = 16'h8421;
    SB_LUT4 b_prev_I_0_63_2_lut (.I0(b_prev), .I1(a_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3806));   // vhdl/quadrature_decoder.vhd(81[18:37])
    defparam b_prev_I_0_63_2_lut.LUT_INIT = 16'h9999;
    SB_DFFE position_1553__i0 (.Q(encoder0_position[0]), .C(n1188), .E(direction_N_3807), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i1 (.Q(encoder0_position[1]), .C(n1188), .E(direction_N_3807), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i2 (.Q(encoder0_position[2]), .C(n1188), .E(direction_N_3807), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i3 (.Q(encoder0_position[3]), .C(n1188), .E(direction_N_3807), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i4 (.Q(encoder0_position[4]), .C(n1188), .E(direction_N_3807), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i5 (.Q(encoder0_position[5]), .C(n1188), .E(direction_N_3807), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i6 (.Q(encoder0_position[6]), .C(n1188), .E(direction_N_3807), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i7 (.Q(encoder0_position[7]), .C(n1188), .E(direction_N_3807), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i8 (.Q(encoder0_position[8]), .C(n1188), .E(direction_N_3807), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i9 (.Q(encoder0_position[9]), .C(n1188), .E(direction_N_3807), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i10 (.Q(encoder0_position[10]), .C(n1188), .E(direction_N_3807), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i11 (.Q(encoder0_position[11]), .C(n1188), .E(direction_N_3807), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i12 (.Q(encoder0_position[12]), .C(n1188), .E(direction_N_3807), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i13 (.Q(encoder0_position[13]), .C(n1188), .E(direction_N_3807), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i14 (.Q(encoder0_position[14]), .C(n1188), .E(direction_N_3807), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i15 (.Q(encoder0_position[15]), .C(n1188), .E(direction_N_3807), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i16 (.Q(encoder0_position[16]), .C(n1188), .E(direction_N_3807), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i17 (.Q(encoder0_position[17]), .C(n1188), .E(direction_N_3807), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i18 (.Q(encoder0_position[18]), .C(n1188), .E(direction_N_3807), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i19 (.Q(encoder0_position[19]), .C(n1188), .E(direction_N_3807), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i20 (.Q(encoder0_position[20]), .C(n1188), .E(direction_N_3807), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i21 (.Q(encoder0_position[21]), .C(n1188), .E(direction_N_3807), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i22 (.Q(encoder0_position[22]), .C(n1188), .E(direction_N_3807), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i23 (.Q(encoder0_position[23]), .C(n1188), .E(direction_N_3807), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i24 (.Q(encoder0_position[24]), .C(n1188), .E(direction_N_3807), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i25 (.Q(encoder0_position[25]), .C(n1188), .E(direction_N_3807), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i26 (.Q(encoder0_position[26]), .C(n1188), .E(direction_N_3807), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i27 (.Q(encoder0_position[27]), .C(n1188), .E(direction_N_3807), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i28 (.Q(encoder0_position[28]), .C(n1188), .E(direction_N_3807), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i29 (.Q(encoder0_position[29]), .C(n1188), .E(direction_N_3807), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i30 (.Q(encoder0_position[30]), .C(n1188), .E(direction_N_3807), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1553__i31 (.Q(encoder0_position[31]), .C(n1188), .E(direction_N_3807), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_LUT4 i15180_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3813), .I2(a_new[1]), 
            .I3(a_prev), .O(n28243));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i15180_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15179_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3813), .I2(b_new[1]), 
            .I3(b_prev), .O(n28242));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i15179_3_lut_4_lut.LUT_INIT = 16'hf780;
    
endmodule
//
// Verilog Description of module \quadrature_decoder(1,500000) 
//

module \quadrature_decoder(1,500000)  (b_prev, GND_net, a_new, direction_N_3807, 
            ENCODER1_B_N_keep, n1188, ENCODER1_A_N_keep, encoder1_position, 
            VCC_net, n28234, n1193) /* synthesis lattice_noprune=1 */ ;
    output b_prev;
    input GND_net;
    output [1:0]a_new;
    output direction_N_3807;
    input ENCODER1_B_N_keep;
    input n1188;
    input ENCODER1_A_N_keep;
    output [31:0]encoder1_position;
    input VCC_net;
    input n28234;
    output n1193;
    
    wire [1:0]b_new;   // vhdl/quadrature_decoder.vhd(41[9:14])
    
    wire direction_N_3810, debounce_cnt, a_prev, a_prev_N_3813, n28240, 
        n28227;
    wire [1:0]a_new_c;   // vhdl/quadrature_decoder.vhd(40[9:14])
    wire [31:0]n133;
    
    wire direction_N_3806, n40452, n40451, n40450, n40449, n40448, 
        n40447, n40446, n40445, n40444, n40443, n40442, n40441, 
        n40440, n40439, n40438, n40437, n40436, n40435, n40434, 
        n40433, n40432, n40431, n40430, n40429, n40428, n40427, 
        n40426, n40425, n40424, n40423, n40422;
    
    SB_LUT4 b_prev_I_0_65_2_lut (.I0(b_prev), .I1(b_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3810));   // vhdl/quadrature_decoder.vhd(80[37:56])
    defparam b_prev_I_0_65_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 debounce_cnt_I_0_4_lut (.I0(debounce_cnt), .I1(a_prev), .I2(direction_N_3810), 
            .I3(a_new[1]), .O(direction_N_3807));   // vhdl/quadrature_decoder.vhd(79[10] 80[64])
    defparam debounce_cnt_I_0_4_lut.LUT_INIT = 16'ha2a8;
    SB_LUT4 i15177_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3813), .I2(b_new[1]), 
            .I3(b_prev), .O(n28240));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i15177_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i15164_3_lut_4_lut (.I0(debounce_cnt), .I1(a_prev_N_3813), .I2(a_new[1]), 
            .I3(a_prev), .O(n28227));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i15164_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_DFF b_new_i0 (.Q(b_new[0]), .C(n1188), .D(ENCODER1_B_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i0 (.Q(a_new_c[0]), .C(n1188), .D(ENCODER1_A_N_keep));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF debounce_cnt_50 (.Q(debounce_cnt), .C(n1188), .D(a_prev_N_3813));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_new_i1 (.Q(a_new[1]), .C(n1188), .D(a_new_c[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF b_new_i1 (.Q(b_new[1]), .C(n1188), .D(b_new[0]));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_LUT4 position_1548_add_4_33_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[31]), .I3(n40452), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 position_1548_add_4_32_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[30]), .I3(n40451), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_32 (.CI(n40451), .I0(direction_N_3806), 
            .I1(encoder1_position[30]), .CO(n40452));
    SB_LUT4 position_1548_add_4_31_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[29]), .I3(n40450), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_31 (.CI(n40450), .I0(direction_N_3806), 
            .I1(encoder1_position[29]), .CO(n40451));
    SB_LUT4 position_1548_add_4_30_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[28]), .I3(n40449), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_30 (.CI(n40449), .I0(direction_N_3806), 
            .I1(encoder1_position[28]), .CO(n40450));
    SB_LUT4 position_1548_add_4_29_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[27]), .I3(n40448), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_29 (.CI(n40448), .I0(direction_N_3806), 
            .I1(encoder1_position[27]), .CO(n40449));
    SB_LUT4 position_1548_add_4_28_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[26]), .I3(n40447), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_28 (.CI(n40447), .I0(direction_N_3806), 
            .I1(encoder1_position[26]), .CO(n40448));
    SB_LUT4 position_1548_add_4_27_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[25]), .I3(n40446), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_27 (.CI(n40446), .I0(direction_N_3806), 
            .I1(encoder1_position[25]), .CO(n40447));
    SB_LUT4 position_1548_add_4_26_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[24]), .I3(n40445), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_26 (.CI(n40445), .I0(direction_N_3806), 
            .I1(encoder1_position[24]), .CO(n40446));
    SB_LUT4 position_1548_add_4_25_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[23]), .I3(n40444), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_25 (.CI(n40444), .I0(direction_N_3806), 
            .I1(encoder1_position[23]), .CO(n40445));
    SB_LUT4 position_1548_add_4_24_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[22]), .I3(n40443), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_24 (.CI(n40443), .I0(direction_N_3806), 
            .I1(encoder1_position[22]), .CO(n40444));
    SB_LUT4 position_1548_add_4_23_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[21]), .I3(n40442), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_23 (.CI(n40442), .I0(direction_N_3806), 
            .I1(encoder1_position[21]), .CO(n40443));
    SB_LUT4 position_1548_add_4_22_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[20]), .I3(n40441), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_22 (.CI(n40441), .I0(direction_N_3806), 
            .I1(encoder1_position[20]), .CO(n40442));
    SB_LUT4 position_1548_add_4_21_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[19]), .I3(n40440), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_21 (.CI(n40440), .I0(direction_N_3806), 
            .I1(encoder1_position[19]), .CO(n40441));
    SB_LUT4 position_1548_add_4_20_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[18]), .I3(n40439), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_20 (.CI(n40439), .I0(direction_N_3806), 
            .I1(encoder1_position[18]), .CO(n40440));
    SB_LUT4 position_1548_add_4_19_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[17]), .I3(n40438), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_19 (.CI(n40438), .I0(direction_N_3806), 
            .I1(encoder1_position[17]), .CO(n40439));
    SB_LUT4 position_1548_add_4_18_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[16]), .I3(n40437), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_18 (.CI(n40437), .I0(direction_N_3806), 
            .I1(encoder1_position[16]), .CO(n40438));
    SB_LUT4 position_1548_add_4_17_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[15]), .I3(n40436), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_17 (.CI(n40436), .I0(direction_N_3806), 
            .I1(encoder1_position[15]), .CO(n40437));
    SB_LUT4 position_1548_add_4_16_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[14]), .I3(n40435), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_16 (.CI(n40435), .I0(direction_N_3806), 
            .I1(encoder1_position[14]), .CO(n40436));
    SB_LUT4 position_1548_add_4_15_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[13]), .I3(n40434), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_15 (.CI(n40434), .I0(direction_N_3806), 
            .I1(encoder1_position[13]), .CO(n40435));
    SB_LUT4 position_1548_add_4_14_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[12]), .I3(n40433), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_14 (.CI(n40433), .I0(direction_N_3806), 
            .I1(encoder1_position[12]), .CO(n40434));
    SB_LUT4 position_1548_add_4_13_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[11]), .I3(n40432), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_13 (.CI(n40432), .I0(direction_N_3806), 
            .I1(encoder1_position[11]), .CO(n40433));
    SB_LUT4 position_1548_add_4_12_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[10]), .I3(n40431), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_12 (.CI(n40431), .I0(direction_N_3806), 
            .I1(encoder1_position[10]), .CO(n40432));
    SB_LUT4 position_1548_add_4_11_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[9]), .I3(n40430), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_11 (.CI(n40430), .I0(direction_N_3806), 
            .I1(encoder1_position[9]), .CO(n40431));
    SB_LUT4 position_1548_add_4_10_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[8]), .I3(n40429), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_10 (.CI(n40429), .I0(direction_N_3806), 
            .I1(encoder1_position[8]), .CO(n40430));
    SB_LUT4 position_1548_add_4_9_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[7]), .I3(n40428), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_9 (.CI(n40428), .I0(direction_N_3806), 
            .I1(encoder1_position[7]), .CO(n40429));
    SB_LUT4 position_1548_add_4_8_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[6]), .I3(n40427), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_8 (.CI(n40427), .I0(direction_N_3806), 
            .I1(encoder1_position[6]), .CO(n40428));
    SB_LUT4 position_1548_add_4_7_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[5]), .I3(n40426), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_7 (.CI(n40426), .I0(direction_N_3806), 
            .I1(encoder1_position[5]), .CO(n40427));
    SB_LUT4 position_1548_add_4_6_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[4]), .I3(n40425), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_6 (.CI(n40425), .I0(direction_N_3806), 
            .I1(encoder1_position[4]), .CO(n40426));
    SB_LUT4 position_1548_add_4_5_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[3]), .I3(n40424), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_5 (.CI(n40424), .I0(direction_N_3806), 
            .I1(encoder1_position[3]), .CO(n40425));
    SB_LUT4 position_1548_add_4_4_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[2]), .I3(n40423), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_4 (.CI(n40423), .I0(direction_N_3806), 
            .I1(encoder1_position[2]), .CO(n40424));
    SB_LUT4 position_1548_add_4_3_lut (.I0(GND_net), .I1(direction_N_3806), 
            .I2(encoder1_position[1]), .I3(n40422), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_3 (.CI(n40422), .I0(direction_N_3806), 
            .I1(encoder1_position[1]), .CO(n40423));
    SB_LUT4 position_1548_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(encoder1_position[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam position_1548_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY position_1548_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(encoder1_position[0]), 
            .CO(n40422));
    SB_LUT4 b_prev_I_0_63_2_lut (.I0(b_prev), .I1(a_new[1]), .I2(GND_net), 
            .I3(GND_net), .O(direction_N_3806));   // vhdl/quadrature_decoder.vhd(81[18:37])
    defparam b_prev_I_0_63_2_lut.LUT_INIT = 16'h9999;
    SB_DFF b_prev_52 (.Q(b_prev), .C(n1188), .D(n28240));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF direction_57 (.Q(n1193), .C(n1188), .D(n28234));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFF a_prev_51 (.Q(a_prev), .C(n1188), .D(n28227));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    SB_DFFE position_1548__i0 (.Q(encoder1_position[0]), .C(n1188), .E(direction_N_3807), 
            .D(n133[0]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_LUT4 i35741_4_lut (.I0(a_new_c[0]), .I1(b_new[0]), .I2(a_new[1]), 
            .I3(b_new[1]), .O(a_prev_N_3813));   // vhdl/quadrature_decoder.vhd(52[3] 89[10])
    defparam i35741_4_lut.LUT_INIT = 16'h8421;
    SB_DFFE position_1548__i1 (.Q(encoder1_position[1]), .C(n1188), .E(direction_N_3807), 
            .D(n133[1]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i2 (.Q(encoder1_position[2]), .C(n1188), .E(direction_N_3807), 
            .D(n133[2]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i3 (.Q(encoder1_position[3]), .C(n1188), .E(direction_N_3807), 
            .D(n133[3]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i4 (.Q(encoder1_position[4]), .C(n1188), .E(direction_N_3807), 
            .D(n133[4]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i5 (.Q(encoder1_position[5]), .C(n1188), .E(direction_N_3807), 
            .D(n133[5]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i6 (.Q(encoder1_position[6]), .C(n1188), .E(direction_N_3807), 
            .D(n133[6]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i7 (.Q(encoder1_position[7]), .C(n1188), .E(direction_N_3807), 
            .D(n133[7]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i8 (.Q(encoder1_position[8]), .C(n1188), .E(direction_N_3807), 
            .D(n133[8]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i9 (.Q(encoder1_position[9]), .C(n1188), .E(direction_N_3807), 
            .D(n133[9]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i10 (.Q(encoder1_position[10]), .C(n1188), .E(direction_N_3807), 
            .D(n133[10]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i11 (.Q(encoder1_position[11]), .C(n1188), .E(direction_N_3807), 
            .D(n133[11]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i12 (.Q(encoder1_position[12]), .C(n1188), .E(direction_N_3807), 
            .D(n133[12]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i13 (.Q(encoder1_position[13]), .C(n1188), .E(direction_N_3807), 
            .D(n133[13]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i14 (.Q(encoder1_position[14]), .C(n1188), .E(direction_N_3807), 
            .D(n133[14]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i15 (.Q(encoder1_position[15]), .C(n1188), .E(direction_N_3807), 
            .D(n133[15]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i16 (.Q(encoder1_position[16]), .C(n1188), .E(direction_N_3807), 
            .D(n133[16]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i17 (.Q(encoder1_position[17]), .C(n1188), .E(direction_N_3807), 
            .D(n133[17]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i18 (.Q(encoder1_position[18]), .C(n1188), .E(direction_N_3807), 
            .D(n133[18]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i19 (.Q(encoder1_position[19]), .C(n1188), .E(direction_N_3807), 
            .D(n133[19]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i20 (.Q(encoder1_position[20]), .C(n1188), .E(direction_N_3807), 
            .D(n133[20]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i21 (.Q(encoder1_position[21]), .C(n1188), .E(direction_N_3807), 
            .D(n133[21]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i22 (.Q(encoder1_position[22]), .C(n1188), .E(direction_N_3807), 
            .D(n133[22]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i23 (.Q(encoder1_position[23]), .C(n1188), .E(direction_N_3807), 
            .D(n133[23]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i24 (.Q(encoder1_position[24]), .C(n1188), .E(direction_N_3807), 
            .D(n133[24]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i25 (.Q(encoder1_position[25]), .C(n1188), .E(direction_N_3807), 
            .D(n133[25]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i26 (.Q(encoder1_position[26]), .C(n1188), .E(direction_N_3807), 
            .D(n133[26]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i27 (.Q(encoder1_position[27]), .C(n1188), .E(direction_N_3807), 
            .D(n133[27]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i28 (.Q(encoder1_position[28]), .C(n1188), .E(direction_N_3807), 
            .D(n133[28]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i29 (.Q(encoder1_position[29]), .C(n1188), .E(direction_N_3807), 
            .D(n133[29]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i30 (.Q(encoder1_position[30]), .C(n1188), .E(direction_N_3807), 
            .D(n133[30]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    SB_DFFE position_1548__i31 (.Q(encoder1_position[31]), .C(n1188), .E(direction_N_3807), 
            .D(n133[31]));   // vhdl/quadrature_decoder.vhd(77[4] 87[11])
    
endmodule
//
// Verilog Description of module pll32MHz
//

module pll32MHz (GND_net, CLK_c, VCC_net, clk32MHz) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input CLK_c;
    input VCC_net;
    output clk32MHz;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    
    SB_PLL40_CORE pll32MHz_inst (.REFERENCECLK(CLK_c), .PLLOUTGLOBAL(clk32MHz), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=51, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=37 */ ;   // verilog/TinyFPGA_B.v(34[10] 37[2])
    defparam pll32MHz_inst.FEEDBACK_PATH = "PHASE_AND_DELAY";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam pll32MHz_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam pll32MHz_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam pll32MHz_inst.FDA_FEEDBACK = 4'b0000;
    defparam pll32MHz_inst.FDA_RELATIVE = 4'b0000;
    defparam pll32MHz_inst.PLLOUT_SELECT = "SHIFTREG_0deg";
    defparam pll32MHz_inst.DIVR = 4'b0000;
    defparam pll32MHz_inst.DIVF = 7'b0000001;
    defparam pll32MHz_inst.DIVQ = 3'b011;
    defparam pll32MHz_inst.FILTER_RANGE = 3'b001;
    defparam pll32MHz_inst.ENABLE_ICEGATE = 1'b0;
    defparam pll32MHz_inst.TEST_MODE = 1'b0;
    defparam pll32MHz_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module motorControl
//

module motorControl (\Kp[3] , GND_net, \Ki[8] , \Kp[13] , \Kp[4] , 
            \Kp[14] , \Ki[9] , \Kp[5] , PWMLimit, \Ki[3] , \Kp[15] , 
            \Ki[10] , \Kp[6] , \Kp[7] , \Kp[8] , \Kp[9] , \Ki[11] , 
            \Kp[10] , \Ki[4] , \Ki[5] , \Ki[0] , \Kp[0] , \Kp[11] , 
            \Ki[6] , \Ki[12] , \Kp[12] , \Ki[7] , \Ki[13] , \Ki[14] , 
            \Ki[15] , \Ki[1] , \Ki[2] , \Kp[1] , \Kp[2] , IntegralLimit, 
            duty, clk32MHz, VCC_net, setpoint, motor_state, n51409) /* synthesis syn_module_defined=1 */ ;
    input \Kp[3] ;
    input GND_net;
    input \Ki[8] ;
    input \Kp[13] ;
    input \Kp[4] ;
    input \Kp[14] ;
    input \Ki[9] ;
    input \Kp[5] ;
    input [23:0]PWMLimit;
    input \Ki[3] ;
    input \Kp[15] ;
    input \Ki[10] ;
    input \Kp[6] ;
    input \Kp[7] ;
    input \Kp[8] ;
    input \Kp[9] ;
    input \Ki[11] ;
    input \Kp[10] ;
    input \Ki[4] ;
    input \Ki[5] ;
    input \Ki[0] ;
    input \Kp[0] ;
    input \Kp[11] ;
    input \Ki[6] ;
    input \Ki[12] ;
    input \Kp[12] ;
    input \Ki[7] ;
    input \Ki[13] ;
    input \Ki[14] ;
    input \Ki[15] ;
    input \Ki[1] ;
    input \Ki[2] ;
    input \Kp[1] ;
    input \Kp[2] ;
    input [23:0]IntegralLimit;
    output [23:0]duty;
    input clk32MHz;
    input VCC_net;
    input [23:0]setpoint;
    input [23:0]motor_state;
    output n51409;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [23:0]n1;
    
    wire n220;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3572 ;
    
    wire n591, n968, n293;
    wire [15:0]n15821;
    wire [14:0]n16365;
    
    wire n241, n39461, n1041;
    wire [20:0]n11628;
    wire [19:0]n12924;
    
    wire n226, n39569, n679, n664, n366, n971;
    wire [23:0]n1_adj_4767;
    
    wire n39570, n256, n40000;
    wire [20:0]n12113;
    
    wire n515, n40001, n1114, n39269, n39270, n752, n737, n439, 
        n512;
    wire [21:0]n9870;
    
    wire n442, n39999, n153, n39568, n585, n658, n39883;
    wire [14:0]n16620;
    
    wire n1117, n39884, n810, n369, n39998, n731, n329, n402, 
        n825;
    wire [47:0]n155;
    wire [47:0]n106;
    
    wire n804, n475, n883, n877, n548, n956, n950, n621, n1023, 
        n1096, n898, n448, n971_adj_4346, n694, n1029, n1044, 
        n1102, n1117_adj_4347, n743, n521, n92, n23_adj_4348, \PID_CONTROLLER.integral_23__N_3620 ;
    wire [23:0]n3616;
    
    wire n767, n165, n1044_adj_4350, n39462, n296, n39997, n77, 
        n8_adj_4351, n840, n150;
    wire [15:0]n16109;
    
    wire n39882, n39881, n238, n223, n296_adj_4352, n168, n39460, 
        n898_adj_4353, n39880, n26_adj_4354, n95, n816;
    wire [23:0]n257;
    
    wire n39268, n101, n39267, n32, n889, n11_adj_4355, n80;
    wire [7:0]n18685;
    wire [6:0]n18812;
    
    wire n630, n39459, n962, n594, n1035, n1108, n557, n39458, 
        n484, n39457, n39266, n39265, n311, n369_adj_4356, n174, 
        n247, n667, n320;
    wire [23:0]n1_adj_4768;
    
    wire n223_adj_4358, n39996, n384, n393, n740, n825_adj_4360, 
        n39879, n150_adj_4361, n39995;
    wire [18:0]n13765;
    
    wire n39567, n39264, n39566, n39565, n411, n39456, n125, n56, 
        n466, n101_adj_4364, n32_adj_4365, n539, n813, n174_adj_4367, 
        n612, n886, n959, n685, n1032, n758, n1105, n831, n198, 
        n271_adj_4369, n904, n977, n344, n247_adj_4370, n39564, 
        n752_adj_4371, n39878;
    wire [23:0]duty_23__N_3548;
    
    wire n1050, n417, n6_adj_4372;
    wire [3:0]n19005;
    wire [4:0]n18945;
    
    wire n98, n29;
    wire [23:0]\PID_CONTROLLER.integral ;   // verilog/motorControl.v(23[23:31])
    
    wire n204, n338, n39455, n265, n39454;
    wire [1:0]n19069;
    
    wire n131, n62, n39263;
    wire [9:0]n18205;
    wire [8:0]n18425;
    
    wire n770, n39358, n679_adj_4374, n39877, n697, n39357, n192, 
        n39453, n624, n39356, n442_adj_4375, n4_adj_4376;
    wire [2:0]n19045;
    
    wire n490, n12_adj_4377, n8_adj_4378, n8_adj_4379, n77_adj_4380, 
        n11_adj_4381, n6_adj_4382, n50, n119, n38742, n18_adj_4383, 
        n551, n39355, n13_adj_4384, n4_adj_4385, n46537, n39262, 
        n122, n53, n320_adj_4387, n171, n457, n39563, n530, n113;
    wire [19:0]n13364;
    
    wire n39994, n39993, n44, n39992;
    wire [13:0]n16845;
    
    wire n1120, n39452, n606, n39876, n244, n317, n39261, n80_adj_4396, 
        n89, n20_adj_4398, n11_adj_4399, n195, n17_adj_4400, n9_adj_4401, 
        n11_adj_4402, n49965, n49961, n51890, n50401, n50216, n39991, 
        n162, n515_adj_4403, n51872, n50212, n603, n235, n50205, 
        n51865, n27, n15_adj_4404, n13_adj_4405, n11_adj_4406, n49859, 
        n21_adj_4407, n19_adj_4408, n17_adj_4409, n9_adj_4410, n49866, 
        n43, n16_adj_4411, n49842, n8_adj_4412, n45, n24_adj_4413, 
        n7_adj_4414, n5_adj_4415, n49876, n50181, n588, n676, n661, 
        n50177, n25_adj_4416, n23_adj_4417, n50543, n31, n29_adj_4418, 
        n50373, n37, n35, n33, n50605, n50219, n51859, n50199, 
        n478, n39354, n51853, n12_adj_4419, n49893, n125_adj_4420, 
        n56_adj_4421, n308, n51877, n10_adj_4422, n1105_adj_4423, 
        n39562, n39260, n749, n533, n39875, n30, n734, n50463, 
        n49905, n381, n51857, n454, n1047, n39451, n50389, n51883, 
        n50555, n51848, n527, n50633, n51845, n198_adj_4425, n600, 
        n16_adj_4426, n1032_adj_4427, n39561, n49878, n822, n271_adj_4428, 
        n895, n24_adj_4429, n807, n6_adj_4430, n50527, n673, n959_adj_4431, 
        n39560, n50528, n49880, n8_adj_4432, n51843, n50475, n50470;
    wire [23:0]\PID_CONTROLLER.integral_23__N_3623 ;
    
    wire n3_adj_4433, n4_adj_4434, n50545, n50546, n12_adj_4435, n405, 
        n39353, n49852, n10_adj_4436, n30_adj_4437, n49854, n974, 
        n39450, n50625, n39259, n50480, n50667, n901, n39449, 
        n886_adj_4439, n39559, n50668, n39, n50652, n6_adj_4440, 
        n332, n39352, n813_adj_4441, n39558, n828, n39448, n50547, 
        n50548, n259, n39351, n49844, n50483, n50478, n41, n49846, 
        n50569, n40, n50571, n4_adj_4442, n50551, n50552, n39258, 
        n49899, n50623, n50472, n50665, n50666, n50654, n49882, 
        n755, n39447, n460, n39874, n186, n39350, n39257, n50563, 
        n740_adj_4445, n39557, n40_adj_4446, \PID_CONTROLLER.integral_23__N_3622 , 
        n50565, n39990, n387, n39873, n667_adj_4447, n39556, n44_adj_4448, 
        n113_adj_4449, n39256, n682, n39446, n594_adj_4452, n39555, 
        n186_adj_4453, n390, n268_adj_4455, n39989, n153_adj_4456, 
        n393_adj_4457, n341, n521_adj_4458, n39554, n226_adj_4459;
    wire [7:0]n18605;
    
    wire n700, n39349, n466_adj_4460, n314, n39872, n463, n627, 
        n39348, n609, n39445, n536, n39444, n414, n554, n39347, 
        n448_adj_4463, n39553, n539_adj_4465, n1102_adj_4467, n39988, 
        n487, n536_adj_4468, n1029_adj_4469, n39987, n375, n39552, 
        n299, n463_adj_4470, n39443, n560, n481, n39346, n241_adj_4472, 
        n39871, n39255, n612_adj_4474, n259_adj_4475, n119_adj_4476, 
        n50_adj_4477, n685_adj_4478, n372, n332_adj_4479, n445, n302, 
        n39551, n39254, n192_adj_4482, n956_adj_4483, n39986, n609_adj_4484, 
        n168_adj_4485, n39870, n408, n39345, n229, n39550, n39253, 
        n390_adj_4487, n39442, n883_adj_4488, n39985, n810_adj_4489, 
        n39984, n518, n405_adj_4490, n758_adj_4491, n682_adj_4492, 
        n265_adj_4493, n317_adj_4494, n39441, n26_adj_4496, n95_adj_4497, 
        n156, n39549, n737_adj_4498, n39983;
    wire [13:0]n17069;
    
    wire n1120_adj_4499, n39869, n335, n39344, n1047_adj_4500, n39868, 
        n39252, n244_adj_4502, n39440, n664_adj_4503, n39982, n262, 
        n39343, n14_adj_4504, n83, n344_adj_4505, n171_adj_4506, n39439, 
        n189, n39342, n39251, n968_adj_4508, n1041_adj_4509, n39250, 
        n880;
    wire [9:0]n18325;
    wire [8:0]n18524;
    
    wire n770_adj_4511, n39548, n953, n697_adj_4512, n39547, n746, 
        n819, n892, n1026, n417_adj_4513, n47, n116, n6_adj_4514;
    wire [3:0]n19029;
    wire [4:0]n18980;
    
    wire n974_adj_4515, n39867, n29_adj_4516, n98_adj_4517;
    wire [6:0]n18749;
    
    wire n630_adj_4518, n39341, n557_adj_4519, n39340;
    wire [1:0]n19077;
    
    wire n591_adj_4520, n39981, n901_adj_4521, n39866, n39249, n624_adj_4523, 
        n39546, n4_adj_4524;
    wire [2:0]n19060;
    
    wire n490_adj_4525, n12_adj_4526;
    wire [12:0]n17265;
    
    wire n1050_adj_4527, n39438, n8_adj_4528, n484_adj_4529, n39339, 
        n977_adj_4530, n39437, n551_adj_4531, n39545, n411_adj_4532, 
        n39338, n39248, n11_adj_4534, n904_adj_4535, n39436, n831_adj_4536, 
        n39435, n39247, n338_adj_4538, n39337, n828_adj_4539, n39865, 
        n755_adj_4540, n39864, n39246, n6_adj_4542, n478_adj_4543, 
        n39544, n39245, n39336, n39863, n39434, n39543, n39980, 
        n39862, n39335, n38783, n18_adj_4544, n13_adj_4545, n39244, 
        n4_adj_4546, n46504, n39979, n965, n1099, n39542, n39978, 
        n39433, n39541, n39432;
    wire [5:0]n18861;
    
    wire n39334, n39243, n39977, n39861, n39333, n39242, n1114_adj_4547, 
        n107, n38, n39431, n107_adj_4549, n38_adj_4551, n1038;
    wire [23:0]duty_23__N_3672;
    
    wire n256_adj_4552;
    wire [23:0]duty_23__N_3647;
    
    wire duty_23__N_3671, n39241, n39332, n39240, n39860, n39430, 
        n39976, n39331, n39429, n39975, n39330, n39239, n39859, 
        n1111, n116_adj_4556, n47_adj_4557, n39540, n189_adj_4558, 
        n180, n180_adj_4559, n262_adj_4560, n39158, n253, n39329, 
        n253_adj_4561, n86, n17_adj_4563, n39238, n39858, n326, 
        n39157, n399;
    wire [18:0]n14164;
    
    wire n39974, n39857, n159, n232, n335_adj_4564, n305, n39237, 
        n39156, n378, n472, n39856, n39973, n451, n326_adj_4565, 
        n408_adj_4566, n39428, n74, n5_adj_4567, n524, n147, n481_adj_4568, 
        n545, n597, n39328, n220_adj_4569, n670, n39972, n618, 
        n39327;
    wire [12:0]n17460;
    
    wire n39855, n743_adj_4570, n691, n554_adj_4571, n816_adj_4572, 
        n889_adj_4573, n764, n399_adj_4574, n837, n910, n962_adj_4575, 
        n293_adj_4576, n472_adj_4577, n39427, n39971, n39326, n39854, 
        n39236, n39853, n39970, n366_adj_4578, n39235, n627_adj_4579, 
        n545_adj_4580, n39325, n1035_adj_4581, n439_adj_4582, n700_adj_4583, 
        n512_adj_4584, n89_adj_4585, n20_adj_4586, n39324, n39852, 
        n39969, n39851, n39968, n39155, n39850, n39967, n104, 
        n39966, n35_adj_4587, n618_adj_4588, n1108_adj_4589, n39849, 
        n39426, n177, n691_adj_4590, n162_adj_4591, n764_adj_4592, 
        n39965, n585_adj_4593, n39848, n39234, n39847, n39233, n39154, 
        n39964, n39846, n39153;
    wire [17:0]n14525;
    
    wire n39533, n39845, n39963, n39844, n39843, n39532, n39531, 
        n39232, n39152, n39530, n39231, n39529, n39528, n39962, 
        n39527, n39230, n39229, n658_adj_4594, n235_adj_4595, n308_adj_4596, 
        n731_adj_4597, n110, n41_adj_4598, n381_adj_4599, n250, n804_adj_4600, 
        n39526, n183, n837_adj_4601, n454_adj_4602, n910_adj_4603, 
        n39151, n39525, n527_adj_4604, n256_adj_4605, n877_adj_4606, 
        n104_adj_4607, n35_adj_4608, n323, n600_adj_4609, n673_adj_4610, 
        n950_adj_4611, n177_adj_4612, n250_adj_4613, n39150, n746_adj_4614, 
        n39961, n83_adj_4615, n39228, n39524, n14_adj_4616, n39227, 
        n39960;
    wire [11:0]n17797;
    
    wire n980, n39842, n39149, n907, n39841, n323_adj_4617, n396, 
        n670_adj_4618, n39523, n375_adj_4619, n39959, n834, n39840, 
        n469, n39226, n597_adj_4620, n39522, n524_adj_4621, n39521, 
        n39225, n761, n39839, n39148, n396_adj_4622;
    wire [0:0]n8832;
    wire [21:0]n9339;
    
    wire n39630, n39629, n451_adj_4623, n39520, n302_adj_4624, n39958;
    wire [10:0]n18084;
    
    wire n840_adj_4625, n39734, n39628, n378_adj_4626, n39519, n767_adj_4627, 
        n39733;
    wire [5:0]n18909;
    
    wire n560_adj_4628, n39414, n487_adj_4629, n39413, n688, n39838, 
        n694_adj_4630, n39732, n39224, n39147, n305_adj_4631, n39518, 
        n414_adj_4632, n39412, n232_adj_4633, n39517, n159_adj_4634, 
        n39516, n39223, n341_adj_4635, n39411, n39222, n268_adj_4636, 
        n39410, n39146, n469_adj_4637, n819_adj_4638, n329_adj_4639, 
        n542, n39627, n892_adj_4641, n1023_adj_4642, n1096_adj_4643, 
        n39145, n17_adj_4644, n86_adj_4645, n39221, n39626;
    wire [16:0]n15209;
    
    wire n39515, n39144, n195_adj_4646, n39409, n39220, n615, n39837, 
        n39514, n39625, n615_adj_4647, n402_adj_4648, n965_adj_4649, 
        n39143, n39219, n39142, n53_adj_4650, n122_adj_4651, n475_adj_4652, 
        n621_adj_4653, n39731, n39513;
    wire [11:0]n17629;
    
    wire n980_adj_4654, n39408, n907_adj_4655, n39407, n39218, n39141, 
        n229_adj_4656, n39957, n39624, n688_adj_4658, n39217, n1111_adj_4659, 
        n39512, n39140, n834_adj_4660, n39406, n548_adj_4661, n39730, 
        n156_adj_4662, n39956, n542_adj_4663, n39836, n1038_adj_4664, 
        n39511, n761_adj_4665, n39405, n39216, n39404, n39139, n39138, 
        n39729, n39215, n39137, n39623, n39510, n39728, n39403, 
        n39622, n39621, n39509, n39214, n39402, n39727, n39136, 
        n39508, n39401, n39213, n39400, n39835, n39212;
    wire [0:0]n9363;
    
    wire n39135, n39834, n39134, n39399, n39211, n39210, n39133, 
        n39507;
    wire [17:0]n14885;
    
    wire n39955, n39398, n39954, n39397, n39620, n39132, n39506, 
        n39131, n39505, n39833, n39953, n39130, n39619, n39726, 
        n39504;
    wire [10:0]n17941;
    
    wire n39396, n39503, n39395, n39129, n39725, n39618, n39832, 
        n39502, n39617, n39952, n39501, n39500, n39616, n39615, 
        n39128, n39394, n39499, n39393, n39831, n39951, n39392, 
        n39614, n39498, n39613, n39950, n39127, n39391, n39497, 
        n39612, n39390, n39611, n39949, n39830, n39829, n39389, 
        n39828, n39948, n39947, n39496, n39827, n39946, n39826, 
        n39945, n39126, n39610, n39944, n39825, n39495, n39609, 
        n39943, n39494, n39388, n39942, n39824, n39125, n39608, 
        n39941, n39607, n39940, n39493, n39939, n39938, n39823, 
        n39606, n39822, n39821, n39387, n39605;
    wire [16:0]n15532;
    
    wire n39937, n39492, n39936, n39124, n39935, n39604, n39820, 
        n39386, n39491, n39603, n50075, n50086, n39934, n50113, 
        n39933, n39602, n39490, n39489, n39488, n39123, n39601, 
        n39932, n39385, n39384, n39122, n39600, n50123, n39931, 
        n39930, n39121, n39929, n39599, n39598, n39487, n39486, 
        n39383, n39120, n50111, n6_adj_4670, n49840, n6_adj_4671, 
        n39928, n39119, n39597, n39485, n39382, n39484, n39927, 
        n39381, n39926, n39118, n39925, n39924, n39596, n39483, 
        n39923, n39595, n39482, n39594, n39922, n39481, n39593, 
        n39921, n39117, n39116, n39480, n39115, n39479, n39278, 
        n39277, n39592, n39114, n39478, n39591, n39477, n39276, 
        n39590, n39113, n39589, n39476, n39588, n39375, n39587, 
        n39586, n39275, n39585, n39475, n39374, n39584, n39583, 
        n39474, n39473, n39582, n39581, n39472, n39580, n40037, 
        n40036, n39373, n40035, n39471, n40034, n40033, n40032, 
        n40031, n39470, n40030, n40029, n40028, n39372, n40027, 
        n39579, n39371, n40026, n39578, n39370, n39274, n40025, 
        n39469, n39369, n39368, n39273, n40024, n39577, n40023, 
        n40022, n39900, n39899, n40021, n40020, n39576, n39468, 
        n39898, n39367, n39272, n40019, n39575, n39467, n39897, 
        n40018, n39896, n39574, n40017, n895_adj_4675, n39895, n147_adj_4676, 
        n40016, n5_adj_4677, n74_adj_4678, n822_adj_4679, n39894, 
        n749_adj_4680, n39893, n518_adj_4681, n39573, n183_adj_4682, 
        n39366, n39271, n606_adj_4684, n39466, n676_adj_4685, n39892, 
        n40015, n603_adj_4686, n39891, n533_adj_4687, n39465, n445_adj_4688, 
        n39572, n530_adj_4690, n39890, n460_adj_4691, n39464, n41_adj_4692, 
        n110_adj_4693, n40014, n457_adj_4694, n39889, n372_adj_4695, 
        n39571, n384_adj_4696, n39888, n40013, n311_adj_4697, n39887, 
        n299_adj_4698, n238_adj_4699, n39886, n387_adj_4700, n39463, 
        n40012, n40011, n40010, n40009, n1099_adj_4701, n40008, 
        n165_adj_4702, n39885, n1026_adj_4703, n40007, n953_adj_4704, 
        n40006, n880_adj_4705, n40005, n807_adj_4706, n40004, n23_adj_4707, 
        n92_adj_4708, n734_adj_4709, n40003, n314_adj_4710, n661_adj_4711, 
        n40002, n588_adj_4712, n39_adj_4713, n41_adj_4714, n45_adj_4715, 
        n37_adj_4716, n29_adj_4717, n31_adj_4718, n43_adj_4719, n35_adj_4720, 
        n23_adj_4721, n25_adj_4722, n33_adj_4723, n9_adj_4724, n17_adj_4725, 
        n19_adj_4726, n21_adj_4727, n11_adj_4728, n13_adj_4729, n15_adj_4730, 
        n27_adj_4731, n49830, n49823, n12_adj_4732, n10_adj_4733, 
        n30_adj_4734, n50148, n50144, n50529, n50357, n50603, n16_adj_4735, 
        n50539, n50540, n8_adj_4736, n24_adj_4737, n50115, n50487, 
        n50486, n4_adj_4738, n50501, n50502, n50128, n50585, n50232, 
        n50647, n50648, n50644, n50117, n50609, n50238, n50611, 
        n41_adj_4739, n39_adj_4740, n45_adj_4741, n43_adj_4742, n37_adj_4743, 
        n29_adj_4744, n31_adj_4745, n21_adj_4746, n23_adj_4747, n25_adj_4748, 
        n17_adj_4749, n19_adj_4750, n9_adj_4751, n35_adj_4752, n33_adj_4753, 
        n11_adj_4754, n13_adj_4755, n38876, n15_adj_4756, n38901, 
        n4_adj_4757, n27_adj_4758, n50101, n38935, n50093, n12_adj_4759, 
        n10_adj_4760, n30_adj_4761, n50337, n50333, n50599, n50435, 
        n50627, n16_adj_4762, n50495, n50496, n8_adj_4763, n24_adj_4764, 
        n50077, n50489, n50240, n4_adj_4765, n50493, n50494, n50088, 
        n50587, n50242, n50649, n50650, n50640, n50079, n50613, 
        n50248, n50615, n4_adj_4766, n38833, n38758;
    
    SB_LUT4 mult_10_i149_2_lut (.I0(\Kp[3] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n220));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i398_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n591));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i651_2_lut (.I0(\Kp[13] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n968));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i198_2_lut (.I0(\Kp[4] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n293));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5857_4_lut (.I0(GND_net), .I1(n16365[1]), .I2(n241), .I3(n39461), 
            .O(n15821[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5857_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i700_2_lut (.I0(\Kp[14] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1041));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5299_4_lut (.I0(GND_net), .I1(n12924[1]), .I2(n226), .I3(n39569), 
            .O(n11628[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i457_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n679));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i447_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n664));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i247_2_lut (.I0(\Kp[5] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n366));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i653_2_lut (.I0(\Kp[13] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n971));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i18_1_lut (.I0(PWMLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[17]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5299_4 (.CI(n39569), .I0(n12924[1]), .I1(n226), .CO(n39570));
    SB_LUT4 mult_11_i173_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n256));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i173_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4077_8 (.CI(n40000), .I0(n12113[5]), .I1(n515), .CO(n40001));
    SB_LUT4 mult_10_i749_2_lut (.I0(\Kp[15] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n1114));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i749_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_16 (.CI(n39269), .I0(GND_net), .I1(n1_adj_4767[14]), 
            .CO(n39270));
    SB_LUT4 mult_11_i506_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n752));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i496_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n737));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i296_2_lut (.I0(\Kp[6] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n439));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i345_2_lut (.I0(\Kp[7] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n512));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4077_7_lut (.I0(GND_net), .I1(n12113[4]), .I2(n442), .I3(n39999), 
            .O(n9870[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5299_3_lut (.I0(GND_net), .I1(n12924[0]), .I2(n153), .I3(n39568), 
            .O(n11628[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4077_7 (.CI(n39999), .I0(n12113[4]), .I1(n442), .CO(n40000));
    SB_LUT4 mult_10_i394_2_lut (.I0(\Kp[8] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n585));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i443_2_lut (.I0(\Kp[9] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n658));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i443_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5873_16 (.CI(n39883), .I0(n16620[13]), .I1(n1117), .CO(n39884));
    SB_LUT4 mult_11_i545_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n810));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_4077_6_lut (.I0(GND_net), .I1(n12113[3]), .I2(n369), .I3(n39998), 
            .O(n9870[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i492_2_lut (.I0(\Kp[10] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n731));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i19_1_lut (.I0(PWMLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[18]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i222_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n329));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i271_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n402));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i555_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n825));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i2_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n155[0]));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i2_2_lut (.I0(\Kp[0] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n106[0]));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i541_2_lut (.I0(\Kp[11] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n804));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i20_1_lut (.I0(PWMLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[19]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i320_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n475));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i320_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i594_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n883));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i590_2_lut (.I0(\Kp[12] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n877));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i369_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n548));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i643_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n956));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i639_2_lut (.I0(\Kp[13] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n950));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i418_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n621));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i688_2_lut (.I0(\Kp[14] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1023));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i737_2_lut (.I0(\Kp[15] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n1096));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i737_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i604_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n898));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i302_2_lut (.I0(\Kp[6] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n448));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i653_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n971_adj_4346));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i653_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i467_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n694));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i692_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1029));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i702_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1044));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i741_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n1102));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i751_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n1117_adj_4347));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i500_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n743));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i351_2_lut (.I0(\Kp[7] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n521));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i63_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n92));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i16_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4348));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20692_2_lut (.I0(n1[15]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[15]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i516_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n767));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i112_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n165));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i21_1_lut (.I0(PWMLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[20]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i702_2_lut (.I0(\Kp[14] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1044_adj_4350));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i702_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4077_6 (.CI(n39998), .I0(n12113[3]), .I1(n369), .CO(n39999));
    SB_CARRY add_5857_4 (.CI(n39461), .I0(n16365[1]), .I1(n241), .CO(n39462));
    SB_LUT4 add_4077_5_lut (.I0(GND_net), .I1(n12113[2]), .I2(n296), .I3(n39997), 
            .O(n9870[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i200_2_lut (.I0(\Kp[4] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n296));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i53_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n77));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i6_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4351));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i565_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n840));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i102_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n150));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5873_15_lut (.I0(GND_net), .I1(n16620[12]), .I2(n1044_adj_4350), 
            .I3(n39882), .O(n16109[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5873_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5873_15 (.CI(n39882), .I0(n16620[12]), .I1(n1044_adj_4350), 
            .CO(n39883));
    SB_LUT4 add_5873_14_lut (.I0(GND_net), .I1(n16620[11]), .I2(n971), 
            .I3(n39881), .O(n16109[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5873_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i161_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n238));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i151_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n223));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i151_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4077_5 (.CI(n39997), .I0(n12113[2]), .I1(n296), .CO(n39998));
    SB_LUT4 mult_11_i200_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n296_adj_4352));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i200_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5857_3_lut (.I0(GND_net), .I1(n16365[0]), .I2(n168), .I3(n39460), 
            .O(n15821[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5857_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5873_14 (.CI(n39881), .I0(n16620[11]), .I1(n971), .CO(n39882));
    SB_CARRY add_5299_3 (.CI(n39568), .I0(n12924[0]), .I1(n153), .CO(n39569));
    SB_LUT4 add_5873_13_lut (.I0(GND_net), .I1(n16620[10]), .I2(n898_adj_4353), 
            .I3(n39880), .O(n16109[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5873_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5873_13 (.CI(n39880), .I0(n16620[10]), .I1(n898_adj_4353), 
            .CO(n39881));
    SB_CARRY add_5857_3 (.CI(n39460), .I0(n16365[0]), .I1(n168), .CO(n39461));
    SB_LUT4 add_5857_2_lut (.I0(GND_net), .I1(n26_adj_4354), .I2(n95), 
            .I3(GND_net), .O(n15821[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5857_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i549_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n816));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_15_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[13]), 
            .I3(n39268), .O(n257[13])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20691_2_lut (.I0(n1[16]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[16]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20691_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_16_add_3_15 (.CI(n39268), .I0(GND_net), .I1(n1_adj_4767[13]), 
            .CO(n39269));
    SB_LUT4 mult_10_i69_2_lut (.I0(\Kp[1] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n101));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_14_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[12]), 
            .I3(n39267), .O(n257[12])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_14 (.CI(n39267), .I0(GND_net), .I1(n1_adj_4767[12]), 
            .CO(n39268));
    SB_LUT4 mult_10_i22_2_lut (.I0(\Kp[0] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n32));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i598_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n889));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5299_2_lut (.I0(GND_net), .I1(n11_adj_4355), .I2(n80), 
            .I3(GND_net), .O(n11628[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5299_2 (.CI(GND_net), .I0(n11_adj_4355), .I1(n80), .CO(n39568));
    SB_CARRY add_5857_2 (.CI(GND_net), .I0(n26_adj_4354), .I1(n95), .CO(n39460));
    SB_LUT4 add_6057_9_lut (.I0(GND_net), .I1(n18812[6]), .I2(n630), .I3(n39459), 
            .O(n18685[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6057_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i647_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n962));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i400_2_lut (.I0(\Kp[8] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n594));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i696_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1035));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i745_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n1108));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20690_2_lut (.I0(n1[17]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[17]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6057_8_lut (.I0(GND_net), .I1(n18812[5]), .I2(n557), .I3(n39458), 
            .O(n18685[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6057_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6057_8 (.CI(n39458), .I0(n18812[5]), .I1(n557), .CO(n39459));
    SB_LUT4 add_6057_7_lut (.I0(GND_net), .I1(n18812[4]), .I2(n484), .I3(n39457), 
            .O(n18685[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6057_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_13_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[11]), 
            .I3(n39266), .O(n257[11])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_13 (.CI(n39266), .I0(GND_net), .I1(n1_adj_4767[11]), 
            .CO(n39267));
    SB_LUT4 unary_minus_16_add_3_12_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[10]), 
            .I3(n39265), .O(n257[10])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i22_1_lut (.I0(PWMLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[21]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i210_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n311));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i249_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n369_adj_4356));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i118_2_lut (.I0(\Kp[2] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n174));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i167_2_lut (.I0(\Kp[3] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n247));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i167_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i449_2_lut (.I0(\Kp[9] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n667));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i216_2_lut (.I0(\Kp[4] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n320));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i1_1_lut (.I0(IntegralLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[0]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_4077_4_lut (.I0(GND_net), .I1(n12113[1]), .I2(n223_adj_4358), 
            .I3(n39996), .O(n9870[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i259_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n384));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20689_2_lut (.I0(n1[18]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[18]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20689_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i265_2_lut (.I0(\Kp[5] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n393));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i265_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i498_2_lut (.I0(\Kp[10] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n740));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i498_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4077_4 (.CI(n39996), .I0(n12113[1]), .I1(n223_adj_4358), 
            .CO(n39997));
    SB_LUT4 add_5873_12_lut (.I0(GND_net), .I1(n16620[9]), .I2(n825_adj_4360), 
            .I3(n39879), .O(n16109[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5873_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4077_3_lut (.I0(GND_net), .I1(n12113[0]), .I2(n150_adj_4361), 
            .I3(n39995), .O(n9870[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_12 (.CI(n39265), .I0(GND_net), .I1(n1_adj_4767[10]), 
            .CO(n39266));
    SB_LUT4 add_5712_21_lut (.I0(GND_net), .I1(n13765[18]), .I2(GND_net), 
            .I3(n39567), .O(n12924[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_11_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[9]), 
            .I3(n39264), .O(n257[9])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6057_7 (.CI(n39457), .I0(n18812[4]), .I1(n484), .CO(n39458));
    SB_LUT4 add_5712_20_lut (.I0(GND_net), .I1(n13765[17]), .I2(GND_net), 
            .I3(n39566), .O(n12924[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5712_20 (.CI(n39566), .I0(n13765[17]), .I1(GND_net), 
            .CO(n39567));
    SB_LUT4 add_5712_19_lut (.I0(GND_net), .I1(n13765[16]), .I2(GND_net), 
            .I3(n39565), .O(n12924[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20688_2_lut (.I0(n1[19]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[19]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i2_1_lut (.I0(IntegralLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[1]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6057_6_lut (.I0(GND_net), .I1(n18812[3]), .I2(n411), .I3(n39456), 
            .O(n18685[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6057_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i85_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n125));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i38_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [18]), 
            .I2(GND_net), .I3(GND_net), .O(n56));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i314_2_lut (.I0(\Kp[6] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n466));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i69_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n101_adj_4364));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i69_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i22_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n32_adj_4365));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i22_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i3_1_lut (.I0(IntegralLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[2]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i363_2_lut (.I0(\Kp[7] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n539));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i547_2_lut (.I0(\Kp[11] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n813));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i118_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n174_adj_4367));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i118_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i412_2_lut (.I0(\Kp[8] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n612));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i596_2_lut (.I0(\Kp[12] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n886));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i645_2_lut (.I0(\Kp[13] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n959));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i461_2_lut (.I0(\Kp[9] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n685));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20687_2_lut (.I0(n1[20]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[20]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20687_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i694_2_lut (.I0(\Kp[14] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1032));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i510_2_lut (.I0(\Kp[10] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n758));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i510_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i743_2_lut (.I0(\Kp[15] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n1105));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i743_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i559_2_lut (.I0(\Kp[11] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n831));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i134_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n198));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i183_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n271_adj_4369));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i183_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i4_1_lut (.I0(IntegralLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[3]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i608_2_lut (.I0(\Kp[12] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n904));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i608_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i5_1_lut (.I0(IntegralLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[4]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i657_2_lut (.I0(\Kp[13] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n977));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i657_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i232_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n344));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i167_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n247_adj_4370));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i167_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4077_3 (.CI(n39995), .I0(n12113[0]), .I1(n150_adj_4361), 
            .CO(n39996));
    SB_CARRY add_6057_6 (.CI(n39456), .I0(n18812[3]), .I1(n411), .CO(n39457));
    SB_CARRY add_5873_12 (.CI(n39879), .I0(n16620[9]), .I1(n825_adj_4360), 
            .CO(n39880));
    SB_CARRY add_5712_19 (.CI(n39565), .I0(n13765[16]), .I1(GND_net), 
            .CO(n39566));
    SB_LUT4 add_5712_18_lut (.I0(GND_net), .I1(n13765[15]), .I2(GND_net), 
            .I3(n39564), .O(n12924[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5873_11_lut (.I0(GND_net), .I1(n16620[8]), .I2(n752_adj_4371), 
            .I3(n39878), .O(n16109[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5873_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5873_11 (.CI(n39878), .I0(n16620[8]), .I1(n752_adj_4371), 
            .CO(n39879));
    SB_DFF result_i0 (.Q(duty[0]), .C(clk32MHz), .D(duty_23__N_3548[0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_10_i706_2_lut (.I0(\Kp[14] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n1050));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i281_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n417));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut (.I0(n6_adj_4372), .I1(\Ki[4] ), .I2(n19005[2]), 
            .I3(\PID_CONTROLLER.integral_23__N_3572 [18]), .O(n18945[3]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut.LUT_INIT = 16'h965a;
    SB_LUT4 mult_10_i67_2_lut (.I0(\Kp[1] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n98));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i67_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i20_2_lut (.I0(\Kp[0] ), .I1(n1[9]), .I2(GND_net), 
            .I3(GND_net), .O(n29));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i20_2_lut.LUT_INIT = 16'h8888;
    SB_DFF \PID_CONTROLLER.integral_i0  (.Q(\PID_CONTROLLER.integral [0]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [0]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 mult_11_i138_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n204));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i138_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6057_5_lut (.I0(GND_net), .I1(n18812[2]), .I2(n338), .I3(n39455), 
            .O(n18685[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6057_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6057_5 (.CI(n39455), .I0(n18812[2]), .I1(n338), .CO(n39456));
    SB_LUT4 add_6057_4_lut (.I0(GND_net), .I1(n18812[1]), .I2(n265), .I3(n39454), 
            .O(n18685[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6057_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25722_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3572 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3572 [21]), .O(n19069[0]));   // verilog/motorControl.v(34[25:36])
    defparam i25722_4_lut.LUT_INIT = 16'h6ca0;
    SB_CARRY unary_minus_16_add_3_11 (.CI(n39264), .I0(GND_net), .I1(n1_adj_4767[9]), 
            .CO(n39265));
    SB_LUT4 mult_11_i89_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [19]), 
            .I2(GND_net), .I3(GND_net), .O(n131));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i89_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i42_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [20]), 
            .I2(GND_net), .I3(GND_net), .O(n62));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i42_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_10_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[8]), 
            .I3(n39263), .O(n257[8])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6013_11_lut (.I0(GND_net), .I1(n18425[8]), .I2(n770), 
            .I3(n39358), .O(n18205[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6013_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5873_10_lut (.I0(GND_net), .I1(n16620[7]), .I2(n679_adj_4374), 
            .I3(n39877), .O(n16109[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5873_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6013_10_lut (.I0(GND_net), .I1(n18425[7]), .I2(n697), 
            .I3(n39357), .O(n18205[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6013_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6057_4 (.CI(n39454), .I0(n18812[1]), .I1(n265), .CO(n39455));
    SB_CARRY add_6013_10 (.CI(n39357), .I0(n18425[7]), .I1(n697), .CO(n39358));
    SB_CARRY add_5712_18 (.CI(n39564), .I0(n13765[15]), .I1(GND_net), 
            .CO(n39565));
    SB_LUT4 add_6057_3_lut (.I0(GND_net), .I1(n18812[0]), .I2(n192), .I3(n39453), 
            .O(n18685[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6057_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6057_3 (.CI(n39453), .I0(n18812[0]), .I1(n192), .CO(n39454));
    SB_LUT4 add_6013_9_lut (.I0(GND_net), .I1(n18425[6]), .I2(n624), .I3(n39356), 
            .O(n18205[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6013_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i298_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n442_adj_4375));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i298_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1522 (.I0(n4_adj_4376), .I1(\Ki[3] ), .I2(n19045[1]), 
            .I3(\PID_CONTROLLER.integral_23__N_3572 [19]), .O(n19005[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1522.LUT_INIT = 16'h965a;
    SB_LUT4 mult_11_i330_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n490));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i330_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6013_9 (.CI(n39356), .I0(n18425[6]), .I1(n624), .CO(n39357));
    SB_LUT4 i2_4_lut_adj_1523 (.I0(\Ki[0] ), .I1(\Ki[3] ), .I2(\PID_CONTROLLER.integral_23__N_3572 [23]), 
            .I3(\PID_CONTROLLER.integral_23__N_3572 [20]), .O(n12_adj_4377));   // verilog/motorControl.v(34[25:36])
    defparam i2_4_lut_adj_1523.LUT_INIT = 16'h9c50;
    SB_LUT4 i25835_4_lut (.I0(n19005[2]), .I1(\Ki[4] ), .I2(n6_adj_4372), 
            .I3(\PID_CONTROLLER.integral_23__N_3572 [18]), .O(n8_adj_4378));   // verilog/motorControl.v(34[25:36])
    defparam i25835_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 add_4077_2_lut (.I0(GND_net), .I1(n8_adj_4379), .I2(n77_adj_4380), 
            .I3(GND_net), .O(n9870[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_4_lut (.I0(\Ki[4] ), .I1(\Ki[2] ), .I2(\PID_CONTROLLER.integral_23__N_3572 [19]), 
            .I3(\PID_CONTROLLER.integral_23__N_3572 [21]), .O(n11_adj_4381));   // verilog/motorControl.v(34[25:36])
    defparam i1_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 i25796_4_lut (.I0(n19045[1]), .I1(\Ki[3] ), .I2(n4_adj_4376), 
            .I3(\PID_CONTROLLER.integral_23__N_3572 [19]), .O(n6_adj_4382));   // verilog/motorControl.v(34[25:36])
    defparam i25796_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 add_6057_2_lut (.I0(GND_net), .I1(n50), .I2(n119), .I3(GND_net), 
            .O(n18685[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6057_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25724_4_lut (.I0(\Ki[0] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3572 [22]), 
            .I3(\PID_CONTROLLER.integral_23__N_3572 [21]), .O(n38742));   // verilog/motorControl.v(34[25:36])
    defparam i25724_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY unary_minus_16_add_3_10 (.CI(n39263), .I0(GND_net), .I1(n1_adj_4767[8]), 
            .CO(n39264));
    SB_LUT4 i8_4_lut (.I0(n6_adj_4382), .I1(n11_adj_4381), .I2(n8_adj_4378), 
            .I3(n12_adj_4377), .O(n18_adj_4383));   // verilog/motorControl.v(34[25:36])
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6013_8_lut (.I0(GND_net), .I1(n18425[5]), .I2(n551), .I3(n39355), 
            .O(n18205[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6013_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i3_4_lut (.I0(\Ki[5] ), .I1(\Ki[1] ), .I2(\PID_CONTROLLER.integral_23__N_3572 [18]), 
            .I3(\PID_CONTROLLER.integral_23__N_3572 [22]), .O(n13_adj_4384));   // verilog/motorControl.v(34[25:36])
    defparam i3_4_lut.LUT_INIT = 16'h6ca0;
    SB_CARRY add_4077_2 (.CI(GND_net), .I0(n8_adj_4379), .I1(n77_adj_4380), 
            .CO(n39995));
    SB_LUT4 i9_4_lut (.I0(n13_adj_4384), .I1(n18_adj_4383), .I2(n38742), 
            .I3(n4_adj_4385), .O(n46537));   // verilog/motorControl.v(34[25:36])
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 unary_minus_16_add_3_9_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[7]), 
            .I3(n39262), .O(n257[7])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_9 (.CI(n39262), .I0(GND_net), .I1(n1_adj_4767[7]), 
            .CO(n39263));
    SB_LUT4 mult_11_i83_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n122));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i36_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [17]), 
            .I2(GND_net), .I3(GND_net), .O(n53));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i216_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n320_adj_4387));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i216_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i116_2_lut (.I0(\Kp[2] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n171));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i23_1_lut (.I0(PWMLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[22]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i24_1_lut (.I0(PWMLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[23]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5873_10 (.CI(n39877), .I0(n16620[7]), .I1(n679_adj_4374), 
            .CO(n39878));
    SB_LUT4 mult_11_i308_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n457));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5712_17_lut (.I0(GND_net), .I1(n13765[14]), .I2(GND_net), 
            .I3(n39563), .O(n12924[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6057_2 (.CI(GND_net), .I0(n50), .I1(n119), .CO(n39453));
    SB_LUT4 mult_11_i357_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n530));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i77_2_lut (.I0(\Kp[1] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n113));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5322_22_lut (.I0(GND_net), .I1(n13364[19]), .I2(GND_net), 
            .I3(n39994), .O(n12113[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5322_21_lut (.I0(GND_net), .I1(n13364[18]), .I2(GND_net), 
            .I3(n39993), .O(n12113[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i30_2_lut (.I0(\Kp[0] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n44));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i30_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5322_21 (.CI(n39993), .I0(n13364[18]), .I1(GND_net), 
            .CO(n39994));
    SB_CARRY add_5712_17 (.CI(n39563), .I0(n13765[14]), .I1(GND_net), 
            .CO(n39564));
    SB_LUT4 add_5322_20_lut (.I0(GND_net), .I1(n13364[17]), .I2(GND_net), 
            .I3(n39992), .O(n12113[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5888_16_lut (.I0(GND_net), .I1(n16845[13]), .I2(n1120), 
            .I3(n39452), .O(n16365[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5888_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20686_2_lut (.I0(n1[21]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[21]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20686_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6013_8 (.CI(n39355), .I0(n18425[5]), .I1(n551), .CO(n39356));
    SB_LUT4 add_5873_9_lut (.I0(GND_net), .I1(n16620[6]), .I2(n606), .I3(n39876), 
            .O(n16109[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5873_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i6_1_lut (.I0(IntegralLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[5]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5873_9 (.CI(n39876), .I0(n16620[6]), .I1(n606), .CO(n39877));
    SB_LUT4 mult_10_i165_2_lut (.I0(\Kp[3] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n244));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20685_2_lut (.I0(n1[22]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[22]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20685_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i214_2_lut (.I0(\Kp[4] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n317));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_add_3_8_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[6]), 
            .I3(n39261), .O(n257[6])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i7_1_lut (.I0(IntegralLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[6]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i55_2_lut (.I0(\Kp[1] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n80_adj_4396));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i61_2_lut (.I0(\Kp[1] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n89));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i14_2_lut (.I0(\Kp[0] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n20_adj_4398));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i8_2_lut (.I0(\Kp[0] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n11_adj_4399));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i132_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n195));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i17_2_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(IntegralLimit[8]), .I2(GND_net), .I3(GND_net), .O(n17_adj_4400));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i9_2_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(IntegralLimit[4]), .I2(GND_net), .I3(GND_net), .O(n9_adj_4401));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i11_2_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(IntegralLimit[5]), .I2(GND_net), .I3(GND_net), .O(n11_adj_4402));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35013_4_lut (.I0(\PID_CONTROLLER.integral [3]), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(IntegralLimit[3]), .I3(IntegralLimit[2]), .O(n49965));
    defparam i35013_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 i35009_3_lut (.I0(n11_adj_4402), .I1(n9_adj_4401), .I2(n49965), 
            .I3(GND_net), .O(n49961));
    defparam i35009_3_lut.LUT_INIT = 16'habab;
    SB_LUT4 IntegralLimit_23__I_0_i13_rep_217_2_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(IntegralLimit[6]), .I2(GND_net), .I3(GND_net), .O(n51890));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i13_rep_217_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35448_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n51890), 
            .I2(IntegralLimit[7]), .I3(n49961), .O(n50401));
    defparam i35448_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i35264_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4400), 
            .I2(IntegralLimit[9]), .I3(n50401), .O(n50216));
    defparam i35264_4_lut.LUT_INIT = 16'hdeff;
    SB_CARRY add_5322_20 (.CI(n39992), .I0(n13364[17]), .I1(GND_net), 
            .CO(n39993));
    SB_LUT4 add_5322_19_lut (.I0(GND_net), .I1(n13364[16]), .I2(GND_net), 
            .I3(n39991), .O(n12113[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i110_2_lut (.I0(\Kp[2] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n162));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i347_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n515_adj_4403));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i21_rep_199_2_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(IntegralLimit[10]), .I2(GND_net), .I3(GND_net), .O(n51872));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i21_rep_199_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35260_4_lut (.I0(\PID_CONTROLLER.integral [9]), .I1(n17_adj_4400), 
            .I2(IntegralLimit[9]), .I3(n9_adj_4401), .O(n50212));
    defparam i35260_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 mult_11_i406_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n603));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i159_2_lut (.I0(\Kp[3] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n235));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35253_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n51872), 
            .I2(IntegralLimit[11]), .I3(n50212), .O(n50205));
    defparam i35253_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 IntegralLimit_23__I_0_i25_rep_192_2_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(IntegralLimit[12]), .I2(GND_net), .I3(GND_net), .O(n51865));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i25_rep_192_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34907_4_lut (.I0(n27), .I1(n15_adj_4404), .I2(n13_adj_4405), 
            .I3(n11_adj_4406), .O(n49859));
    defparam i34907_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34914_4_lut (.I0(n21_adj_4407), .I1(n19_adj_4408), .I2(n17_adj_4409), 
            .I3(n9_adj_4410), .O(n49866));
    defparam i34914_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i16_3_lut  (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(\PID_CONTROLLER.integral [21]), .I2(n43), .I3(GND_net), 
            .O(n16_adj_4411));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i16_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i34890_2_lut (.I0(n43), .I1(n19_adj_4408), .I2(GND_net), .I3(GND_net), 
            .O(n49842));
    defparam i34890_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i8_3_lut  (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(\PID_CONTROLLER.integral [8]), .I2(n17_adj_4409), .I3(GND_net), 
            .O(n8_adj_4412));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i8_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i24_3_lut  (.I0(n16_adj_4411), 
            .I1(\PID_CONTROLLER.integral [22]), .I2(n45), .I3(GND_net), 
            .O(n24_adj_4413));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i24_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 i34924_2_lut (.I0(n7_adj_4414), .I1(n5_adj_4415), .I2(GND_net), 
            .I3(GND_net), .O(n49876));
    defparam i34924_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i35229_4_lut (.I0(n13_adj_4405), .I1(n11_adj_4406), .I2(n9_adj_4410), 
            .I3(n49876), .O(n50181));
    defparam i35229_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 mult_11_i396_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n588));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i455_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n676));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i445_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n661));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35225_4_lut (.I0(n19_adj_4408), .I1(n17_adj_4409), .I2(n15_adj_4404), 
            .I3(n50181), .O(n50177));
    defparam i35225_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35590_4_lut (.I0(n25_adj_4416), .I1(n23_adj_4417), .I2(n21_adj_4407), 
            .I3(n50177), .O(n50543));
    defparam i35590_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35420_4_lut (.I0(n31), .I1(n29_adj_4418), .I2(n27), .I3(n50543), 
            .O(n50373));
    defparam i35420_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35652_4_lut (.I0(n37), .I1(n35), .I2(n33), .I3(n50373), 
            .O(n50605));
    defparam i35652_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35267_4_lut (.I0(\PID_CONTROLLER.integral [7]), .I1(n51890), 
            .I2(IntegralLimit[7]), .I3(n11_adj_4402), .O(n50219));
    defparam i35267_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i27_rep_186_2_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(IntegralLimit[13]), .I2(GND_net), .I3(GND_net), .O(n51859));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i27_rep_186_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35247_4_lut (.I0(\PID_CONTROLLER.integral [14]), .I1(n51859), 
            .I2(IntegralLimit[14]), .I3(n50219), .O(n50199));
    defparam i35247_4_lut.LUT_INIT = 16'hdeff;
    SB_LUT4 add_6013_7_lut (.I0(GND_net), .I1(n18425[4]), .I2(n478), .I3(n39354), 
            .O(n18205[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6013_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i31_rep_180_2_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(IntegralLimit[15]), .I2(GND_net), .I3(GND_net), .O(n51853));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i31_rep_180_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY unary_minus_16_add_3_8 (.CI(n39261), .I0(GND_net), .I1(n1_adj_4767[6]), 
            .CO(n39262));
    SB_LUT4 IntegralLimit_23__I_0_i12_3_lut (.I0(IntegralLimit[7]), .I1(IntegralLimit[16]), 
            .I2(\PID_CONTROLLER.integral [16]), .I3(GND_net), .O(n12_adj_4419));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i12_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34941_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(IntegralLimit[16]), .I3(IntegralLimit[7]), .O(n49893));
    defparam i34941_4_lut.LUT_INIT = 16'h7bde;
    SB_LUT4 mult_10_i85_2_lut (.I0(\Kp[1] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n125_adj_4420));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i85_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i38_2_lut (.I0(\Kp[0] ), .I1(n1[18]), .I2(GND_net), 
            .I3(GND_net), .O(n56_adj_4421));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i38_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i208_2_lut (.I0(\Kp[4] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n308));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i35_rep_204_2_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(IntegralLimit[17]), .I2(GND_net), .I3(GND_net), .O(n51877));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i35_rep_204_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 IntegralLimit_23__I_0_i10_3_lut (.I0(IntegralLimit[5]), .I1(IntegralLimit[6]), 
            .I2(\PID_CONTROLLER.integral [6]), .I3(GND_net), .O(n10_adj_4422));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i10_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5712_16_lut (.I0(GND_net), .I1(n13765[13]), .I2(n1105_adj_4423), 
            .I3(n39562), .O(n12924[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_7_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[5]), 
            .I3(n39260), .O(n257[5])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i504_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n749));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5873_8_lut (.I0(GND_net), .I1(n16620[5]), .I2(n533), .I3(n39875), 
            .O(n16109[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5873_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i30_3_lut (.I0(n12_adj_4419), .I1(IntegralLimit[17]), 
            .I2(\PID_CONTROLLER.integral [17]), .I3(GND_net), .O(n30));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i30_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i494_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n734));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35510_4_lut (.I0(\PID_CONTROLLER.integral [11]), .I1(n51872), 
            .I2(IntegralLimit[11]), .I3(n50216), .O(n50463));
    defparam i35510_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i34953_4_lut (.I0(\PID_CONTROLLER.integral [13]), .I1(n51865), 
            .I2(IntegralLimit[13]), .I3(n50463), .O(n49905));
    defparam i34953_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 mult_10_i257_2_lut (.I0(\Kp[5] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n381));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i29_rep_184_2_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(IntegralLimit[14]), .I2(GND_net), .I3(GND_net), .O(n51857));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i29_rep_184_2_lut.LUT_INIT = 16'h6666;
    SB_CARRY add_5712_16 (.CI(n39562), .I0(n13765[13]), .I1(n1105_adj_4423), 
            .CO(n39563));
    SB_LUT4 mult_10_i306_2_lut (.I0(\Kp[6] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n454));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5888_15_lut (.I0(GND_net), .I1(n16845[12]), .I2(n1047), 
            .I3(n39451), .O(n16365[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5888_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35436_4_lut (.I0(\PID_CONTROLLER.integral [15]), .I1(n51857), 
            .I2(IntegralLimit[15]), .I3(n49905), .O(n50389));
    defparam i35436_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i33_rep_210_2_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(IntegralLimit[16]), .I2(GND_net), .I3(GND_net), .O(n51883));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i33_rep_210_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35602_4_lut (.I0(\PID_CONTROLLER.integral [17]), .I1(n51883), 
            .I2(IntegralLimit[17]), .I3(n50389), .O(n50555));
    defparam i35602_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i37_rep_175_2_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(IntegralLimit[18]), .I2(GND_net), .I3(GND_net), .O(n51848));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i37_rep_175_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i355_2_lut (.I0(\Kp[7] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n527));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35680_4_lut (.I0(\PID_CONTROLLER.integral [19]), .I1(n51848), 
            .I2(IntegralLimit[19]), .I3(n50555), .O(n50633));
    defparam i35680_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 IntegralLimit_23__I_0_i41_rep_172_2_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(IntegralLimit[20]), .I2(GND_net), .I3(GND_net), .O(n51845));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i41_rep_172_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 mult_10_i134_2_lut (.I0(\Kp[2] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n198_adj_4425));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i134_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i404_2_lut (.I0(\Kp[8] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n600));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i16_3_lut (.I0(IntegralLimit[9]), .I1(IntegralLimit[21]), 
            .I2(\PID_CONTROLLER.integral [21]), .I3(GND_net), .O(n16_adj_4426));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i16_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 add_5712_15_lut (.I0(GND_net), .I1(n13765[12]), .I2(n1032_adj_4427), 
            .I3(n39561), .O(n12924[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34926_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(IntegralLimit[21]), .I3(IntegralLimit[9]), .O(n49878));
    defparam i34926_4_lut.LUT_INIT = 16'h7bde;
    SB_CARRY add_6013_7 (.CI(n39354), .I0(n18425[4]), .I1(n478), .CO(n39355));
    SB_LUT4 mult_11_i553_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n822));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i183_2_lut (.I0(\Kp[3] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n271_adj_4428));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i183_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5888_15 (.CI(n39451), .I0(n16845[12]), .I1(n1047), .CO(n39452));
    SB_LUT4 mult_11_i602_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n895));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i602_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i24_3_lut (.I0(n16_adj_4426), .I1(IntegralLimit[22]), 
            .I2(\PID_CONTROLLER.integral [22]), .I3(GND_net), .O(n24_adj_4429));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i24_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_11_i543_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n807));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i543_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5712_15 (.CI(n39561), .I0(n13765[12]), .I1(n1032_adj_4427), 
            .CO(n39562));
    SB_LUT4 IntegralLimit_23__I_0_i6_3_lut (.I0(IntegralLimit[2]), .I1(IntegralLimit[3]), 
            .I2(\PID_CONTROLLER.integral [3]), .I3(GND_net), .O(n6_adj_4430));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i6_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35574_3_lut (.I0(n6_adj_4430), .I1(IntegralLimit[10]), .I2(\PID_CONTROLLER.integral [10]), 
            .I3(GND_net), .O(n50527));   // verilog/motorControl.v(31[10:34])
    defparam i35574_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mult_10_i453_2_lut (.I0(\Kp[9] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n673));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5712_14_lut (.I0(GND_net), .I1(n13765[11]), .I2(n959_adj_4431), 
            .I3(n39560), .O(n12924[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35575_3_lut (.I0(n50527), .I1(IntegralLimit[11]), .I2(\PID_CONTROLLER.integral [11]), 
            .I3(GND_net), .O(n50528));   // verilog/motorControl.v(31[10:34])
    defparam i35575_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i34928_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n51865), 
            .I2(IntegralLimit[21]), .I3(n50205), .O(n49880));
    defparam i34928_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i35522_4_lut (.I0(n24_adj_4429), .I1(n8_adj_4432), .I2(n51843), 
            .I3(n49878), .O(n50475));   // verilog/motorControl.v(31[10:34])
    defparam i35522_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY unary_minus_16_add_3_7 (.CI(n39260), .I0(GND_net), .I1(n1_adj_4767[5]), 
            .CO(n39261));
    SB_LUT4 i35517_3_lut (.I0(n50528), .I1(IntegralLimit[12]), .I2(\PID_CONTROLLER.integral [12]), 
            .I3(GND_net), .O(n50470));   // verilog/motorControl.v(31[10:34])
    defparam i35517_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i4_4_lut  (.I0(\PID_CONTROLLER.integral_23__N_3623 [0]), 
            .I1(\PID_CONTROLLER.integral [1]), .I2(n3_adj_4433), .I3(\PID_CONTROLLER.integral [0]), 
            .O(n4_adj_4434));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i4_4_lut .LUT_INIT = 16'hc5c0;
    SB_CARRY add_5322_19 (.CI(n39991), .I0(n13364[16]), .I1(GND_net), 
            .CO(n39992));
    SB_LUT4 i35592_3_lut (.I0(n4_adj_4434), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n27), .I3(GND_net), .O(n50545));   // verilog/motorControl.v(31[38:63])
    defparam i35592_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35593_3_lut (.I0(n50545), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n29_adj_4418), .I3(GND_net), .O(n50546));   // verilog/motorControl.v(31[38:63])
    defparam i35593_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i12_3_lut  (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(\PID_CONTROLLER.integral [16]), .I2(n33), .I3(GND_net), 
            .O(n12_adj_4435));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i12_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 add_6013_6_lut (.I0(GND_net), .I1(n18425[3]), .I2(n405), .I3(n39353), 
            .O(n18205[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6013_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34900_2_lut (.I0(n33), .I1(n15_adj_4404), .I2(GND_net), .I3(GND_net), 
            .O(n49852));
    defparam i34900_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i10_3_lut  (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(\PID_CONTROLLER.integral [6]), .I2(n13_adj_4405), .I3(GND_net), 
            .O(n10_adj_4436));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i10_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i30_3_lut  (.I0(n12_adj_4435), 
            .I1(\PID_CONTROLLER.integral [17]), .I2(n35), .I3(GND_net), 
            .O(n30_adj_4437));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i30_3_lut .LUT_INIT = 16'hcaca;
    SB_CARRY add_5712_14 (.CI(n39560), .I0(n13765[11]), .I1(n959_adj_4431), 
            .CO(n39561));
    SB_LUT4 i34902_4_lut (.I0(n33), .I1(n31), .I2(n29_adj_4418), .I3(n49859), 
            .O(n49854));
    defparam i34902_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 add_5888_14_lut (.I0(GND_net), .I1(n16845[11]), .I2(n974), 
            .I3(n39450), .O(n16365[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5888_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35672_4_lut (.I0(n30_adj_4437), .I1(n10_adj_4436), .I2(n35), 
            .I3(n49852), .O(n50625));   // verilog/motorControl.v(31[38:63])
    defparam i35672_4_lut.LUT_INIT = 16'haaac;
    SB_CARRY add_5888_14 (.CI(n39450), .I0(n16845[11]), .I1(n974), .CO(n39451));
    SB_LUT4 unary_minus_16_add_3_6_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[4]), 
            .I3(n39259), .O(n257[4])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35527_3_lut (.I0(n50546), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n31), .I3(GND_net), .O(n50480));   // verilog/motorControl.v(31[38:63])
    defparam i35527_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35714_4_lut (.I0(n50480), .I1(n50625), .I2(n35), .I3(n49854), 
            .O(n50667));   // verilog/motorControl.v(31[38:63])
    defparam i35714_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_5888_13_lut (.I0(GND_net), .I1(n16845[10]), .I2(n901), 
            .I3(n39449), .O(n16365[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5888_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5712_13_lut (.I0(GND_net), .I1(n13765[10]), .I2(n886_adj_4439), 
            .I3(n39559), .O(n12924[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35715_3_lut (.I0(n50667), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n37), .I3(GND_net), .O(n50668));   // verilog/motorControl.v(31[38:63])
    defparam i35715_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5873_8 (.CI(n39875), .I0(n16620[5]), .I1(n533), .CO(n39876));
    SB_LUT4 i35699_3_lut (.I0(n50668), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n39), .I3(GND_net), .O(n50652));   // verilog/motorControl.v(31[38:63])
    defparam i35699_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6013_6 (.CI(n39353), .I0(n18425[3]), .I1(n405), .CO(n39354));
    SB_LUT4 \PID_CONTROLLER.integral_23__I_0_i6_3_lut  (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(\PID_CONTROLLER.integral [3]), .I2(n7_adj_4414), .I3(GND_net), 
            .O(n6_adj_4440));   // verilog/motorControl.v(31[38:63])
    defparam \PID_CONTROLLER.integral_23__I_0_i6_3_lut .LUT_INIT = 16'hcaca;
    SB_LUT4 add_6013_5_lut (.I0(GND_net), .I1(n18425[2]), .I2(n332), .I3(n39352), 
            .O(n18205[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6013_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5888_13 (.CI(n39449), .I0(n16845[10]), .I1(n901), .CO(n39450));
    SB_CARRY add_5712_13 (.CI(n39559), .I0(n13765[10]), .I1(n886_adj_4439), 
            .CO(n39560));
    SB_LUT4 add_5712_12_lut (.I0(GND_net), .I1(n13765[9]), .I2(n813_adj_4441), 
            .I3(n39558), .O(n12924[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5888_12_lut (.I0(GND_net), .I1(n16845[9]), .I2(n828), 
            .I3(n39448), .O(n16365[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5888_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_6 (.CI(n39259), .I0(GND_net), .I1(n1_adj_4767[4]), 
            .CO(n39260));
    SB_LUT4 i35594_3_lut (.I0(n6_adj_4440), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n21_adj_4407), .I3(GND_net), .O(n50547));   // verilog/motorControl.v(31[38:63])
    defparam i35594_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6013_5 (.CI(n39352), .I0(n18425[2]), .I1(n332), .CO(n39353));
    SB_LUT4 i35595_3_lut (.I0(n50547), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n23_adj_4417), .I3(GND_net), .O(n50548));   // verilog/motorControl.v(31[38:63])
    defparam i35595_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_6013_4_lut (.I0(GND_net), .I1(n18425[1]), .I2(n259), .I3(n39351), 
            .O(n18205[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6013_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34892_4_lut (.I0(n43), .I1(n25_adj_4416), .I2(n23_adj_4417), 
            .I3(n49866), .O(n49844));
    defparam i34892_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35530_4_lut (.I0(n24_adj_4413), .I1(n8_adj_4412), .I2(n45), 
            .I3(n49842), .O(n50483));   // verilog/motorControl.v(31[38:63])
    defparam i35530_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35525_3_lut (.I0(n50548), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n25_adj_4416), .I3(GND_net), .O(n50478));   // verilog/motorControl.v(31[38:63])
    defparam i35525_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34894_4_lut (.I0(n43), .I1(n41), .I2(n39), .I3(n50605), 
            .O(n49846));
    defparam i34894_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35616_4_lut (.I0(n50478), .I1(n50483), .I2(n45), .I3(n49844), 
            .O(n50569));   // verilog/motorControl.v(31[38:63])
    defparam i35616_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35685_3_lut (.I0(n50652), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n41), .I3(GND_net), .O(n40));   // verilog/motorControl.v(31[38:63])
    defparam i35685_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35618_4_lut (.I0(n40), .I1(n50569), .I2(n45), .I3(n49846), 
            .O(n50571));   // verilog/motorControl.v(31[38:63])
    defparam i35618_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 IntegralLimit_23__I_0_i4_4_lut (.I0(\PID_CONTROLLER.integral [0]), 
            .I1(IntegralLimit[1]), .I2(\PID_CONTROLLER.integral [1]), .I3(IntegralLimit[0]), 
            .O(n4_adj_4442));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i35598_3_lut (.I0(n4_adj_4442), .I1(IntegralLimit[13]), .I2(\PID_CONTROLLER.integral [13]), 
            .I3(GND_net), .O(n50551));   // verilog/motorControl.v(31[10:34])
    defparam i35598_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35599_3_lut (.I0(n50551), .I1(IntegralLimit[14]), .I2(\PID_CONTROLLER.integral [14]), 
            .I3(GND_net), .O(n50552));   // verilog/motorControl.v(31[10:34])
    defparam i35599_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 unary_minus_16_add_3_5_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[3]), 
            .I3(n39258), .O(n257[3])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i34947_4_lut (.I0(\PID_CONTROLLER.integral [16]), .I1(n51853), 
            .I2(IntegralLimit[16]), .I3(n50199), .O(n49899));
    defparam i34947_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 i35670_4_lut (.I0(n30), .I1(n10_adj_4422), .I2(n51877), .I3(n49893), 
            .O(n50623));   // verilog/motorControl.v(31[10:34])
    defparam i35670_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35519_3_lut (.I0(n50552), .I1(IntegralLimit[15]), .I2(\PID_CONTROLLER.integral [15]), 
            .I3(GND_net), .O(n50472));   // verilog/motorControl.v(31[10:34])
    defparam i35519_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35712_4_lut (.I0(n50472), .I1(n50623), .I2(n51877), .I3(n49899), 
            .O(n50665));   // verilog/motorControl.v(31[10:34])
    defparam i35712_4_lut.LUT_INIT = 16'hccca;
    SB_CARRY add_5712_12 (.CI(n39558), .I0(n13765[9]), .I1(n813_adj_4441), 
            .CO(n39559));
    SB_LUT4 i35713_3_lut (.I0(n50665), .I1(IntegralLimit[18]), .I2(\PID_CONTROLLER.integral [18]), 
            .I3(GND_net), .O(n50666));   // verilog/motorControl.v(31[10:34])
    defparam i35713_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35701_3_lut (.I0(n50666), .I1(IntegralLimit[19]), .I2(\PID_CONTROLLER.integral [19]), 
            .I3(GND_net), .O(n50654));   // verilog/motorControl.v(31[10:34])
    defparam i35701_3_lut.LUT_INIT = 16'h8e8e;
    SB_CARRY unary_minus_16_add_3_5 (.CI(n39258), .I0(GND_net), .I1(n1_adj_4767[3]), 
            .CO(n39259));
    SB_CARRY add_5888_12 (.CI(n39448), .I0(n16845[9]), .I1(n828), .CO(n39449));
    SB_LUT4 i34930_4_lut (.I0(\PID_CONTROLLER.integral [21]), .I1(n51845), 
            .I2(IntegralLimit[21]), .I3(n50633), .O(n49882));
    defparam i34930_4_lut.LUT_INIT = 16'h5a7b;
    SB_LUT4 add_5888_11_lut (.I0(GND_net), .I1(n16845[8]), .I2(n755), 
            .I3(n39447), .O(n16365[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5888_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5873_7_lut (.I0(GND_net), .I1(n16620[4]), .I2(n460), .I3(n39874), 
            .O(n16109[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5873_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6013_4 (.CI(n39351), .I0(n18425[1]), .I1(n259), .CO(n39352));
    SB_LUT4 add_6013_3_lut (.I0(GND_net), .I1(n18425[0]), .I2(n186), .I3(n39350), 
            .O(n18205[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6013_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_4_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[2]), 
            .I3(n39257), .O(n257[2])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 IntegralLimit_23__I_0_i45_rep_170_2_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(IntegralLimit[22]), .I2(GND_net), .I3(GND_net), .O(n51843));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i45_rep_170_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35610_4_lut (.I0(n50470), .I1(n50475), .I2(n51843), .I3(n49880), 
            .O(n50563));   // verilog/motorControl.v(31[10:34])
    defparam i35610_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 add_5712_11_lut (.I0(GND_net), .I1(n13765[8]), .I2(n740_adj_4445), 
            .I3(n39557), .O(n12924[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_4 (.CI(n39257), .I0(GND_net), .I1(n1_adj_4767[2]), 
            .CO(n39258));
    SB_LUT4 i35683_3_lut (.I0(n50654), .I1(IntegralLimit[20]), .I2(\PID_CONTROLLER.integral [20]), 
            .I3(GND_net), .O(n40_adj_4446));   // verilog/motorControl.v(31[10:34])
    defparam i35683_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35619_3_lut (.I0(n50571), .I1(\PID_CONTROLLER.integral_23__N_3623 [23]), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3622 ));   // verilog/motorControl.v(31[38:63])
    defparam i35619_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i35612_4_lut (.I0(n40_adj_4446), .I1(n50563), .I2(n51843), 
            .I3(n49882), .O(n50565));   // verilog/motorControl.v(31[10:34])
    defparam i35612_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 \PID_CONTROLLER.integral_23__I_831_4_lut  (.I0(n50565), .I1(\PID_CONTROLLER.integral_23__N_3622 ), 
            .I2(\PID_CONTROLLER.integral [23]), .I3(IntegralLimit[23]), 
            .O(\PID_CONTROLLER.integral_23__N_3620 ));   // verilog/motorControl.v(31[10:63])
    defparam \PID_CONTROLLER.integral_23__I_831_4_lut .LUT_INIT = 16'h80c8;
    SB_LUT4 add_5322_18_lut (.I0(GND_net), .I1(n13364[15]), .I2(GND_net), 
            .I3(n39990), .O(n12113[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5873_7 (.CI(n39874), .I0(n16620[4]), .I1(n460), .CO(n39875));
    SB_LUT4 add_5873_6_lut (.I0(GND_net), .I1(n16620[3]), .I2(n387), .I3(n39873), 
            .O(n16109[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5873_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5712_11 (.CI(n39557), .I0(n13765[8]), .I1(n740_adj_4445), 
            .CO(n39558));
    SB_CARRY add_6013_3 (.CI(n39350), .I0(n18425[0]), .I1(n186), .CO(n39351));
    SB_CARRY add_5888_11 (.CI(n39447), .I0(n16845[8]), .I1(n755), .CO(n39448));
    SB_LUT4 add_5712_10_lut (.I0(GND_net), .I1(n13765[7]), .I2(n667_adj_4447), 
            .I3(n39556), .O(n12924[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6013_2_lut (.I0(GND_net), .I1(n44_adj_4448), .I2(n113_adj_4449), 
            .I3(GND_net), .O(n18205[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6013_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5712_10 (.CI(n39556), .I0(n13765[7]), .I1(n667_adj_4447), 
            .CO(n39557));
    SB_LUT4 unary_minus_16_add_3_3_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[1]), 
            .I3(n39256), .O(n257[1])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5888_10_lut (.I0(GND_net), .I1(n16845[7]), .I2(n682), 
            .I3(n39446), .O(n16365[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5888_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5873_6 (.CI(n39873), .I0(n16620[3]), .I1(n387), .CO(n39874));
    SB_CARRY add_5322_18 (.CI(n39990), .I0(n13364[15]), .I1(GND_net), 
            .CO(n39991));
    SB_LUT4 i20684_2_lut (.I0(n1[23]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[23]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20684_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5712_9_lut (.I0(GND_net), .I1(n13765[6]), .I2(n594_adj_4452), 
            .I3(n39555), .O(n12924[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i126_2_lut (.I0(\Kp[2] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n186_adj_4453));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i126_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i263_2_lut (.I0(\Kp[5] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n390));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i8_1_lut (.I0(IntegralLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[7]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i181_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n268_adj_4455));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5322_17_lut (.I0(GND_net), .I1(n13364[14]), .I2(GND_net), 
            .I3(n39989), .O(n12113[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6013_2 (.CI(GND_net), .I0(n44_adj_4448), .I1(n113_adj_4449), 
            .CO(n39350));
    SB_LUT4 mult_10_i104_2_lut (.I0(\Kp[2] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n153_adj_4456));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i104_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5322_17 (.CI(n39989), .I0(n13364[14]), .I1(GND_net), 
            .CO(n39990));
    SB_LUT4 mult_11_i265_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n393_adj_4457));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i265_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5712_9 (.CI(n39555), .I0(n13765[6]), .I1(n594_adj_4452), 
            .CO(n39556));
    SB_LUT4 mult_11_i230_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n341));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i230_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5888_10 (.CI(n39446), .I0(n16845[7]), .I1(n682), .CO(n39447));
    SB_LUT4 add_5712_8_lut (.I0(GND_net), .I1(n13765[5]), .I2(n521_adj_4458), 
            .I3(n39554), .O(n12924[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_3 (.CI(n39256), .I0(GND_net), .I1(n1_adj_4767[1]), 
            .CO(n39257));
    SB_LUT4 mult_10_i153_2_lut (.I0(\Kp[3] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n226_adj_4459));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i153_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5712_8 (.CI(n39554), .I0(n13765[5]), .I1(n521_adj_4458), 
            .CO(n39555));
    SB_LUT4 add_6032_10_lut (.I0(GND_net), .I1(n18605[7]), .I2(n700), 
            .I3(n39349), .O(n18425[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6032_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i314_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n466_adj_4460));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i314_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5873_5_lut (.I0(GND_net), .I1(n16620[2]), .I2(n314), .I3(n39872), 
            .O(n16109[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5873_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i312_2_lut (.I0(\Kp[6] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n463));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6032_9_lut (.I0(GND_net), .I1(n18605[6]), .I2(n627), .I3(n39348), 
            .O(n18425[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6032_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5888_9_lut (.I0(GND_net), .I1(n16845[6]), .I2(n609), .I3(n39445), 
            .O(n16365[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5888_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5888_9 (.CI(n39445), .I0(n16845[6]), .I1(n609), .CO(n39446));
    SB_CARRY add_5873_5 (.CI(n39872), .I0(n16620[2]), .I1(n314), .CO(n39873));
    SB_LUT4 add_5888_8_lut (.I0(GND_net), .I1(n16845[5]), .I2(n536), .I3(n39444), 
            .O(n16365[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5888_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i9_1_lut (.I0(IntegralLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[8]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i279_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n414));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i279_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6032_9 (.CI(n39348), .I0(n18605[6]), .I1(n627), .CO(n39349));
    SB_LUT4 add_6032_8_lut (.I0(GND_net), .I1(n18605[5]), .I2(n554), .I3(n39347), 
            .O(n18425[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6032_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5888_8 (.CI(n39444), .I0(n16845[5]), .I1(n536), .CO(n39445));
    SB_LUT4 unary_minus_16_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[0]), 
            .I3(VCC_net), .O(n257[0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5712_7_lut (.I0(GND_net), .I1(n13765[4]), .I2(n448_adj_4463), 
            .I3(n39553), .O(n12924[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i10_1_lut (.I0(IntegralLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[9]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i363_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n539_adj_4465));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i363_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i11_1_lut (.I0(IntegralLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[10]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5322_16_lut (.I0(GND_net), .I1(n13364[13]), .I2(n1102_adj_4467), 
            .I3(n39988), .O(n12113[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5322_16 (.CI(n39988), .I0(n13364[13]), .I1(n1102_adj_4467), 
            .CO(n39989));
    SB_LUT4 mult_11_i328_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n487));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i361_2_lut (.I0(\Kp[7] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n536_adj_4468));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i361_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6032_8 (.CI(n39347), .I0(n18605[5]), .I1(n554), .CO(n39348));
    SB_LUT4 add_5322_15_lut (.I0(GND_net), .I1(n13364[12]), .I2(n1029_adj_4469), 
            .I3(n39987), .O(n12113[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4767[0]), 
            .CO(n39256));
    SB_CARRY add_5712_7 (.CI(n39553), .I0(n13765[4]), .I1(n448_adj_4463), 
            .CO(n39554));
    SB_LUT4 add_5712_6_lut (.I0(GND_net), .I1(n13765[3]), .I2(n375), .I3(n39552), 
            .O(n12924[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i202_2_lut (.I0(\Kp[4] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n299));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i202_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5712_6 (.CI(n39552), .I0(n13765[3]), .I1(n375), .CO(n39553));
    SB_LUT4 add_5888_7_lut (.I0(GND_net), .I1(n16845[4]), .I2(n463_adj_4470), 
            .I3(n39443), .O(n16365[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5888_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i12_1_lut (.I0(IntegralLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[11]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i377_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n560));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i377_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5888_7 (.CI(n39443), .I0(n16845[4]), .I1(n463_adj_4470), 
            .CO(n39444));
    SB_LUT4 add_6032_7_lut (.I0(GND_net), .I1(n18605[4]), .I2(n481), .I3(n39346), 
            .O(n18425[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6032_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5873_4_lut (.I0(GND_net), .I1(n16620[1]), .I2(n241_adj_4472), 
            .I3(n39871), .O(n16109[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5873_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4768[23]), 
            .I3(n39255), .O(\PID_CONTROLLER.integral_23__N_3623 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i412_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n612_adj_4474));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i412_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i175_2_lut (.I0(\Kp[3] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n259_adj_4475));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i81_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n119_adj_4476));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i34_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [16]), 
            .I2(GND_net), .I3(GND_net), .O(n50_adj_4477));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i461_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n685_adj_4478));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i461_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i251_2_lut (.I0(\Kp[5] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n372));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i224_2_lut (.I0(\Kp[4] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n332_adj_4479));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i300_2_lut (.I0(\Kp[6] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n445));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i300_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6032_7 (.CI(n39346), .I0(n18605[4]), .I1(n481), .CO(n39347));
    SB_LUT4 add_5712_5_lut (.I0(GND_net), .I1(n13765[2]), .I2(n302), .I3(n39551), 
            .O(n12924[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5322_15 (.CI(n39987), .I0(n13364[12]), .I1(n1029_adj_4469), 
            .CO(n39988));
    SB_LUT4 unary_minus_5_inv_0_i13_1_lut (.I0(IntegralLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[12]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5873_4 (.CI(n39871), .I0(n16620[1]), .I1(n241_adj_4472), 
            .CO(n39872));
    SB_LUT4 unary_minus_5_add_3_24_lut (.I0(\PID_CONTROLLER.integral [22]), 
            .I1(GND_net), .I2(n1_adj_4768[22]), .I3(n39254), .O(n45)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i130_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n192_adj_4482));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5322_14_lut (.I0(GND_net), .I1(n13364[11]), .I2(n956_adj_4483), 
            .I3(n39986), .O(n12113[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i410_2_lut (.I0(\Kp[8] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n609_adj_4484));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5873_3_lut (.I0(GND_net), .I1(n16620[0]), .I2(n168_adj_4485), 
            .I3(n39870), .O(n16109[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5873_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5712_5 (.CI(n39551), .I0(n13765[2]), .I1(n302), .CO(n39552));
    SB_LUT4 add_6032_6_lut (.I0(GND_net), .I1(n18605[3]), .I2(n408), .I3(n39345), 
            .O(n18425[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6032_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5712_4_lut (.I0(GND_net), .I1(n13765[1]), .I2(n229), .I3(n39550), 
            .O(n12924[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_24 (.CI(n39254), .I0(GND_net), .I1(n1_adj_4768[22]), 
            .CO(n39255));
    SB_LUT4 unary_minus_5_add_3_23_lut (.I0(\PID_CONTROLLER.integral [21]), 
            .I1(GND_net), .I2(n1_adj_4768[21]), .I3(n39253), .O(n43)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_23_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5888_6_lut (.I0(GND_net), .I1(n16845[3]), .I2(n390_adj_4487), 
            .I3(n39442), .O(n16365[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5888_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5322_14 (.CI(n39986), .I0(n13364[11]), .I1(n956_adj_4483), 
            .CO(n39987));
    SB_CARRY add_5888_6 (.CI(n39442), .I0(n16845[3]), .I1(n390_adj_4487), 
            .CO(n39443));
    SB_LUT4 add_5322_13_lut (.I0(GND_net), .I1(n13364[10]), .I2(n883_adj_4488), 
            .I3(n39985), .O(n12113[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5322_13 (.CI(n39985), .I0(n13364[10]), .I1(n883_adj_4488), 
            .CO(n39986));
    SB_LUT4 add_5322_12_lut (.I0(GND_net), .I1(n13364[9]), .I2(n810_adj_4489), 
            .I3(n39984), .O(n12113[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5712_4 (.CI(n39550), .I0(n13765[1]), .I1(n229), .CO(n39551));
    SB_LUT4 mult_10_i349_2_lut (.I0(\Kp[7] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n518));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i273_2_lut (.I0(\Kp[5] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n405_adj_4490));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i273_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i510_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n758_adj_4491));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i510_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5873_3 (.CI(n39870), .I0(n16620[0]), .I1(n168_adj_4485), 
            .CO(n39871));
    SB_LUT4 mult_10_i459_2_lut (.I0(\Kp[9] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n682_adj_4492));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i179_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n265_adj_4493));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5888_5_lut (.I0(GND_net), .I1(n16845[2]), .I2(n317_adj_4494), 
            .I3(n39441), .O(n16365[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5888_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i14_1_lut (.I0(IntegralLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[13]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5873_2_lut (.I0(GND_net), .I1(n26_adj_4496), .I2(n95_adj_4497), 
            .I3(GND_net), .O(n16109[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5873_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5712_3_lut (.I0(GND_net), .I1(n13765[0]), .I2(n156), .I3(n39549), 
            .O(n12924[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6032_6 (.CI(n39345), .I0(n18605[3]), .I1(n408), .CO(n39346));
    SB_CARRY add_5322_12 (.CI(n39984), .I0(n13364[9]), .I1(n810_adj_4489), 
            .CO(n39985));
    SB_CARRY add_5873_2 (.CI(GND_net), .I0(n26_adj_4496), .I1(n95_adj_4497), 
            .CO(n39870));
    SB_LUT4 add_5322_11_lut (.I0(GND_net), .I1(n13364[8]), .I2(n737_adj_4498), 
            .I3(n39983), .O(n12113[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5888_5 (.CI(n39441), .I0(n16845[2]), .I1(n317_adj_4494), 
            .CO(n39442));
    SB_CARRY add_5322_11 (.CI(n39983), .I0(n13364[8]), .I1(n737_adj_4498), 
            .CO(n39984));
    SB_LUT4 add_5903_16_lut (.I0(GND_net), .I1(n17069[13]), .I2(n1120_adj_4499), 
            .I3(n39869), .O(n16620[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5903_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6032_5_lut (.I0(GND_net), .I1(n18605[2]), .I2(n335), .I3(n39344), 
            .O(n18425[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6032_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5903_15_lut (.I0(GND_net), .I1(n17069[12]), .I2(n1047_adj_4500), 
            .I3(n39868), .O(n16620[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5903_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_23 (.CI(n39253), .I0(GND_net), .I1(n1_adj_4768[21]), 
            .CO(n39254));
    SB_CARRY add_5903_15 (.CI(n39868), .I0(n17069[12]), .I1(n1047_adj_4500), 
            .CO(n39869));
    SB_LUT4 unary_minus_5_add_3_22_lut (.I0(\PID_CONTROLLER.integral [20]), 
            .I1(GND_net), .I2(n1_adj_4768[20]), .I3(n39252), .O(n41)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_22_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6032_5 (.CI(n39344), .I0(n18605[2]), .I1(n335), .CO(n39345));
    SB_LUT4 add_5888_4_lut (.I0(GND_net), .I1(n16845[1]), .I2(n244_adj_4502), 
            .I3(n39440), .O(n16365[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5888_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5322_10_lut (.I0(GND_net), .I1(n13364[7]), .I2(n664_adj_4503), 
            .I3(n39982), .O(n12113[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5712_3 (.CI(n39549), .I0(n13765[0]), .I1(n156), .CO(n39550));
    SB_CARRY unary_minus_5_add_3_22 (.CI(n39252), .I0(GND_net), .I1(n1_adj_4768[20]), 
            .CO(n39253));
    SB_LUT4 add_6032_4_lut (.I0(GND_net), .I1(n18605[1]), .I2(n262), .I3(n39343), 
            .O(n18425[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6032_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5888_4 (.CI(n39440), .I0(n16845[1]), .I1(n244_adj_4502), 
            .CO(n39441));
    SB_LUT4 add_5712_2_lut (.I0(GND_net), .I1(n14_adj_4504), .I2(n83), 
            .I3(GND_net), .O(n12924[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5712_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i232_2_lut (.I0(\Kp[4] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n344_adj_4505));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i232_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5888_3_lut (.I0(GND_net), .I1(n16845[0]), .I2(n171_adj_4506), 
            .I3(n39439), .O(n16365[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5888_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6032_4 (.CI(n39343), .I0(n18605[1]), .I1(n262), .CO(n39344));
    SB_LUT4 add_6032_3_lut (.I0(GND_net), .I1(n18605[0]), .I2(n189), .I3(n39342), 
            .O(n18425[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6032_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_21_lut (.I0(\PID_CONTROLLER.integral [19]), 
            .I1(GND_net), .I2(n1_adj_4768[19]), .I3(n39251), .O(n39)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_21_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_21 (.CI(n39251), .I0(GND_net), .I1(n1_adj_4768[19]), 
            .CO(n39252));
    SB_CARRY add_6032_3 (.CI(n39342), .I0(n18605[0]), .I1(n189), .CO(n39343));
    SB_CARRY add_5712_2 (.CI(GND_net), .I0(n14_adj_4504), .I1(n83), .CO(n39549));
    SB_LUT4 mult_11_i651_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n968_adj_4508));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i651_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i700_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1041_adj_4509));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i700_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5322_10 (.CI(n39982), .I0(n13364[7]), .I1(n664_adj_4503), 
            .CO(n39983));
    SB_LUT4 unary_minus_5_add_3_20_lut (.I0(\PID_CONTROLLER.integral [18]), 
            .I1(GND_net), .I2(n1_adj_4768[18]), .I3(n39250), .O(n37)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_20_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i592_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n880));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6023_11_lut (.I0(GND_net), .I1(n18524[8]), .I2(n770_adj_4511), 
            .I3(n39548), .O(n18325[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6023_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i641_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n953));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6023_10_lut (.I0(GND_net), .I1(n18524[7]), .I2(n697_adj_4512), 
            .I3(n39547), .O(n18325[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6023_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i502_2_lut (.I0(\Kp[10] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n746));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i502_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5888_3 (.CI(n39439), .I0(n16845[0]), .I1(n171_adj_4506), 
            .CO(n39440));
    SB_LUT4 mult_10_i551_2_lut (.I0(\Kp[11] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n819));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i600_2_lut (.I0(\Kp[12] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n892));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i690_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1026));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i281_2_lut (.I0(\Kp[5] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n417_adj_4513));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i281_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6032_2_lut (.I0(GND_net), .I1(n47), .I2(n116), .I3(GND_net), 
            .O(n18425[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6032_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut_adj_1524 (.I0(n6_adj_4514), .I1(\Kp[4] ), .I2(n19029[2]), 
            .I3(n1[18]), .O(n18980[3]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1524.LUT_INIT = 16'h965a;
    SB_CARRY add_6032_2 (.CI(GND_net), .I0(n47), .I1(n116), .CO(n39342));
    SB_CARRY add_6023_10 (.CI(n39547), .I0(n18524[7]), .I1(n697_adj_4512), 
            .CO(n39548));
    SB_CARRY unary_minus_5_add_3_20 (.CI(n39250), .I0(GND_net), .I1(n1_adj_4768[18]), 
            .CO(n39251));
    SB_LUT4 add_5903_14_lut (.I0(GND_net), .I1(n17069[11]), .I2(n974_adj_4515), 
            .I3(n39867), .O(n16620[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5903_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5888_2_lut (.I0(GND_net), .I1(n29_adj_4516), .I2(n98_adj_4517), 
            .I3(GND_net), .O(n16365[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5888_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6049_9_lut (.I0(GND_net), .I1(n18749[6]), .I2(n630_adj_4518), 
            .I3(n39341), .O(n18605[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6049_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6049_8_lut (.I0(GND_net), .I1(n18749[5]), .I2(n557_adj_4519), 
            .I3(n39340), .O(n18605[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6049_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5888_2 (.CI(GND_net), .I0(n29_adj_4516), .I1(n98_adj_4517), 
            .CO(n39439));
    SB_LUT4 i25760_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n19077[0]));   // verilog/motorControl.v(34[16:22])
    defparam i25760_4_lut.LUT_INIT = 16'h6ca0;
    SB_LUT4 add_5322_9_lut (.I0(GND_net), .I1(n13364[6]), .I2(n591_adj_4520), 
            .I3(n39981), .O(n12113[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6049_8 (.CI(n39340), .I0(n18749[5]), .I1(n557_adj_4519), 
            .CO(n39341));
    SB_CARRY add_5903_14 (.CI(n39867), .I0(n17069[11]), .I1(n974_adj_4515), 
            .CO(n39868));
    SB_LUT4 add_5903_13_lut (.I0(GND_net), .I1(n17069[10]), .I2(n901_adj_4521), 
            .I3(n39866), .O(n16620[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5903_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_19_lut (.I0(\PID_CONTROLLER.integral [17]), 
            .I1(GND_net), .I2(n1_adj_4768[17]), .I3(n39249), .O(n35)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_19_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5322_9 (.CI(n39981), .I0(n13364[6]), .I1(n591_adj_4520), 
            .CO(n39982));
    SB_LUT4 add_6023_9_lut (.I0(GND_net), .I1(n18524[6]), .I2(n624_adj_4523), 
            .I3(n39546), .O(n18325[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6023_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6023_9 (.CI(n39546), .I0(n18524[6]), .I1(n624_adj_4523), 
            .CO(n39547));
    SB_LUT4 i2_4_lut_adj_1525 (.I0(n4_adj_4524), .I1(\Kp[3] ), .I2(n19060[1]), 
            .I3(n1[19]), .O(n19029[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1525.LUT_INIT = 16'h965a;
    SB_CARRY unary_minus_5_add_3_19 (.CI(n39249), .I0(GND_net), .I1(n1_adj_4768[17]), 
            .CO(n39250));
    SB_LUT4 mult_10_i330_2_lut (.I0(\Kp[6] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n490_adj_4525));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i330_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1526 (.I0(\Kp[0] ), .I1(\Kp[3] ), .I2(n1[23]), 
            .I3(n1[20]), .O(n12_adj_4526));   // verilog/motorControl.v(34[16:22])
    defparam i2_4_lut_adj_1526.LUT_INIT = 16'h9c50;
    SB_CARRY add_5903_13 (.CI(n39866), .I0(n17069[10]), .I1(n901_adj_4521), 
            .CO(n39867));
    SB_LUT4 add_5917_15_lut (.I0(GND_net), .I1(n17265[12]), .I2(n1050_adj_4527), 
            .I3(n39438), .O(n16845[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5917_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25928_4_lut (.I0(n19029[2]), .I1(\Kp[4] ), .I2(n6_adj_4514), 
            .I3(n1[18]), .O(n8_adj_4528));   // verilog/motorControl.v(34[16:22])
    defparam i25928_4_lut.LUT_INIT = 16'he8a0;
    SB_LUT4 add_6049_7_lut (.I0(GND_net), .I1(n18749[4]), .I2(n484_adj_4529), 
            .I3(n39339), .O(n18605[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6049_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5917_14_lut (.I0(GND_net), .I1(n17265[11]), .I2(n977_adj_4530), 
            .I3(n39437), .O(n16845[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5917_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6023_8_lut (.I0(GND_net), .I1(n18524[5]), .I2(n551_adj_4531), 
            .I3(n39545), .O(n18325[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6023_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6049_7 (.CI(n39339), .I0(n18749[4]), .I1(n484_adj_4529), 
            .CO(n39340));
    SB_CARRY add_5917_14 (.CI(n39437), .I0(n17265[11]), .I1(n977_adj_4530), 
            .CO(n39438));
    SB_LUT4 add_6049_6_lut (.I0(GND_net), .I1(n18749[3]), .I2(n411_adj_4532), 
            .I3(n39338), .O(n18605[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6049_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_18_lut (.I0(\PID_CONTROLLER.integral [16]), 
            .I1(GND_net), .I2(n1_adj_4768[16]), .I3(n39248), .O(n33)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_18_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_18 (.CI(n39248), .I0(GND_net), .I1(n1_adj_4768[16]), 
            .CO(n39249));
    SB_DFF \PID_CONTROLLER.integral_i23  (.Q(\PID_CONTROLLER.integral [23]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 i1_4_lut_adj_1527 (.I0(\Kp[4] ), .I1(\Kp[2] ), .I2(n1[19]), 
            .I3(n1[21]), .O(n11_adj_4534));   // verilog/motorControl.v(34[16:22])
    defparam i1_4_lut_adj_1527.LUT_INIT = 16'h6ca0;
    SB_DFF \PID_CONTROLLER.integral_i22  (.Q(\PID_CONTROLLER.integral [22]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i21  (.Q(\PID_CONTROLLER.integral [21]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i20  (.Q(\PID_CONTROLLER.integral [20]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i19  (.Q(\PID_CONTROLLER.integral [19]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i18  (.Q(\PID_CONTROLLER.integral [18]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i17  (.Q(\PID_CONTROLLER.integral [17]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i16  (.Q(\PID_CONTROLLER.integral [16]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i15  (.Q(\PID_CONTROLLER.integral [15]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i14  (.Q(\PID_CONTROLLER.integral [14]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i13  (.Q(\PID_CONTROLLER.integral [13]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i12  (.Q(\PID_CONTROLLER.integral [12]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_5917_13_lut (.I0(GND_net), .I1(n17265[10]), .I2(n904_adj_4535), 
            .I3(n39436), .O(n16845[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5917_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF \PID_CONTROLLER.integral_i11  (.Q(\PID_CONTROLLER.integral [11]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i10  (.Q(\PID_CONTROLLER.integral [10]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i9  (.Q(\PID_CONTROLLER.integral [9]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i8  (.Q(\PID_CONTROLLER.integral [8]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i7  (.Q(\PID_CONTROLLER.integral [7]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i6  (.Q(\PID_CONTROLLER.integral [6]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i5  (.Q(\PID_CONTROLLER.integral [5]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i4  (.Q(\PID_CONTROLLER.integral [4]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i3  (.Q(\PID_CONTROLLER.integral [3]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i2  (.Q(\PID_CONTROLLER.integral [2]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF \PID_CONTROLLER.integral_i1  (.Q(\PID_CONTROLLER.integral [1]), 
           .C(clk32MHz), .D(\PID_CONTROLLER.integral_23__N_3572 [1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i23 (.Q(duty[23]), .C(clk32MHz), .D(duty_23__N_3548[23]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i22 (.Q(duty[22]), .C(clk32MHz), .D(duty_23__N_3548[22]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i21 (.Q(duty[21]), .C(clk32MHz), .D(duty_23__N_3548[21]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i20 (.Q(duty[20]), .C(clk32MHz), .D(duty_23__N_3548[20]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i19 (.Q(duty[19]), .C(clk32MHz), .D(duty_23__N_3548[19]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i18 (.Q(duty[18]), .C(clk32MHz), .D(duty_23__N_3548[18]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i17 (.Q(duty[17]), .C(clk32MHz), .D(duty_23__N_3548[17]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i16 (.Q(duty[16]), .C(clk32MHz), .D(duty_23__N_3548[16]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i15 (.Q(duty[15]), .C(clk32MHz), .D(duty_23__N_3548[15]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i14 (.Q(duty[14]), .C(clk32MHz), .D(duty_23__N_3548[14]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i13 (.Q(duty[13]), .C(clk32MHz), .D(duty_23__N_3548[13]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i12 (.Q(duty[12]), .C(clk32MHz), .D(duty_23__N_3548[12]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i11 (.Q(duty[11]), .C(clk32MHz), .D(duty_23__N_3548[11]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i10 (.Q(duty[10]), .C(clk32MHz), .D(duty_23__N_3548[10]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i9 (.Q(duty[9]), .C(clk32MHz), .D(duty_23__N_3548[9]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i8 (.Q(duty[8]), .C(clk32MHz), .D(duty_23__N_3548[8]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_5917_13 (.CI(n39436), .I0(n17265[10]), .I1(n904_adj_4535), 
            .CO(n39437));
    SB_DFF result_i7 (.Q(duty[7]), .C(clk32MHz), .D(duty_23__N_3548[7]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i6 (.Q(duty[6]), .C(clk32MHz), .D(duty_23__N_3548[6]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i5 (.Q(duty[5]), .C(clk32MHz), .D(duty_23__N_3548[5]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i4 (.Q(duty[4]), .C(clk32MHz), .D(duty_23__N_3548[4]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i3 (.Q(duty[3]), .C(clk32MHz), .D(duty_23__N_3548[3]));   // verilog/motorControl.v(29[14] 48[8])
    SB_DFF result_i2 (.Q(duty[2]), .C(clk32MHz), .D(duty_23__N_3548[2]));   // verilog/motorControl.v(29[14] 48[8])
    SB_LUT4 add_5917_12_lut (.I0(GND_net), .I1(n17265[9]), .I2(n831_adj_4536), 
            .I3(n39435), .O(n16845[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5917_12_lut.LUT_INIT = 16'hC33C;
    SB_DFF result_i1 (.Q(duty[1]), .C(clk32MHz), .D(duty_23__N_3548[1]));   // verilog/motorControl.v(29[14] 48[8])
    SB_CARRY add_6049_6 (.CI(n39338), .I0(n18749[3]), .I1(n411_adj_4532), 
            .CO(n39339));
    SB_LUT4 unary_minus_5_add_3_17_lut (.I0(\PID_CONTROLLER.integral [15]), 
            .I1(GND_net), .I2(n1_adj_4768[15]), .I3(n39247), .O(n31)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_17_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6049_5_lut (.I0(GND_net), .I1(n18749[2]), .I2(n338_adj_4538), 
            .I3(n39337), .O(n18605[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6049_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_17 (.CI(n39247), .I0(GND_net), .I1(n1_adj_4768[15]), 
            .CO(n39248));
    SB_CARRY add_6049_5 (.CI(n39337), .I0(n18749[2]), .I1(n338_adj_4538), 
            .CO(n39338));
    SB_LUT4 add_5903_12_lut (.I0(GND_net), .I1(n17069[9]), .I2(n828_adj_4539), 
            .I3(n39865), .O(n16620[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5903_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5903_12 (.CI(n39865), .I0(n17069[9]), .I1(n828_adj_4539), 
            .CO(n39866));
    SB_LUT4 add_5903_11_lut (.I0(GND_net), .I1(n17069[8]), .I2(n755_adj_4540), 
            .I3(n39864), .O(n16620[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5903_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_16_lut (.I0(\PID_CONTROLLER.integral [14]), 
            .I1(GND_net), .I2(n1_adj_4768[14]), .I3(n39246), .O(n29_adj_4418)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_16_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6023_8 (.CI(n39545), .I0(n18524[5]), .I1(n551_adj_4531), 
            .CO(n39546));
    SB_LUT4 i25889_4_lut (.I0(n19060[1]), .I1(\Kp[3] ), .I2(n4_adj_4524), 
            .I3(n1[19]), .O(n6_adj_4542));   // verilog/motorControl.v(34[16:22])
    defparam i25889_4_lut.LUT_INIT = 16'he8a0;
    SB_CARRY unary_minus_5_add_3_16 (.CI(n39246), .I0(GND_net), .I1(n1_adj_4768[14]), 
            .CO(n39247));
    SB_LUT4 add_6023_7_lut (.I0(GND_net), .I1(n18524[4]), .I2(n478_adj_4543), 
            .I3(n39544), .O(n18325[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6023_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5903_11 (.CI(n39864), .I0(n17069[8]), .I1(n755_adj_4540), 
            .CO(n39865));
    SB_CARRY add_5917_12 (.CI(n39435), .I0(n17265[9]), .I1(n831_adj_4536), 
            .CO(n39436));
    SB_CARRY add_6023_7 (.CI(n39544), .I0(n18524[4]), .I1(n478_adj_4543), 
            .CO(n39545));
    SB_LUT4 unary_minus_5_add_3_15_lut (.I0(\PID_CONTROLLER.integral [13]), 
            .I1(GND_net), .I2(n1_adj_4768[13]), .I3(n39245), .O(n27)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_15_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6049_4_lut (.I0(GND_net), .I1(n18749[1]), .I2(n265_adj_4493), 
            .I3(n39336), .O(n18605[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6049_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6049_4 (.CI(n39336), .I0(n18749[1]), .I1(n265_adj_4493), 
            .CO(n39337));
    SB_LUT4 add_5903_10_lut (.I0(GND_net), .I1(n17069[7]), .I2(n682_adj_4492), 
            .I3(n39863), .O(n16620[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5903_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_15 (.CI(n39245), .I0(GND_net), .I1(n1_adj_4768[13]), 
            .CO(n39246));
    SB_CARRY add_5903_10 (.CI(n39863), .I0(n17069[7]), .I1(n682_adj_4492), 
            .CO(n39864));
    SB_LUT4 add_5917_11_lut (.I0(GND_net), .I1(n17265[8]), .I2(n758_adj_4491), 
            .I3(n39434), .O(n16845[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5917_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6023_6_lut (.I0(GND_net), .I1(n18524[3]), .I2(n405_adj_4490), 
            .I3(n39543), .O(n18325[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6023_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5322_8_lut (.I0(GND_net), .I1(n13364[5]), .I2(n518), .I3(n39980), 
            .O(n12113[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5903_9_lut (.I0(GND_net), .I1(n17069[6]), .I2(n609_adj_4484), 
            .I3(n39862), .O(n16620[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5903_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5322_8 (.CI(n39980), .I0(n13364[5]), .I1(n518), .CO(n39981));
    SB_LUT4 add_6049_3_lut (.I0(GND_net), .I1(n18749[0]), .I2(n192_adj_4482), 
            .I3(n39335), .O(n18605[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6049_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i25762_4_lut (.I0(\Kp[0] ), .I1(\Kp[1] ), .I2(n1[22]), .I3(n1[21]), 
            .O(n38783));   // verilog/motorControl.v(34[16:22])
    defparam i25762_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i8_4_lut_adj_1528 (.I0(n6_adj_4542), .I1(n11_adj_4534), .I2(n8_adj_4528), 
            .I3(n12_adj_4526), .O(n18_adj_4544));   // verilog/motorControl.v(34[16:22])
    defparam i8_4_lut_adj_1528.LUT_INIT = 16'h6996;
    SB_CARRY add_5917_11 (.CI(n39434), .I0(n17265[8]), .I1(n758_adj_4491), 
            .CO(n39435));
    SB_LUT4 i3_4_lut_adj_1529 (.I0(\Kp[5] ), .I1(\Kp[1] ), .I2(n1[18]), 
            .I3(n1[22]), .O(n13_adj_4545));   // verilog/motorControl.v(34[16:22])
    defparam i3_4_lut_adj_1529.LUT_INIT = 16'h6ca0;
    SB_CARRY add_6023_6 (.CI(n39543), .I0(n18524[3]), .I1(n405_adj_4490), 
            .CO(n39544));
    SB_LUT4 unary_minus_5_add_3_14_lut (.I0(\PID_CONTROLLER.integral [12]), 
            .I1(GND_net), .I2(n1_adj_4768[12]), .I3(n39244), .O(n25_adj_4416)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_14_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_5903_9 (.CI(n39862), .I0(n17069[6]), .I1(n609_adj_4484), 
            .CO(n39863));
    SB_LUT4 i9_4_lut_adj_1530 (.I0(n13_adj_4545), .I1(n18_adj_4544), .I2(n38783), 
            .I3(n4_adj_4546), .O(n46504));   // verilog/motorControl.v(34[16:22])
    defparam i9_4_lut_adj_1530.LUT_INIT = 16'h6996;
    SB_LUT4 add_5322_7_lut (.I0(GND_net), .I1(n13364[4]), .I2(n445), .I3(n39979), 
            .O(n12113[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5322_7 (.CI(n39979), .I0(n13364[4]), .I1(n445), .CO(n39980));
    SB_CARRY add_6049_3 (.CI(n39335), .I0(n18749[0]), .I1(n192_adj_4482), 
            .CO(n39336));
    SB_LUT4 mult_10_i649_2_lut (.I0(\Kp[13] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n965));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i739_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n1099));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6023_5_lut (.I0(GND_net), .I1(n18524[2]), .I2(n332_adj_4479), 
            .I3(n39542), .O(n18325[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6023_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6023_5 (.CI(n39542), .I0(n18524[2]), .I1(n332_adj_4479), 
            .CO(n39543));
    SB_LUT4 add_5322_6_lut (.I0(GND_net), .I1(n13364[3]), .I2(n372), .I3(n39978), 
            .O(n12113[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5917_10_lut (.I0(GND_net), .I1(n17265[7]), .I2(n685_adj_4478), 
            .I3(n39433), .O(n16845[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5917_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6049_2_lut (.I0(GND_net), .I1(n50_adj_4477), .I2(n119_adj_4476), 
            .I3(GND_net), .O(n18605[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6049_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_14 (.CI(n39244), .I0(GND_net), .I1(n1_adj_4768[12]), 
            .CO(n39245));
    SB_CARRY add_5917_10 (.CI(n39433), .I0(n17265[7]), .I1(n685_adj_4478), 
            .CO(n39434));
    SB_LUT4 add_6023_4_lut (.I0(GND_net), .I1(n18524[1]), .I2(n259_adj_4475), 
            .I3(n39541), .O(n18325[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6023_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5322_6 (.CI(n39978), .I0(n13364[3]), .I1(n372), .CO(n39979));
    SB_LUT4 add_5917_9_lut (.I0(GND_net), .I1(n17265[6]), .I2(n612_adj_4474), 
            .I3(n39432), .O(n16845[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5917_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6049_2 (.CI(GND_net), .I0(n50_adj_4477), .I1(n119_adj_4476), 
            .CO(n39335));
    SB_LUT4 add_6064_8_lut (.I0(GND_net), .I1(n18861[5]), .I2(n560), .I3(n39334), 
            .O(n18749[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6064_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_13_lut (.I0(\PID_CONTROLLER.integral [11]), 
            .I1(GND_net), .I2(n1_adj_4768[11]), .I3(n39243), .O(n23_adj_4417)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_13_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5322_5_lut (.I0(GND_net), .I1(n13364[2]), .I2(n299), .I3(n39977), 
            .O(n12113[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5903_8_lut (.I0(GND_net), .I1(n17069[5]), .I2(n536_adj_4468), 
            .I3(n39861), .O(n16620[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5903_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5903_8 (.CI(n39861), .I0(n17069[5]), .I1(n536_adj_4468), 
            .CO(n39862));
    SB_LUT4 mult_10_i322_2_lut (.I0(\Kp[6] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n478_adj_4543));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i15_1_lut (.I0(IntegralLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[14]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5322_5 (.CI(n39977), .I0(n13364[2]), .I1(n299), .CO(n39978));
    SB_CARRY add_5917_9 (.CI(n39432), .I0(n17265[6]), .I1(n612_adj_4474), 
            .CO(n39433));
    SB_LUT4 add_6064_7_lut (.I0(GND_net), .I1(n18861[4]), .I2(n487), .I3(n39333), 
            .O(n18749[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6064_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i508_2_lut (.I0(\Kp[10] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n755_adj_4540));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i508_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_13 (.CI(n39243), .I0(GND_net), .I1(n1_adj_4768[11]), 
            .CO(n39244));
    SB_LUT4 unary_minus_5_add_3_12_lut (.I0(\PID_CONTROLLER.integral [10]), 
            .I1(GND_net), .I2(n1_adj_4768[10]), .I3(n39242), .O(n21_adj_4407)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_12_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_i749_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1114_adj_4547));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i749_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i557_2_lut (.I0(\Kp[11] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n828_adj_4539));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i73_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n107));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i26_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n38));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5917_8_lut (.I0(GND_net), .I1(n17265[5]), .I2(n539_adj_4465), 
            .I3(n39431), .O(n16845[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5917_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i228_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n338_adj_4538));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i73_2_lut (.I0(\Kp[1] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n107_adj_4549));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i73_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i26_2_lut (.I0(\Kp[0] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n38_adj_4551));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i26_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i698_2_lut (.I0(\Kp[14] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1038));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i698_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6064_7 (.CI(n39333), .I0(n18861[4]), .I1(n487), .CO(n39334));
    SB_LUT4 unary_minus_5_inv_0_i16_1_lut (.I0(IntegralLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[15]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mux_17_i2_3_lut (.I0(duty_23__N_3672[1]), .I1(n257[1]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_5_add_3_12 (.CI(n39242), .I0(GND_net), .I1(n1_adj_4768[10]), 
            .CO(n39243));
    SB_LUT4 duty_23__I_0_i2_3_lut (.I0(duty_23__N_3647[1]), .I1(PWMLimit[1]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[1]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i559_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n831_adj_4536));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i559_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_11_lut (.I0(\PID_CONTROLLER.integral [9]), 
            .I1(GND_net), .I2(n1_adj_4768[9]), .I3(n39241), .O(n19_adj_4408)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_11_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_6064_6_lut (.I0(GND_net), .I1(n18861[3]), .I2(n414), .I3(n39332), 
            .O(n18749[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6064_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i3_3_lut (.I0(duty_23__N_3672[2]), .I1(n257[2]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_6023_4 (.CI(n39541), .I0(n18524[1]), .I1(n259_adj_4475), 
            .CO(n39542));
    SB_LUT4 duty_23__I_0_i3_3_lut (.I0(duty_23__N_3647[2]), .I1(PWMLimit[2]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[2]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i4_3_lut (.I0(duty_23__N_3672[3]), .I1(n257[3]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY unary_minus_5_add_3_11 (.CI(n39241), .I0(GND_net), .I1(n1_adj_4768[9]), 
            .CO(n39242));
    SB_CARRY add_6064_6 (.CI(n39332), .I0(n18861[3]), .I1(n414), .CO(n39333));
    SB_LUT4 duty_23__I_0_i4_3_lut (.I0(duty_23__N_3647[3]), .I1(PWMLimit[3]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[3]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_add_3_10_lut (.I0(\PID_CONTROLLER.integral [8]), 
            .I1(GND_net), .I2(n1_adj_4768[8]), .I3(n39240), .O(n17_adj_4409)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_10_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mux_17_i5_3_lut (.I0(duty_23__N_3672[4]), .I1(n257[4]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i5_3_lut (.I0(duty_23__N_3647[4]), .I1(PWMLimit[4]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[4]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i6_3_lut (.I0(duty_23__N_3672[5]), .I1(n257[5]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i6_3_lut (.I0(duty_23__N_3647[5]), .I1(PWMLimit[5]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[5]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i7_3_lut (.I0(duty_23__N_3672[6]), .I1(n257[6]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i7_3_lut (.I0(duty_23__N_3647[6]), .I1(PWMLimit[6]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[6]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i8_3_lut (.I0(duty_23__N_3672[7]), .I1(n257[7]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i8_3_lut (.I0(duty_23__N_3647[7]), .I1(PWMLimit[7]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[7]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i9_3_lut (.I0(duty_23__N_3672[8]), .I1(n257[8]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i9_3_lut (.I0(duty_23__N_3647[8]), .I1(PWMLimit[8]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[8]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i10_3_lut (.I0(duty_23__N_3672[9]), .I1(n257[9]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i10_3_lut (.I0(duty_23__N_3647[9]), .I1(PWMLimit[9]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[9]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5917_8 (.CI(n39431), .I0(n17265[5]), .I1(n539_adj_4465), 
            .CO(n39432));
    SB_LUT4 mux_17_i11_3_lut (.I0(duty_23__N_3672[10]), .I1(n257[10]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i11_3_lut (.I0(duty_23__N_3647[10]), .I1(PWMLimit[10]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[10]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5903_7_lut (.I0(GND_net), .I1(n17069[4]), .I2(n463), .I3(n39860), 
            .O(n16620[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5903_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i12_3_lut (.I0(duty_23__N_3672[11]), .I1(n257[11]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_5917_7_lut (.I0(GND_net), .I1(n17265[4]), .I2(n466_adj_4460), 
            .I3(n39430), .O(n16845[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5917_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5322_4_lut (.I0(GND_net), .I1(n13364[1]), .I2(n226_adj_4459), 
            .I3(n39976), .O(n12113[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6064_5_lut (.I0(GND_net), .I1(n18861[2]), .I2(n341), .I3(n39331), 
            .O(n18749[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6064_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5917_7 (.CI(n39430), .I0(n17265[4]), .I1(n466_adj_4460), 
            .CO(n39431));
    SB_CARRY add_6064_5 (.CI(n39331), .I0(n18861[2]), .I1(n341), .CO(n39332));
    SB_LUT4 add_5917_6_lut (.I0(GND_net), .I1(n17265[3]), .I2(n393_adj_4457), 
            .I3(n39429), .O(n16845[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5917_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_10 (.CI(n39240), .I0(GND_net), .I1(n1_adj_4768[8]), 
            .CO(n39241));
    SB_CARRY add_5322_4 (.CI(n39976), .I0(n13364[1]), .I1(n226_adj_4459), 
            .CO(n39977));
    SB_LUT4 add_5322_3_lut (.I0(GND_net), .I1(n13364[0]), .I2(n153_adj_4456), 
            .I3(n39975), .O(n12113[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6064_4_lut (.I0(GND_net), .I1(n18861[1]), .I2(n268_adj_4455), 
            .I3(n39330), .O(n18749[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6064_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_0_i12_3_lut (.I0(duty_23__N_3647[11]), .I1(PWMLimit[11]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[11]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 unary_minus_5_add_3_9_lut (.I0(\PID_CONTROLLER.integral [7]), 
            .I1(GND_net), .I2(n1_adj_4768[7]), .I3(n39239), .O(n15_adj_4404)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_9_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mux_17_i13_3_lut (.I0(duty_23__N_3672[12]), .I1(n257[12]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i13_3_lut (.I0(duty_23__N_3647[12]), .I1(PWMLimit[12]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[12]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i14_3_lut (.I0(duty_23__N_3672[13]), .I1(n257[13]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i14_3_lut (.I0(duty_23__N_3647[13]), .I1(PWMLimit[13]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[13]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i15_3_lut (.I0(duty_23__N_3672[14]), .I1(n257[14]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i15_3_lut (.I0(duty_23__N_3647[14]), .I1(PWMLimit[14]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[14]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i16_3_lut (.I0(duty_23__N_3672[15]), .I1(n257[15]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i16_3_lut (.I0(duty_23__N_3647[15]), .I1(PWMLimit[15]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[15]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i17_3_lut (.I0(duty_23__N_3672[16]), .I1(n257[16]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5903_7 (.CI(n39860), .I0(n17069[4]), .I1(n463), .CO(n39861));
    SB_LUT4 duty_23__I_0_i17_3_lut (.I0(duty_23__N_3647[16]), .I1(PWMLimit[16]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[16]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_5322_3 (.CI(n39975), .I0(n13364[0]), .I1(n153_adj_4456), 
            .CO(n39976));
    SB_LUT4 add_5903_6_lut (.I0(GND_net), .I1(n17069[3]), .I2(n390), .I3(n39859), 
            .O(n16620[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5903_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_17_i18_3_lut (.I0(duty_23__N_3672[17]), .I1(n257[17]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i18_3_lut (.I0(duty_23__N_3647[17]), .I1(PWMLimit[17]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[17]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i19_3_lut (.I0(duty_23__N_3672[18]), .I1(n257[18]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i19_3_lut (.I0(duty_23__N_3647[18]), .I1(PWMLimit[18]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[18]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i20_3_lut (.I0(duty_23__N_3672[19]), .I1(n257[19]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i20_3_lut (.I0(duty_23__N_3647[19]), .I1(PWMLimit[19]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[19]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i21_3_lut (.I0(duty_23__N_3672[20]), .I1(n257[20]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i21_3_lut (.I0(duty_23__N_3647[20]), .I1(PWMLimit[20]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[20]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i22_3_lut (.I0(duty_23__N_3672[21]), .I1(n257[21]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i22_3_lut (.I0(duty_23__N_3647[21]), .I1(PWMLimit[21]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[21]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i23_3_lut (.I0(duty_23__N_3672[22]), .I1(n257[22]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i23_3_lut (.I0(duty_23__N_3647[22]), .I1(PWMLimit[22]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[22]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_17_i24_3_lut (.I0(duty_23__N_3672[23]), .I1(n257[23]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i24_3_lut (.I0(duty_23__N_3647[23]), .I1(PWMLimit[23]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[23]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_11_i608_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n904_adj_4535));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i608_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6064_4 (.CI(n39330), .I0(n18861[1]), .I1(n268_adj_4455), 
            .CO(n39331));
    SB_LUT4 unary_minus_5_inv_0_i17_1_lut (.I0(IntegralLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[16]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_5_add_3_9 (.CI(n39239), .I0(GND_net), .I1(n1_adj_4768[7]), 
            .CO(n39240));
    SB_LUT4 mult_11_i277_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n411_adj_4532));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i371_2_lut (.I0(\Kp[7] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n551_adj_4531));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i371_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i657_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n977_adj_4530));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i657_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5903_6 (.CI(n39859), .I0(n17069[3]), .I1(n390), .CO(n39860));
    SB_LUT4 mult_10_i747_2_lut (.I0(\Kp[15] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n1111));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i326_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n484_adj_4529));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i79_2_lut (.I0(\Kp[1] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n116_adj_4556));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i32_2_lut (.I0(\Kp[0] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n47_adj_4557));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6023_3_lut (.I0(GND_net), .I1(n18524[0]), .I2(n186_adj_4453), 
            .I3(n39540), .O(n18325[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6023_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i128_2_lut (.I0(\Kp[2] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n189_adj_4558));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i122_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n180));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i122_2_lut (.I0(\Kp[2] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n180_adj_4559));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i122_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i706_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n1050_adj_4527));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i177_2_lut (.I0(\Kp[3] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n262_adj_4560));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_710_25_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [23]), 
            .I2(n3616[23]), .I3(n39158), .O(\PID_CONTROLLER.integral_23__N_3572 [23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i153_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n226));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i153_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i420_2_lut (.I0(\Kp[8] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n624_adj_4523));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i171_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n253));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6064_3_lut (.I0(GND_net), .I1(n18861[0]), .I2(n195), .I3(n39329), 
            .O(n18749[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6064_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i171_2_lut (.I0(\Kp[3] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n253_adj_4561));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i171_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i59_2_lut (.I0(\Kp[1] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n86));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i12_2_lut (.I0(\Kp[0] ), .I1(n1[5]), .I2(GND_net), 
            .I3(GND_net), .O(n17_adj_4563));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i18_1_lut (.I0(IntegralLimit[17]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[17]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i18_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5322_2_lut (.I0(GND_net), .I1(n11_adj_4399), .I2(n80_adj_4396), 
            .I3(GND_net), .O(n12113[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5322_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5322_2 (.CI(GND_net), .I0(n11_adj_4399), .I1(n80_adj_4396), 
            .CO(n39975));
    SB_LUT4 unary_minus_5_add_3_8_lut (.I0(\PID_CONTROLLER.integral [6]), 
            .I1(GND_net), .I2(n1_adj_4768[6]), .I3(n39238), .O(n13_adj_4405)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_8_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_5903_5_lut (.I0(GND_net), .I1(n17069[2]), .I2(n317), .I3(n39858), 
            .O(n16620[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5903_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5903_5 (.CI(n39858), .I0(n17069[2]), .I1(n317), .CO(n39859));
    SB_LUT4 mult_10_i220_2_lut (.I0(\Kp[4] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n326));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_710_24_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [22]), 
            .I2(n3616[22]), .I3(n39157), .O(\PID_CONTROLLER.integral_23__N_3572 [22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_8 (.CI(n39238), .I0(GND_net), .I1(n1_adj_4768[6]), 
            .CO(n39239));
    SB_LUT4 mult_10_i606_2_lut (.I0(\Kp[12] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n901_adj_4521));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i606_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_710_24 (.CI(n39157), .I0(\PID_CONTROLLER.integral [22]), 
            .I1(n3616[22]), .CO(n39158));
    SB_LUT4 mult_10_i269_2_lut (.I0(\Kp[5] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n399));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5732_21_lut (.I0(GND_net), .I1(n14164[18]), .I2(GND_net), 
            .I3(n39974), .O(n13364[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5903_4_lut (.I0(GND_net), .I1(n17069[1]), .I2(n244), .I3(n39857), 
            .O(n16620[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5903_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i398_2_lut (.I0(\Kp[8] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n591_adj_4520));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i398_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i108_2_lut (.I0(\Kp[2] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n159));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i108_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6064_3 (.CI(n39329), .I0(n18861[0]), .I1(n195), .CO(n39330));
    SB_LUT4 mult_10_i157_2_lut (.I0(\Kp[3] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n232));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i226_2_lut (.I0(\Kp[4] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n335_adj_4564));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i226_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i375_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n557_adj_4519));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i424_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n630_adj_4518));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i206_2_lut (.I0(\Kp[4] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n305));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i206_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6023_3 (.CI(n39540), .I0(n18524[0]), .I1(n186_adj_4453), 
            .CO(n39541));
    SB_LUT4 unary_minus_5_add_3_7_lut (.I0(\PID_CONTROLLER.integral [5]), 
            .I1(GND_net), .I2(n1_adj_4768[5]), .I3(n39237), .O(n11_adj_4406)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_7_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_710_23_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [21]), 
            .I2(n3616[21]), .I3(n39156), .O(\PID_CONTROLLER.integral_23__N_3572 [21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6023_2_lut (.I0(GND_net), .I1(n44), .I2(n113), .I3(GND_net), 
            .O(n18325[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6023_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6023_2 (.CI(GND_net), .I0(n44), .I1(n113), .CO(n39540));
    SB_LUT4 mult_10_i255_2_lut (.I0(\Kp[5] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n378));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i318_2_lut (.I0(\Kp[6] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n472));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i318_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5903_4 (.CI(n39857), .I0(n17069[1]), .I1(n244), .CO(n39858));
    SB_LUT4 add_5903_3_lut (.I0(GND_net), .I1(n17069[0]), .I2(n171), .I3(n39856), 
            .O(n16620[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5903_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5732_20_lut (.I0(GND_net), .I1(n14164[17]), .I2(GND_net), 
            .I3(n39973), .O(n13364[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5732_20 (.CI(n39973), .I0(n14164[17]), .I1(GND_net), 
            .CO(n39974));
    SB_LUT4 mult_10_i304_2_lut (.I0(\Kp[6] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n451));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i304_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5917_6 (.CI(n39429), .I0(n17265[3]), .I1(n393_adj_4457), 
            .CO(n39430));
    SB_LUT4 mult_11_i220_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n326_adj_4565));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i220_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i275_2_lut (.I0(\Kp[5] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n408_adj_4566));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5917_5_lut (.I0(GND_net), .I1(n17265[2]), .I2(n320_adj_4387), 
            .I3(n39428), .O(n16845[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5917_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i51_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n74));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i4_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5_adj_4567));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6064_2_lut (.I0(GND_net), .I1(n53), .I2(n122), .I3(GND_net), 
            .O(n18749[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6064_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i353_2_lut (.I0(\Kp[7] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n524));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i100_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n147));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i324_2_lut (.I0(\Kp[6] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n481_adj_4568));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i367_2_lut (.I0(\Kp[7] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n545));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i367_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6064_2 (.CI(GND_net), .I0(n53), .I1(n122), .CO(n39329));
    SB_LUT4 mult_10_i402_2_lut (.I0(\Kp[8] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n597));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6077_7_lut (.I0(GND_net), .I1(n46537), .I2(n490), .I3(n39328), 
            .O(n18861[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6077_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i67_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n98_adj_4517));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i67_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5903_3 (.CI(n39856), .I0(n17069[0]), .I1(n171), .CO(n39857));
    SB_LUT4 mult_11_i20_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [9]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4516));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i20_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i149_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n220_adj_4569));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i149_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i451_2_lut (.I0(\Kp[9] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n670));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5732_19_lut (.I0(GND_net), .I1(n14164[16]), .I2(GND_net), 
            .I3(n39972), .O(n13364[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i655_2_lut (.I0(\Kp[13] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n974_adj_4515));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5903_2_lut (.I0(GND_net), .I1(n29), .I2(n98), .I3(GND_net), 
            .O(n16620[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5903_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i416_2_lut (.I0(\Kp[8] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n618));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i79_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n116));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i79_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i32_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [15]), 
            .I2(GND_net), .I3(GND_net), .O(n47));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i32_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i469_2_lut (.I0(\Kp[9] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n697_adj_4512));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i518_2_lut (.I0(\Kp[10] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n770_adj_4511));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6077_6_lut (.I0(GND_net), .I1(n18945[3]), .I2(n417), .I3(n39327), 
            .O(n18861[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6077_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_inv_0_i19_1_lut (.I0(IntegralLimit[18]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[18]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i19_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5903_2 (.CI(GND_net), .I0(n29), .I1(n98), .CO(n39856));
    SB_LUT4 unary_minus_5_inv_0_i20_1_lut (.I0(IntegralLimit[19]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[19]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i20_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY unary_minus_5_add_3_7 (.CI(n39237), .I0(GND_net), .I1(n1_adj_4768[5]), 
            .CO(n39238));
    SB_LUT4 add_5931_15_lut (.I0(GND_net), .I1(n17460[12]), .I2(n1050), 
            .I3(n39855), .O(n17069[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5931_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i128_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n189));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i128_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i500_2_lut (.I0(\Kp[10] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n743_adj_4570));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i500_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i116_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n171_adj_4506));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i116_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i465_2_lut (.I0(\Kp[9] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n691));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i465_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i373_2_lut (.I0(\Kp[7] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n554_adj_4571));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i549_2_lut (.I0(\Kp[11] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n816_adj_4572));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i549_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i598_2_lut (.I0(\Kp[12] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n889_adj_4573));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i598_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i514_2_lut (.I0(\Kp[10] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n764));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i269_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n399_adj_4574));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i269_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i563_2_lut (.I0(\Kp[11] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n837));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i612_2_lut (.I0(\Kp[12] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n910));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i647_2_lut (.I0(\Kp[13] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n962_adj_4575));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i647_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i198_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n293_adj_4576));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i198_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i318_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n472_adj_4577));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i318_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_710_23 (.CI(n39156), .I0(\PID_CONTROLLER.integral [21]), 
            .I1(n3616[21]), .CO(n39157));
    SB_CARRY add_5732_19 (.CI(n39972), .I0(n14164[16]), .I1(GND_net), 
            .CO(n39973));
    SB_CARRY add_6077_6 (.CI(n39327), .I0(n18945[3]), .I1(n417), .CO(n39328));
    SB_CARRY add_5917_5 (.CI(n39428), .I0(n17265[2]), .I1(n320_adj_4387), 
            .CO(n39429));
    SB_LUT4 add_5917_4_lut (.I0(GND_net), .I1(n17265[1]), .I2(n247_adj_4370), 
            .I3(n39427), .O(n16845[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5917_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5732_18_lut (.I0(GND_net), .I1(n14164[15]), .I2(GND_net), 
            .I3(n39971), .O(n13364[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6077_5_lut (.I0(GND_net), .I1(n18945[2]), .I2(n344), .I3(n39326), 
            .O(n18861[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6077_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5931_14_lut (.I0(GND_net), .I1(n17460[11]), .I2(n977), 
            .I3(n39854), .O(n17069[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5931_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_6_lut (.I0(\PID_CONTROLLER.integral [4]), 
            .I1(GND_net), .I2(n1_adj_4768[4]), .I3(n39236), .O(n9_adj_4410)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_6_lut.LUT_INIT = 16'h6996;
    SB_CARRY add_6077_5 (.CI(n39326), .I0(n18945[2]), .I1(n344), .CO(n39327));
    SB_CARRY add_5931_14 (.CI(n39854), .I0(n17460[11]), .I1(n977), .CO(n39855));
    SB_CARRY add_5732_18 (.CI(n39971), .I0(n14164[15]), .I1(GND_net), 
            .CO(n39972));
    SB_CARRY add_5917_4 (.CI(n39427), .I0(n17265[1]), .I1(n247_adj_4370), 
            .CO(n39428));
    SB_LUT4 add_5931_13_lut (.I0(GND_net), .I1(n17460[10]), .I2(n904), 
            .I3(n39853), .O(n17069[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5931_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i57_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n83));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i10_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n14_adj_4504));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i177_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n262));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i177_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i447_2_lut (.I0(\Kp[9] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n664_adj_4503));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i447_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i165_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n244_adj_4502));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i165_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i21_1_lut (.I0(IntegralLimit[20]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[20]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i21_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i704_2_lut (.I0(\Kp[14] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1047_adj_4500));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i704_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5931_13 (.CI(n39853), .I0(n17460[10]), .I1(n904), .CO(n39854));
    SB_LUT4 add_5732_17_lut (.I0(GND_net), .I1(n14164[14]), .I2(GND_net), 
            .I3(n39970), .O(n13364[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i226_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n335));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i226_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_6 (.CI(n39236), .I0(GND_net), .I1(n1_adj_4768[4]), 
            .CO(n39237));
    SB_LUT4 mult_11_i247_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n366_adj_4578));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i247_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_add_3_5_lut (.I0(\PID_CONTROLLER.integral [3]), 
            .I1(GND_net), .I2(n1_adj_4768[3]), .I3(n39235), .O(n7_adj_4414)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_5_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_i422_2_lut (.I0(\Kp[8] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n627_adj_4579));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i367_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n545_adj_4580));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i367_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6077_4_lut (.I0(GND_net), .I1(n18945[1]), .I2(n271_adj_4369), 
            .I3(n39325), .O(n18861[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6077_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i696_2_lut (.I0(\Kp[14] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1035_adj_4581));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i296_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n439_adj_4582));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i296_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i471_2_lut (.I0(\Kp[9] ), .I1(n1[14]), .I2(GND_net), 
            .I3(GND_net), .O(n700_adj_4583));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i345_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n512_adj_4584));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i345_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i61_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n89_adj_4585));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i61_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i753_2_lut (.I0(\Kp[15] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n1120_adj_4499));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i753_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i496_2_lut (.I0(\Kp[10] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n737_adj_4498));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i496_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i106_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n156));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i106_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i14_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [6]), 
            .I2(GND_net), .I3(GND_net), .O(n20_adj_4586));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i14_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i65_2_lut (.I0(\Kp[1] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n95_adj_4497));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i18_2_lut (.I0(\Kp[0] ), .I1(n1[8]), .I2(GND_net), 
            .I3(GND_net), .O(n26_adj_4496));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i18_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY unary_minus_5_add_3_5 (.CI(n39235), .I0(GND_net), .I1(n1_adj_4768[3]), 
            .CO(n39236));
    SB_CARRY add_6077_4 (.CI(n39325), .I0(n18945[1]), .I1(n271_adj_4369), 
            .CO(n39326));
    SB_LUT4 mult_11_i214_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n317_adj_4494));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i214_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6077_3_lut (.I0(GND_net), .I1(n18945[0]), .I2(n198), .I3(n39324), 
            .O(n18861[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6077_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i545_2_lut (.I0(\Kp[11] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n810_adj_4489));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i545_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i594_2_lut (.I0(\Kp[12] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n883_adj_4488));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i594_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i263_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n390_adj_4487));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i263_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5931_12_lut (.I0(GND_net), .I1(n17460[9]), .I2(n831), 
            .I3(n39852), .O(n17069[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5931_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5732_17 (.CI(n39970), .I0(n14164[14]), .I1(GND_net), 
            .CO(n39971));
    SB_LUT4 add_5732_16_lut (.I0(GND_net), .I1(n14164[13]), .I2(n1105), 
            .I3(n39969), .O(n13364[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5931_12 (.CI(n39852), .I0(n17460[9]), .I1(n831), .CO(n39853));
    SB_LUT4 add_5931_11_lut (.I0(GND_net), .I1(n17460[8]), .I2(n758), 
            .I3(n39851), .O(n17069[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5931_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5732_16 (.CI(n39969), .I0(n14164[13]), .I1(n1105), .CO(n39970));
    SB_LUT4 add_5732_15_lut (.I0(GND_net), .I1(n14164[12]), .I2(n1032), 
            .I3(n39968), .O(n13364[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5732_15 (.CI(n39968), .I0(n14164[12]), .I1(n1032), .CO(n39969));
    SB_CARRY add_5931_11 (.CI(n39851), .I0(n17460[8]), .I1(n758), .CO(n39852));
    SB_LUT4 add_710_22_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [20]), 
            .I2(n3616[20]), .I3(n39155), .O(\PID_CONTROLLER.integral_23__N_3572 [20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5931_10_lut (.I0(GND_net), .I1(n17460[7]), .I2(n685), 
            .I3(n39850), .O(n17069[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5931_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5732_14_lut (.I0(GND_net), .I1(n14164[11]), .I2(n959), 
            .I3(n39967), .O(n13364[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5732_14 (.CI(n39967), .I0(n14164[11]), .I1(n959), .CO(n39968));
    SB_CARRY add_5931_10 (.CI(n39850), .I0(n17460[7]), .I1(n685), .CO(n39851));
    SB_LUT4 mult_10_i71_2_lut (.I0(\Kp[1] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n104));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5732_13_lut (.I0(GND_net), .I1(n14164[10]), .I2(n886), 
            .I3(n39966), .O(n13364[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i24_2_lut (.I0(\Kp[0] ), .I1(n1[11]), .I2(GND_net), 
            .I3(GND_net), .O(n35_adj_4587));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i416_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n618_adj_4588));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i416_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i745_2_lut (.I0(\Kp[15] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n1108_adj_4589));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i745_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5931_9_lut (.I0(GND_net), .I1(n17460[6]), .I2(n612), .I3(n39849), 
            .O(n17069[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5931_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5732_13 (.CI(n39966), .I0(n14164[10]), .I1(n886), .CO(n39967));
    SB_CARRY add_5931_9 (.CI(n39849), .I0(n17460[6]), .I1(n612), .CO(n39850));
    SB_LUT4 add_5917_3_lut (.I0(GND_net), .I1(n17265[0]), .I2(n174_adj_4367), 
            .I3(n39426), .O(n16845[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5917_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i120_2_lut (.I0(\Kp[2] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n177));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i465_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n691_adj_4590));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i465_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6077_3 (.CI(n39324), .I0(n18945[0]), .I1(n198), .CO(n39325));
    SB_LUT4 mult_11_i110_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n162_adj_4591));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i110_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i514_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n764_adj_4592));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i514_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5732_12_lut (.I0(GND_net), .I1(n14164[9]), .I2(n813), 
            .I3(n39965), .O(n13364[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i394_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n585_adj_4593));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i394_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i22_1_lut (.I0(IntegralLimit[21]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[21]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i22_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5732_12 (.CI(n39965), .I0(n14164[9]), .I1(n813), .CO(n39966));
    SB_LUT4 add_5931_8_lut (.I0(GND_net), .I1(n17460[5]), .I2(n539), .I3(n39848), 
            .O(n17069[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5931_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5917_3 (.CI(n39426), .I0(n17265[0]), .I1(n174_adj_4367), 
            .CO(n39427));
    SB_CARRY add_5931_8 (.CI(n39848), .I0(n17460[5]), .I1(n539), .CO(n39849));
    SB_LUT4 unary_minus_5_add_3_4_lut (.I0(\PID_CONTROLLER.integral [2]), 
            .I1(GND_net), .I2(n1_adj_4768[2]), .I3(n39234), .O(n5_adj_4415)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_4_lut.LUT_INIT = 16'h6996;
    SB_CARRY unary_minus_5_add_3_4 (.CI(n39234), .I0(GND_net), .I1(n1_adj_4768[2]), 
            .CO(n39235));
    SB_LUT4 add_5917_2_lut (.I0(GND_net), .I1(n32_adj_4365), .I2(n101_adj_4364), 
            .I3(GND_net), .O(n16845[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5917_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_710_22 (.CI(n39155), .I0(\PID_CONTROLLER.integral [20]), 
            .I1(n3616[20]), .CO(n39156));
    SB_LUT4 add_5931_7_lut (.I0(GND_net), .I1(n17460[4]), .I2(n466), .I3(n39847), 
            .O(n17069[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5931_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6077_2_lut (.I0(GND_net), .I1(n56), .I2(n125), .I3(GND_net), 
            .O(n18861[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6077_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_3_lut (.I0(\PID_CONTROLLER.integral [1]), 
            .I1(GND_net), .I2(n1_adj_4768[1]), .I3(n39233), .O(n3_adj_4433)) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_3_lut.LUT_INIT = 16'h6996;
    SB_LUT4 add_710_21_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [19]), 
            .I2(n3616[19]), .I3(n39154), .O(\PID_CONTROLLER.integral_23__N_3572 [19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_710_21 (.CI(n39154), .I0(\PID_CONTROLLER.integral [19]), 
            .I1(n3616[19]), .CO(n39155));
    SB_CARRY add_5931_7 (.CI(n39847), .I0(n17460[4]), .I1(n466), .CO(n39848));
    SB_LUT4 add_5732_11_lut (.I0(GND_net), .I1(n14164[8]), .I2(n740), 
            .I3(n39964), .O(n13364[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5931_6_lut (.I0(GND_net), .I1(n17460[3]), .I2(n393), .I3(n39846), 
            .O(n17069[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5931_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5931_6 (.CI(n39846), .I0(n17460[3]), .I1(n393), .CO(n39847));
    SB_LUT4 add_710_20_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [18]), 
            .I2(n3616[18]), .I3(n39153), .O(\PID_CONTROLLER.integral_23__N_3572 [18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5917_2 (.CI(GND_net), .I0(n32_adj_4365), .I1(n101_adj_4364), 
            .CO(n39426));
    SB_CARRY add_6077_2 (.CI(GND_net), .I0(n56), .I1(n125), .CO(n39324));
    SB_CARRY unary_minus_5_add_3_3 (.CI(n39233), .I0(GND_net), .I1(n1_adj_4768[1]), 
            .CO(n39234));
    SB_LUT4 add_5752_20_lut (.I0(GND_net), .I1(n14525[17]), .I2(GND_net), 
            .I3(n39533), .O(n13765[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_5_add_3_2_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4768[0]), 
            .I3(VCC_net), .O(\PID_CONTROLLER.integral_23__N_3623 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_5_add_3_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_5_add_3_2 (.CI(VCC_net), .I0(GND_net), .I1(n1_adj_4768[0]), 
            .CO(n39233));
    SB_CARRY add_5732_11 (.CI(n39964), .I0(n14164[8]), .I1(n740), .CO(n39965));
    SB_LUT4 add_5931_5_lut (.I0(GND_net), .I1(n17460[2]), .I2(n320), .I3(n39845), 
            .O(n17069[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5931_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_710_20 (.CI(n39153), .I0(\PID_CONTROLLER.integral [18]), 
            .I1(n3616[18]), .CO(n39154));
    SB_CARRY add_5931_5 (.CI(n39845), .I0(n17460[2]), .I1(n320), .CO(n39846));
    SB_LUT4 add_5732_10_lut (.I0(GND_net), .I1(n14164[7]), .I2(n667), 
            .I3(n39963), .O(n13364[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5931_4_lut (.I0(GND_net), .I1(n17460[1]), .I2(n247), .I3(n39844), 
            .O(n17069[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5931_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5931_4 (.CI(n39844), .I0(n17460[1]), .I1(n247), .CO(n39845));
    SB_LUT4 add_5931_3_lut (.I0(GND_net), .I1(n17460[0]), .I2(n174), .I3(n39843), 
            .O(n17069[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5931_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5752_19_lut (.I0(GND_net), .I1(n14525[16]), .I2(GND_net), 
            .I3(n39532), .O(n13765[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i155_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n229));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i275_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n408));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i275_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i114_2_lut (.I0(\Kp[2] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n168_adj_4485));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i114_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5752_19 (.CI(n39532), .I0(n14525[16]), .I1(GND_net), 
            .CO(n39533));
    SB_LUT4 add_5752_18_lut (.I0(GND_net), .I1(n14525[15]), .I2(GND_net), 
            .I3(n39531), .O(n13765[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5752_18 (.CI(n39531), .I0(n14525[15]), .I1(GND_net), 
            .CO(n39532));
    SB_LUT4 sub_3_add_2_25_lut (.I0(GND_net), .I1(setpoint[23]), .I2(motor_state[23]), 
            .I3(n39232), .O(n1[23])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_710_19_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [17]), 
            .I2(n3616[17]), .I3(n39152), .O(\PID_CONTROLLER.integral_23__N_3572 [17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5752_17_lut (.I0(GND_net), .I1(n14525[14]), .I2(GND_net), 
            .I3(n39530), .O(n13765[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_24_lut (.I0(GND_net), .I1(setpoint[22]), .I2(motor_state[22]), 
            .I3(n39231), .O(n1[22])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i643_2_lut (.I0(\Kp[13] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n956_adj_4483));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i643_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_5_inv_0_i23_1_lut (.I0(IntegralLimit[22]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[22]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i204_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n302));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i204_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5752_17 (.CI(n39530), .I0(n14525[14]), .I1(GND_net), 
            .CO(n39531));
    SB_LUT4 add_5752_16_lut (.I0(GND_net), .I1(n14525[13]), .I2(n1108), 
            .I3(n39529), .O(n13765[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5732_10 (.CI(n39963), .I0(n14164[7]), .I1(n667), .CO(n39964));
    SB_CARRY add_5752_16 (.CI(n39529), .I0(n14525[13]), .I1(n1108), .CO(n39530));
    SB_LUT4 unary_minus_5_inv_0_i24_1_lut (.I0(IntegralLimit[23]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4768[23]));   // verilog/motorControl.v(31[48:62])
    defparam unary_minus_5_inv_0_i24_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_5752_15_lut (.I0(GND_net), .I1(n14525[12]), .I2(n1035), 
            .I3(n39528), .O(n13765[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5732_9_lut (.I0(GND_net), .I1(n14164[6]), .I2(n594), .I3(n39962), 
            .O(n13364[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_24 (.CI(n39231), .I0(setpoint[22]), .I1(motor_state[22]), 
            .CO(n39232));
    SB_CARRY add_5752_15 (.CI(n39528), .I0(n14525[12]), .I1(n1035), .CO(n39529));
    SB_LUT4 add_5752_14_lut (.I0(GND_net), .I1(n14525[11]), .I2(n962), 
            .I3(n39527), .O(n13765[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_23_lut (.I0(GND_net), .I1(setpoint[21]), .I2(motor_state[21]), 
            .I3(n39230), .O(n1[21])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5752_14 (.CI(n39527), .I0(n14525[11]), .I1(n962), .CO(n39528));
    SB_CARRY add_710_19 (.CI(n39152), .I0(\PID_CONTROLLER.integral [17]), 
            .I1(n3616[17]), .CO(n39153));
    SB_CARRY sub_3_add_2_23 (.CI(n39230), .I0(setpoint[21]), .I1(motor_state[21]), 
            .CO(n39231));
    SB_CARRY add_5732_9 (.CI(n39962), .I0(n14164[6]), .I1(n594), .CO(n39963));
    SB_CARRY add_5931_3 (.CI(n39843), .I0(n17460[0]), .I1(n174), .CO(n39844));
    SB_LUT4 mult_10_i163_2_lut (.I0(\Kp[3] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n241_adj_4472));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_22_lut (.I0(GND_net), .I1(setpoint[20]), .I2(motor_state[20]), 
            .I3(n39229), .O(n1[20])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i443_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n658_adj_4594));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i443_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i324_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n481));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i324_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i159_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n235_adj_4595));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i159_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i208_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n308_adj_4596));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i208_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i312_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n463_adj_4470));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i312_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i253_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n375));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i692_2_lut (.I0(\Kp[14] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1029_adj_4469));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i692_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i492_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n731_adj_4597));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i492_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i75_2_lut (.I0(\Kp[1] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n110));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i28_2_lut (.I0(\Kp[0] ), .I1(n1[13]), .I2(GND_net), 
            .I3(GND_net), .O(n41_adj_4598));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i741_2_lut (.I0(\Kp[15] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n1102_adj_4467));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i741_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i302_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n448_adj_4463));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i302_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i1_1_lut (.I0(PWMLimit[0]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[0]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i257_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n381_adj_4599));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i257_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i373_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n554));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i373_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i361_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n536));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i361_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i169_2_lut (.I0(\Kp[3] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n250));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i169_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i541_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n804_adj_4600));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i541_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5752_13_lut (.I0(GND_net), .I1(n14525[10]), .I2(n889), 
            .I3(n39526), .O(n13765[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i410_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n609));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i410_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i124_2_lut (.I0(\Kp[2] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n183));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i422_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n627));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i422_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i563_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n837_adj_4601));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i563_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i306_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n454_adj_4602));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i306_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5931_2_lut (.I0(GND_net), .I1(n32), .I2(n101), .I3(GND_net), 
            .O(n17069[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5931_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i612_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n910_adj_4603));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i612_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_710_18_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [16]), 
            .I2(n3616[16]), .I3(n39151), .O(\PID_CONTROLLER.integral_23__N_3572 [16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5752_13 (.CI(n39526), .I0(n14525[10]), .I1(n889), .CO(n39527));
    SB_LUT4 add_5752_12_lut (.I0(GND_net), .I1(n14525[9]), .I2(n816), 
            .I3(n39525), .O(n13765[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i355_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n527_adj_4604));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i355_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i173_2_lut (.I0(\Kp[3] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n256_adj_4605));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i173_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i590_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n877_adj_4606));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i590_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i71_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n104_adj_4607));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i71_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i24_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [11]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4608));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i24_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i218_2_lut (.I0(\Kp[4] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n323));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i404_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n600_adj_4609));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i404_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i212_2_lut (.I0(\Kp[4] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n314));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i36456_1_lut (.I0(duty[23]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n51409));   // verilog/motorControl.v(29[14] 48[8])
    defparam i36456_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i453_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n673_adj_4610));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i453_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i471_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n700));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i471_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i351_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n521_adj_4458));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i351_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i400_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n594_adj_4452));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i400_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i459_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n682));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i459_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i2_1_lut (.I0(PWMLimit[1]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[1]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i2_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_710_18 (.CI(n39151), .I0(\PID_CONTROLLER.integral [16]), 
            .I1(n3616[16]), .CO(n39152));
    SB_CARRY sub_3_add_2_22 (.CI(n39229), .I0(setpoint[20]), .I1(motor_state[20]), 
            .CO(n39230));
    SB_CARRY add_5752_12 (.CI(n39525), .I0(n14525[9]), .I1(n816), .CO(n39526));
    SB_LUT4 mult_11_i639_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n950_adj_4611));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i639_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i120_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n177_adj_4612));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i120_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i169_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n250_adj_4613));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i169_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5931_2 (.CI(GND_net), .I0(n32), .I1(n101), .CO(n39843));
    SB_LUT4 add_710_17_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [15]), 
            .I2(n3616[15]), .I3(n39150), .O(\PID_CONTROLLER.integral_23__N_3572 [15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i502_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n746_adj_4614));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i502_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i77_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n113_adj_4449));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i77_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i30_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [14]), 
            .I2(GND_net), .I3(GND_net), .O(n44_adj_4448));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i30_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5732_8_lut (.I0(GND_net), .I1(n14164[5]), .I2(n521), .I3(n39961), 
            .O(n13364[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i57_2_lut (.I0(\Kp[1] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n83_adj_4615));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i57_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_21_lut (.I0(GND_net), .I1(setpoint[19]), .I2(motor_state[19]), 
            .I3(n39228), .O(n1[19])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_21 (.CI(n39228), .I0(setpoint[19]), .I1(motor_state[19]), 
            .CO(n39229));
    SB_LUT4 add_5752_11_lut (.I0(GND_net), .I1(n14525[8]), .I2(n743), 
            .I3(n39524), .O(n13765[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i10_2_lut (.I0(\Kp[0] ), .I1(n1[4]), .I2(GND_net), 
            .I3(GND_net), .O(n14_adj_4616));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i10_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i449_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n667_adj_4447));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i449_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_20_lut (.I0(GND_net), .I1(setpoint[18]), .I2(motor_state[18]), 
            .I3(n39227), .O(n1[18])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_710_17 (.CI(n39150), .I0(\PID_CONTROLLER.integral [15]), 
            .I1(n3616[15]), .CO(n39151));
    SB_CARRY add_5732_8 (.CI(n39961), .I0(n14164[5]), .I1(n521), .CO(n39962));
    SB_LUT4 add_5732_7_lut (.I0(GND_net), .I1(n14164[4]), .I2(n448), .I3(n39960), 
            .O(n13364[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i261_2_lut (.I0(\Kp[5] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n387));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i261_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5752_11 (.CI(n39524), .I0(n14525[8]), .I1(n743), .CO(n39525));
    SB_LUT4 add_5957_14_lut (.I0(GND_net), .I1(n17797[11]), .I2(n980), 
            .I3(n39842), .O(n17460[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_710_16_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [14]), 
            .I2(n3616[14]), .I3(n39149), .O(\PID_CONTROLLER.integral_23__N_3572 [14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_20 (.CI(n39227), .I0(setpoint[18]), .I1(motor_state[18]), 
            .CO(n39228));
    SB_CARRY add_5732_7 (.CI(n39960), .I0(n14164[4]), .I1(n448), .CO(n39961));
    SB_LUT4 add_5957_13_lut (.I0(GND_net), .I1(n17797[10]), .I2(n907), 
            .I3(n39841), .O(n17460[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_710_16 (.CI(n39149), .I0(\PID_CONTROLLER.integral [14]), 
            .I1(n3616[14]), .CO(n39150));
    SB_CARRY add_5957_13 (.CI(n39841), .I0(n17797[10]), .I1(n907), .CO(n39842));
    SB_LUT4 mult_11_i218_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n323_adj_4617));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i218_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i267_2_lut (.I0(\Kp[5] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n396));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5752_10_lut (.I0(GND_net), .I1(n14525[7]), .I2(n670_adj_4618), 
            .I3(n39523), .O(n13765[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5732_6_lut (.I0(GND_net), .I1(n14164[3]), .I2(n375_adj_4619), 
            .I3(n39959), .O(n13364[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5752_10 (.CI(n39523), .I0(n14525[7]), .I1(n670_adj_4618), 
            .CO(n39524));
    SB_CARRY add_5732_6 (.CI(n39959), .I0(n14164[3]), .I1(n375_adj_4619), 
            .CO(n39960));
    SB_LUT4 add_5957_12_lut (.I0(GND_net), .I1(n17797[9]), .I2(n834), 
            .I3(n39840), .O(n17460[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5957_12 (.CI(n39840), .I0(n17797[9]), .I1(n834), .CO(n39841));
    SB_LUT4 mult_10_i316_2_lut (.I0(\Kp[6] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n469));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_19_lut (.I0(GND_net), .I1(setpoint[17]), .I2(motor_state[17]), 
            .I3(n39226), .O(n1[17])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5752_9_lut (.I0(GND_net), .I1(n14525[6]), .I2(n597_adj_4620), 
            .I3(n39522), .O(n13765[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_19 (.CI(n39226), .I0(setpoint[17]), .I1(motor_state[17]), 
            .CO(n39227));
    SB_CARRY add_5752_9 (.CI(n39522), .I0(n14525[6]), .I1(n597_adj_4620), 
            .CO(n39523));
    SB_LUT4 add_5752_8_lut (.I0(GND_net), .I1(n14525[5]), .I2(n524_adj_4621), 
            .I3(n39521), .O(n13765[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_18_lut (.I0(GND_net), .I1(setpoint[16]), .I2(motor_state[16]), 
            .I3(n39225), .O(n1[16])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_18 (.CI(n39225), .I0(setpoint[16]), .I1(motor_state[16]), 
            .CO(n39226));
    SB_LUT4 add_5957_11_lut (.I0(GND_net), .I1(n17797[8]), .I2(n761), 
            .I3(n39839), .O(n17460[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5752_8 (.CI(n39521), .I0(n14525[5]), .I1(n524_adj_4621), 
            .CO(n39522));
    SB_LUT4 add_710_15_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [13]), 
            .I2(n3616[13]), .I3(n39148), .O(\PID_CONTROLLER.integral_23__N_3572 [13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20558_2_lut (.I0(n1[0]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[0]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20558_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i267_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n396_adj_4622));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i267_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_24_lut (.I0(\PID_CONTROLLER.integral_23__N_3572 [23]), 
            .I1(n9339[21]), .I2(GND_net), .I3(n39630), .O(n8832[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_11_add_1225_23_lut (.I0(GND_net), .I1(n9339[20]), .I2(GND_net), 
            .I3(n39629), .O(n155[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5752_7_lut (.I0(GND_net), .I1(n14525[4]), .I2(n451_adj_4623), 
            .I3(n39520), .O(n13765[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_23 (.CI(n39629), .I0(n9339[20]), .I1(GND_net), 
            .CO(n39630));
    SB_LUT4 add_5732_5_lut (.I0(GND_net), .I1(n14164[2]), .I2(n302_adj_4624), 
            .I3(n39958), .O(n13364[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5752_7 (.CI(n39520), .I0(n14525[4]), .I1(n451_adj_4623), 
            .CO(n39521));
    SB_LUT4 add_6003_12_lut (.I0(GND_net), .I1(n18325[9]), .I2(n840_adj_4625), 
            .I3(n39734), .O(n18084[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6003_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_22_lut (.I0(GND_net), .I1(n9339[19]), .I2(GND_net), 
            .I3(n39628), .O(n155[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_710_15 (.CI(n39148), .I0(\PID_CONTROLLER.integral [13]), 
            .I1(n3616[13]), .CO(n39149));
    SB_CARRY add_5732_5 (.CI(n39958), .I0(n14164[2]), .I1(n302_adj_4624), 
            .CO(n39959));
    SB_CARRY add_5957_11 (.CI(n39839), .I0(n17797[8]), .I1(n761), .CO(n39840));
    SB_LUT4 add_5752_6_lut (.I0(GND_net), .I1(n14525[3]), .I2(n378_adj_4626), 
            .I3(n39519), .O(n13765[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5752_6 (.CI(n39519), .I0(n14525[3]), .I1(n378_adj_4626), 
            .CO(n39520));
    SB_LUT4 add_6003_11_lut (.I0(GND_net), .I1(n18325[8]), .I2(n767_adj_4627), 
            .I3(n39733), .O(n18084[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6003_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6003_11 (.CI(n39733), .I0(n18325[8]), .I1(n767_adj_4627), 
            .CO(n39734));
    SB_LUT4 add_6071_8_lut (.I0(GND_net), .I1(n18909[5]), .I2(n560_adj_4628), 
            .I3(n39414), .O(n18812[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6071_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6071_7_lut (.I0(GND_net), .I1(n18909[4]), .I2(n487_adj_4629), 
            .I3(n39413), .O(n18812[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6071_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5957_10_lut (.I0(GND_net), .I1(n17797[7]), .I2(n688), 
            .I3(n39838), .O(n17460[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6003_10_lut (.I0(GND_net), .I1(n18325[7]), .I2(n694_adj_4630), 
            .I3(n39732), .O(n18084[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6003_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_17_lut (.I0(GND_net), .I1(setpoint[15]), .I2(motor_state[15]), 
            .I3(n39224), .O(n1[15])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_710_14_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [12]), 
            .I2(n3616[12]), .I3(n39147), .O(\PID_CONTROLLER.integral_23__N_3572 [12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_22 (.CI(n39628), .I0(n9339[19]), .I1(GND_net), 
            .CO(n39629));
    SB_CARRY sub_3_add_2_17 (.CI(n39224), .I0(setpoint[15]), .I1(motor_state[15]), 
            .CO(n39225));
    SB_LUT4 add_5752_5_lut (.I0(GND_net), .I1(n14525[2]), .I2(n305_adj_4631), 
            .I3(n39518), .O(n13765[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6071_7 (.CI(n39413), .I0(n18909[4]), .I1(n487_adj_4629), 
            .CO(n39414));
    SB_LUT4 add_6071_6_lut (.I0(GND_net), .I1(n18909[3]), .I2(n414_adj_4632), 
            .I3(n39412), .O(n18812[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6071_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5752_5 (.CI(n39518), .I0(n14525[2]), .I1(n305_adj_4631), 
            .CO(n39519));
    SB_CARRY add_710_14 (.CI(n39147), .I0(\PID_CONTROLLER.integral [12]), 
            .I1(n3616[12]), .CO(n39148));
    SB_LUT4 add_5752_4_lut (.I0(GND_net), .I1(n14525[1]), .I2(n232_adj_4633), 
            .I3(n39517), .O(n13765[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5752_4 (.CI(n39517), .I0(n14525[1]), .I1(n232_adj_4633), 
            .CO(n39518));
    SB_CARRY add_6071_6 (.CI(n39412), .I0(n18909[3]), .I1(n414_adj_4632), 
            .CO(n39413));
    SB_LUT4 add_5752_3_lut (.I0(GND_net), .I1(n14525[0]), .I2(n159_adj_4634), 
            .I3(n39516), .O(n13765[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_16_lut (.I0(GND_net), .I1(setpoint[14]), .I2(motor_state[14]), 
            .I3(n39223), .O(n1[14])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6071_5_lut (.I0(GND_net), .I1(n18909[2]), .I2(n341_adj_4635), 
            .I3(n39411), .O(n18812[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6071_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_16 (.CI(n39223), .I0(setpoint[14]), .I1(motor_state[14]), 
            .CO(n39224));
    SB_LUT4 sub_3_add_2_15_lut (.I0(GND_net), .I1(setpoint[13]), .I2(motor_state[13]), 
            .I3(n39222), .O(n1[13])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6071_5 (.CI(n39411), .I0(n18909[2]), .I1(n341_adj_4635), 
            .CO(n39412));
    SB_LUT4 add_6071_4_lut (.I0(GND_net), .I1(n18909[1]), .I2(n268_adj_4636), 
            .I3(n39410), .O(n18812[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6071_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_15 (.CI(n39222), .I0(setpoint[13]), .I1(motor_state[13]), 
            .CO(n39223));
    SB_LUT4 add_710_13_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [11]), 
            .I2(n3616[11]), .I3(n39146), .O(\PID_CONTROLLER.integral_23__N_3572 [11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_710_13 (.CI(n39146), .I0(\PID_CONTROLLER.integral [11]), 
            .I1(n3616[11]), .CO(n39147));
    SB_LUT4 mult_11_i163_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n241));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i163_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i316_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n469_adj_4637));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i316_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i551_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n819_adj_4638));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i551_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20708_2_lut (.I0(n1[1]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[1]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20708_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i222_2_lut (.I0(\Kp[4] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n329_adj_4639));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i222_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i365_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n542));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_21_lut (.I0(GND_net), .I1(n9339[18]), .I2(GND_net), 
            .I3(n39627), .O(n155[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i600_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n892_adj_4641));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i600_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i688_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1023_adj_4642));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i688_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i737_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [0]), 
            .I2(GND_net), .I3(GND_net), .O(n1096_adj_4643));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i737_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5752_3 (.CI(n39516), .I0(n14525[0]), .I1(n159_adj_4634), 
            .CO(n39517));
    SB_LUT4 add_710_12_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [10]), 
            .I2(n3616[10]), .I3(n39145), .O(\PID_CONTROLLER.integral_23__N_3572 [10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5752_2_lut (.I0(GND_net), .I1(n17_adj_4644), .I2(n86_adj_4645), 
            .I3(GND_net), .O(n13765[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5752_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_14_lut (.I0(GND_net), .I1(setpoint[12]), .I2(motor_state[12]), 
            .I3(n39221), .O(n1[12])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6071_4 (.CI(n39410), .I0(n18909[1]), .I1(n268_adj_4636), 
            .CO(n39411));
    SB_CARRY add_5957_10 (.CI(n39838), .I0(n17797[7]), .I1(n688), .CO(n39839));
    SB_CARRY add_710_12 (.CI(n39145), .I0(\PID_CONTROLLER.integral [10]), 
            .I1(n3616[10]), .CO(n39146));
    SB_CARRY mult_11_add_1225_21 (.CI(n39627), .I0(n9339[18]), .I1(GND_net), 
            .CO(n39628));
    SB_LUT4 mult_11_add_1225_20_lut (.I0(GND_net), .I1(n9339[17]), .I2(GND_net), 
            .I3(n39626), .O(n155[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5752_2 (.CI(GND_net), .I0(n17_adj_4644), .I1(n86_adj_4645), 
            .CO(n39516));
    SB_LUT4 add_5789_19_lut (.I0(GND_net), .I1(n15209[16]), .I2(GND_net), 
            .I3(n39515), .O(n14525[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5789_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_20 (.CI(n39626), .I0(n9339[17]), .I1(GND_net), 
            .CO(n39627));
    SB_CARRY add_6003_10 (.CI(n39732), .I0(n18325[7]), .I1(n694_adj_4630), 
            .CO(n39733));
    SB_CARRY sub_3_add_2_14 (.CI(n39221), .I0(setpoint[12]), .I1(motor_state[12]), 
            .CO(n39222));
    SB_LUT4 add_710_11_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [9]), 
            .I2(n3616[9]), .I3(n39144), .O(\PID_CONTROLLER.integral_23__N_3572 [9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6071_3_lut (.I0(GND_net), .I1(n18909[0]), .I2(n195_adj_4646), 
            .I3(n39409), .O(n18812[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6071_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6071_3 (.CI(n39409), .I0(n18909[0]), .I1(n195_adj_4646), 
            .CO(n39410));
    SB_LUT4 sub_3_add_2_13_lut (.I0(GND_net), .I1(setpoint[11]), .I2(motor_state[11]), 
            .I3(n39220), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_13 (.CI(n39220), .I0(setpoint[11]), .I1(motor_state[11]), 
            .CO(n39221));
    SB_LUT4 add_5957_9_lut (.I0(GND_net), .I1(n17797[6]), .I2(n615), .I3(n39837), 
            .O(n17460[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i498_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n740_adj_4445));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i498_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5789_18_lut (.I0(GND_net), .I1(n15209[15]), .I2(GND_net), 
            .I3(n39514), .O(n14525[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5789_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_710_11 (.CI(n39144), .I0(\PID_CONTROLLER.integral [9]), 
            .I1(n3616[9]), .CO(n39145));
    SB_LUT4 mult_11_add_1225_19_lut (.I0(GND_net), .I1(n9339[16]), .I2(GND_net), 
            .I3(n39625), .O(n155[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5789_18 (.CI(n39514), .I0(n15209[15]), .I1(GND_net), 
            .CO(n39515));
    SB_LUT4 mult_11_i414_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n615_adj_4647));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i271_2_lut (.I0(\Kp[5] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n402_adj_4648));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i271_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i3_1_lut (.I0(PWMLimit[2]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[2]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i3_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i649_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n965_adj_4649));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i649_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20707_2_lut (.I0(n1[2]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[2]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20707_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_710_10_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [8]), 
            .I2(n3616[8]), .I3(n39143), .O(\PID_CONTROLLER.integral_23__N_3572 [8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_12_lut (.I0(GND_net), .I1(setpoint[10]), .I2(motor_state[10]), 
            .I3(n39219), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_710_10 (.CI(n39143), .I0(\PID_CONTROLLER.integral [8]), 
            .I1(n3616[8]), .CO(n39144));
    SB_LUT4 add_710_9_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [7]), 
            .I2(n3616[7]), .I3(n39142), .O(\PID_CONTROLLER.integral_23__N_3572 [7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6071_2_lut (.I0(GND_net), .I1(n53_adj_4650), .I2(n122_adj_4651), 
            .I3(GND_net), .O(n18812[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6071_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6071_2 (.CI(GND_net), .I0(n53_adj_4650), .I1(n122_adj_4651), 
            .CO(n39409));
    SB_LUT4 mult_10_i320_2_lut (.I0(\Kp[6] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n475_adj_4652));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i320_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_12 (.CI(n39219), .I0(setpoint[10]), .I1(motor_state[10]), 
            .CO(n39220));
    SB_LUT4 add_6003_9_lut (.I0(GND_net), .I1(n18325[6]), .I2(n621_adj_4653), 
            .I3(n39731), .O(n18084[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6003_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5789_17_lut (.I0(GND_net), .I1(n15209[14]), .I2(GND_net), 
            .I3(n39513), .O(n14525[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5789_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_710_9 (.CI(n39142), .I0(\PID_CONTROLLER.integral [7]), 
            .I1(n3616[7]), .CO(n39143));
    SB_CARRY mult_11_add_1225_19 (.CI(n39625), .I0(n9339[16]), .I1(GND_net), 
            .CO(n39626));
    SB_LUT4 i20706_2_lut (.I0(n1[3]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[3]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20706_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5944_14_lut (.I0(GND_net), .I1(n17629[11]), .I2(n980_adj_4654), 
            .I3(n39408), .O(n17265[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5944_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5944_13_lut (.I0(GND_net), .I1(n17629[10]), .I2(n907_adj_4655), 
            .I3(n39407), .O(n17265[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5944_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_11_lut (.I0(GND_net), .I1(setpoint[9]), .I2(motor_state[9]), 
            .I3(n39218), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_11 (.CI(n39218), .I0(setpoint[9]), .I1(motor_state[9]), 
            .CO(n39219));
    SB_CARRY add_5944_13 (.CI(n39407), .I0(n17629[10]), .I1(n907_adj_4655), 
            .CO(n39408));
    SB_LUT4 add_710_8_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [6]), 
            .I2(n3616[6]), .I3(n39141), .O(\PID_CONTROLLER.integral_23__N_3572 [6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5732_4_lut (.I0(GND_net), .I1(n14164[1]), .I2(n229_adj_4656), 
            .I3(n39957), .O(n13364[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6003_9 (.CI(n39731), .I0(n18325[6]), .I1(n621_adj_4653), 
            .CO(n39732));
    SB_CARRY add_5789_17 (.CI(n39513), .I0(n15209[14]), .I1(GND_net), 
            .CO(n39514));
    SB_LUT4 i20705_2_lut (.I0(n1[4]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[4]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20705_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_18_lut (.I0(GND_net), .I1(n9339[15]), .I2(GND_net), 
            .I3(n39624), .O(n155[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i463_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n688_adj_4658));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i463_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_710_8 (.CI(n39141), .I0(\PID_CONTROLLER.integral [6]), 
            .I1(n3616[6]), .CO(n39142));
    SB_LUT4 sub_3_add_2_10_lut (.I0(GND_net), .I1(setpoint[8]), .I2(motor_state[8]), 
            .I3(n39217), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_10 (.CI(n39217), .I0(setpoint[8]), .I1(motor_state[8]), 
            .CO(n39218));
    SB_LUT4 add_5789_16_lut (.I0(GND_net), .I1(n15209[13]), .I2(n1111_adj_4659), 
            .I3(n39512), .O(n14525[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5789_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5732_4 (.CI(n39957), .I0(n14164[1]), .I1(n229_adj_4656), 
            .CO(n39958));
    SB_LUT4 add_710_7_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [5]), 
            .I2(n3616[5]), .I3(n39140), .O(\PID_CONTROLLER.integral_23__N_3572 [5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_710_7 (.CI(n39140), .I0(\PID_CONTROLLER.integral [5]), 
            .I1(n3616[5]), .CO(n39141));
    SB_LUT4 add_5944_12_lut (.I0(GND_net), .I1(n17629[9]), .I2(n834_adj_4660), 
            .I3(n39406), .O(n17265[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5944_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5957_9 (.CI(n39837), .I0(n17797[6]), .I1(n615), .CO(n39838));
    SB_LUT4 add_6003_8_lut (.I0(GND_net), .I1(n18325[5]), .I2(n548_adj_4661), 
            .I3(n39730), .O(n18084[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6003_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5732_3_lut (.I0(GND_net), .I1(n14164[0]), .I2(n156_adj_4662), 
            .I3(n39956), .O(n13364[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5957_8_lut (.I0(GND_net), .I1(n17797[5]), .I2(n542_adj_4663), 
            .I3(n39836), .O(n17460[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i126_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n186));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i126_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5789_16 (.CI(n39512), .I0(n15209[13]), .I1(n1111_adj_4659), 
            .CO(n39513));
    SB_LUT4 add_5789_15_lut (.I0(GND_net), .I1(n15209[12]), .I2(n1038_adj_4664), 
            .I3(n39511), .O(n14525[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5789_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5944_12 (.CI(n39406), .I0(n17629[9]), .I1(n834_adj_4660), 
            .CO(n39407));
    SB_CARRY mult_11_add_1225_18 (.CI(n39624), .I0(n9339[15]), .I1(GND_net), 
            .CO(n39625));
    SB_CARRY add_6003_8 (.CI(n39730), .I0(n18325[5]), .I1(n548_adj_4661), 
            .CO(n39731));
    SB_LUT4 add_5944_11_lut (.I0(GND_net), .I1(n17629[8]), .I2(n761_adj_4665), 
            .I3(n39405), .O(n17265[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5944_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5944_11 (.CI(n39405), .I0(n17629[8]), .I1(n761_adj_4665), 
            .CO(n39406));
    SB_CARRY add_5789_15 (.CI(n39511), .I0(n15209[12]), .I1(n1038_adj_4664), 
            .CO(n39512));
    SB_LUT4 sub_3_add_2_9_lut (.I0(GND_net), .I1(setpoint[7]), .I2(motor_state[7]), 
            .I3(n39216), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_9 (.CI(n39216), .I0(setpoint[7]), .I1(motor_state[7]), 
            .CO(n39217));
    SB_CARRY add_5957_8 (.CI(n39836), .I0(n17797[5]), .I1(n542_adj_4663), 
            .CO(n39837));
    SB_LUT4 add_5944_10_lut (.I0(GND_net), .I1(n17629[7]), .I2(n688_adj_4658), 
            .I3(n39404), .O(n17265[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5944_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_710_6_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [4]), 
            .I2(n3616[4]), .I3(n39139), .O(\PID_CONTROLLER.integral_23__N_3572 [4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5944_10 (.CI(n39404), .I0(n17629[7]), .I1(n688_adj_4658), 
            .CO(n39405));
    SB_CARRY add_710_6 (.CI(n39139), .I0(\PID_CONTROLLER.integral [4]), 
            .I1(n3616[4]), .CO(n39140));
    SB_LUT4 add_710_5_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [3]), 
            .I2(n3616[3]), .I3(n39138), .O(\PID_CONTROLLER.integral_23__N_3572 [3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6003_7_lut (.I0(GND_net), .I1(n18325[4]), .I2(n475_adj_4652), 
            .I3(n39729), .O(n18084[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6003_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_8_lut (.I0(GND_net), .I1(setpoint[6]), .I2(motor_state[6]), 
            .I3(n39215), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_8 (.CI(n39215), .I0(setpoint[6]), .I1(motor_state[6]), 
            .CO(n39216));
    SB_LUT4 mult_10_i310_2_lut (.I0(\Kp[6] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n460));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i508_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n755));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i508_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_6003_7 (.CI(n39729), .I0(n18325[4]), .I1(n475_adj_4652), 
            .CO(n39730));
    SB_CARRY add_710_5 (.CI(n39138), .I0(\PID_CONTROLLER.integral [3]), 
            .I1(n3616[3]), .CO(n39139));
    SB_LUT4 add_710_4_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [2]), 
            .I2(n3616[2]), .I3(n39137), .O(\PID_CONTROLLER.integral_23__N_3572 [2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_17_lut (.I0(GND_net), .I1(n9339[14]), .I2(GND_net), 
            .I3(n39623), .O(n155[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5789_14_lut (.I0(GND_net), .I1(n15209[11]), .I2(n965_adj_4649), 
            .I3(n39510), .O(n14525[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5789_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i4_1_lut (.I0(PWMLimit[3]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[3]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i4_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 add_6003_6_lut (.I0(GND_net), .I1(n18325[3]), .I2(n402_adj_4648), 
            .I3(n39728), .O(n18084[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6003_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5944_9_lut (.I0(GND_net), .I1(n17629[6]), .I2(n615_adj_4647), 
            .I3(n39403), .O(n17265[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5944_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_710_4 (.CI(n39137), .I0(\PID_CONTROLLER.integral [2]), 
            .I1(n3616[2]), .CO(n39138));
    SB_CARRY mult_11_add_1225_17 (.CI(n39623), .I0(n9339[14]), .I1(GND_net), 
            .CO(n39624));
    SB_CARRY add_6003_6 (.CI(n39728), .I0(n18325[3]), .I1(n402_adj_4648), 
            .CO(n39729));
    SB_LUT4 mult_11_add_1225_16_lut (.I0(GND_net), .I1(n9339[13]), .I2(n1096_adj_4643), 
            .I3(n39622), .O(n155[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_16 (.CI(n39622), .I0(n9339[13]), .I1(n1096_adj_4643), 
            .CO(n39623));
    SB_LUT4 mult_11_add_1225_15_lut (.I0(GND_net), .I1(n9339[12]), .I2(n1023_adj_4642), 
            .I3(n39621), .O(n155[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5789_14 (.CI(n39510), .I0(n15209[11]), .I1(n965_adj_4649), 
            .CO(n39511));
    SB_LUT4 add_5789_13_lut (.I0(GND_net), .I1(n15209[10]), .I2(n892_adj_4641), 
            .I3(n39509), .O(n14525[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5789_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_7_lut (.I0(GND_net), .I1(setpoint[5]), .I2(motor_state[5]), 
            .I3(n39214), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5944_9 (.CI(n39403), .I0(n17629[6]), .I1(n615_adj_4647), 
            .CO(n39404));
    SB_LUT4 add_5944_8_lut (.I0(GND_net), .I1(n17629[5]), .I2(n542), .I3(n39402), 
            .O(n17265[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5944_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5789_13 (.CI(n39509), .I0(n15209[10]), .I1(n892_adj_4641), 
            .CO(n39510));
    SB_CARRY sub_3_add_2_7 (.CI(n39214), .I0(setpoint[5]), .I1(motor_state[5]), 
            .CO(n39215));
    SB_CARRY add_5944_8 (.CI(n39402), .I0(n17629[5]), .I1(n542), .CO(n39403));
    SB_LUT4 add_6003_5_lut (.I0(GND_net), .I1(n18325[2]), .I2(n329_adj_4639), 
            .I3(n39727), .O(n18084[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6003_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_15 (.CI(n39621), .I0(n9339[12]), .I1(n1023_adj_4642), 
            .CO(n39622));
    SB_LUT4 add_710_3_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [1]), 
            .I2(n3616[1]), .I3(n39136), .O(\PID_CONTROLLER.integral_23__N_3572 [1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5789_12_lut (.I0(GND_net), .I1(n15209[9]), .I2(n819_adj_4638), 
            .I3(n39508), .O(n14525[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5789_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5732_3 (.CI(n39956), .I0(n14164[0]), .I1(n156_adj_4662), 
            .CO(n39957));
    SB_LUT4 add_5944_7_lut (.I0(GND_net), .I1(n17629[4]), .I2(n469_adj_4637), 
            .I3(n39401), .O(n17265[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5944_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_710_3 (.CI(n39136), .I0(\PID_CONTROLLER.integral [1]), 
            .I1(n3616[1]), .CO(n39137));
    SB_CARRY add_5944_7 (.CI(n39401), .I0(n17629[4]), .I1(n469_adj_4637), 
            .CO(n39402));
    SB_LUT4 sub_3_add_2_6_lut (.I0(GND_net), .I1(setpoint[4]), .I2(motor_state[4]), 
            .I3(n39213), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5944_6_lut (.I0(GND_net), .I1(n17629[3]), .I2(n396_adj_4622), 
            .I3(n39400), .O(n17265[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5944_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_710_2_lut (.I0(GND_net), .I1(\PID_CONTROLLER.integral [0]), 
            .I2(n3616[0]), .I3(GND_net), .O(\PID_CONTROLLER.integral_23__N_3572 [0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_710_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_6 (.CI(n39213), .I0(setpoint[4]), .I1(motor_state[4]), 
            .CO(n39214));
    SB_LUT4 add_5957_7_lut (.I0(GND_net), .I1(n17797[4]), .I2(n469), .I3(n39835), 
            .O(n17460[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5944_6 (.CI(n39400), .I0(n17629[3]), .I1(n396_adj_4622), 
            .CO(n39401));
    SB_CARRY add_710_2 (.CI(GND_net), .I0(\PID_CONTROLLER.integral [0]), 
            .I1(n3616[0]), .CO(n39136));
    SB_CARRY add_5957_7 (.CI(n39835), .I0(n17797[4]), .I1(n469), .CO(n39836));
    SB_LUT4 mult_11_i512_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n761_adj_4665));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i698_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1038_adj_4664));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_5_lut (.I0(GND_net), .I1(setpoint[3]), .I2(motor_state[3]), 
            .I3(n39212), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_25_lut (.I0(GND_net), .I1(n9363[0]), .I2(n8832[0]), 
            .I3(n39135), .O(duty_23__N_3672[23])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i365_2_lut (.I0(\Kp[7] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n542_adj_4663));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i365_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5957_6_lut (.I0(GND_net), .I1(n17797[3]), .I2(n396), .I3(n39834), 
            .O(n17460[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5789_12 (.CI(n39508), .I0(n15209[9]), .I1(n819_adj_4638), 
            .CO(n39509));
    SB_LUT4 mult_10_i106_2_lut (.I0(\Kp[2] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n156_adj_4662));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i106_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_3_add_2_5 (.CI(n39212), .I0(setpoint[3]), .I1(motor_state[3]), 
            .CO(n39213));
    SB_LUT4 add_12_24_lut (.I0(GND_net), .I1(n106[22]), .I2(n155[22]), 
            .I3(n39134), .O(duty_23__N_3672[22])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_24_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5944_5_lut (.I0(GND_net), .I1(n17629[2]), .I2(n323_adj_4617), 
            .I3(n39399), .O(n17265[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5944_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_4_lut (.I0(GND_net), .I1(setpoint[2]), .I2(motor_state[2]), 
            .I3(n39211), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_4 (.CI(n39211), .I0(setpoint[2]), .I1(motor_state[2]), 
            .CO(n39212));
    SB_CARRY add_12_24 (.CI(n39134), .I0(n106[22]), .I1(n155[22]), .CO(n39135));
    SB_LUT4 mult_11_i175_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n259));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i175_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5732_2_lut (.I0(GND_net), .I1(n14_adj_4616), .I2(n83_adj_4615), 
            .I3(GND_net), .O(n13364[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5732_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i369_2_lut (.I0(\Kp[7] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n548_adj_4661));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i369_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i561_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n834_adj_4660));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i249_2_lut (.I0(\Kp[5] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n369));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i249_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20704_2_lut (.I0(n1[5]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[5]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i747_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n1111_adj_4659));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i747_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 sub_3_add_2_3_lut (.I0(GND_net), .I1(setpoint[1]), .I2(motor_state[1]), 
            .I3(n39210), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_23_lut (.I0(GND_net), .I1(n106[21]), .I2(n155[21]), 
            .I3(n39133), .O(duty_23__N_3672[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6003_5 (.CI(n39727), .I0(n18325[2]), .I1(n329_adj_4639), 
            .CO(n39728));
    SB_CARRY add_5944_5 (.CI(n39399), .I0(n17629[2]), .I1(n323_adj_4617), 
            .CO(n39400));
    SB_LUT4 add_5789_11_lut (.I0(GND_net), .I1(n15209[8]), .I2(n746_adj_4614), 
            .I3(n39507), .O(n14525[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5789_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_3 (.CI(n39210), .I0(setpoint[1]), .I1(motor_state[1]), 
            .CO(n39211));
    SB_CARRY add_5732_2 (.CI(GND_net), .I0(n14_adj_4616), .I1(n83_adj_4615), 
            .CO(n39956));
    SB_LUT4 add_5771_20_lut (.I0(GND_net), .I1(n14885[17]), .I2(GND_net), 
            .I3(n39955), .O(n14164[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5944_4_lut (.I0(GND_net), .I1(n17629[1]), .I2(n250_adj_4613), 
            .I3(n39398), .O(n17265[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5944_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5771_19_lut (.I0(GND_net), .I1(n14885[16]), .I2(GND_net), 
            .I3(n39954), .O(n14164[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_23 (.CI(n39133), .I0(n106[21]), .I1(n155[21]), .CO(n39134));
    SB_CARRY add_5944_4 (.CI(n39398), .I0(n17629[1]), .I1(n250_adj_4613), 
            .CO(n39399));
    SB_CARRY add_5789_11 (.CI(n39507), .I0(n15209[8]), .I1(n746_adj_4614), 
            .CO(n39508));
    SB_LUT4 mult_11_i557_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n828));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i557_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5944_3_lut (.I0(GND_net), .I1(n17629[0]), .I2(n177_adj_4612), 
            .I3(n39397), .O(n17265[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5944_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i547_2_lut (.I0(\Ki[11] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n813_adj_4441));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i547_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i224_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n332));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i224_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i596_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n886_adj_4439));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i596_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i606_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n901));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i606_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_14_lut (.I0(GND_net), .I1(n9339[11]), .I2(n950_adj_4611), 
            .I3(n39620), .O(n155[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_3_add_2_2_lut (.I0(GND_net), .I1(setpoint[0]), .I2(motor_state[0]), 
            .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_3_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_22_lut (.I0(GND_net), .I1(n106[20]), .I2(n155[20]), 
            .I3(n39132), .O(duty_23__N_3672[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5789_10_lut (.I0(GND_net), .I1(n15209[7]), .I2(n673_adj_4610), 
            .I3(n39506), .O(n14525[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5789_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_3_add_2_2 (.CI(VCC_net), .I0(setpoint[0]), .I1(motor_state[0]), 
            .CO(n39210));
    SB_CARRY add_5789_10 (.CI(n39506), .I0(n15209[7]), .I1(n673_adj_4610), 
            .CO(n39507));
    SB_LUT4 unary_minus_16_inv_0_i5_1_lut (.I0(PWMLimit[4]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[4]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i5_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5957_6 (.CI(n39834), .I0(n17797[3]), .I1(n396), .CO(n39835));
    SB_LUT4 mult_11_i655_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n974));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i655_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i273_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n405));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i273_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_22 (.CI(n39132), .I0(n106[20]), .I1(n155[20]), .CO(n39133));
    SB_CARRY add_5771_19 (.CI(n39954), .I0(n14885[16]), .I1(GND_net), 
            .CO(n39955));
    SB_LUT4 add_12_21_lut (.I0(GND_net), .I1(n106[19]), .I2(n155[19]), 
            .I3(n39131), .O(duty_23__N_3672[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_14 (.CI(n39620), .I0(n9339[11]), .I1(n950_adj_4611), 
            .CO(n39621));
    SB_CARRY add_5944_3 (.CI(n39397), .I0(n17629[0]), .I1(n177_adj_4612), 
            .CO(n39398));
    SB_LUT4 add_5789_9_lut (.I0(GND_net), .I1(n15209[6]), .I2(n600_adj_4609), 
            .I3(n39505), .O(n14525[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5789_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5957_5_lut (.I0(GND_net), .I1(n17797[2]), .I2(n323), .I3(n39833), 
            .O(n17460[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5789_9 (.CI(n39505), .I0(n15209[6]), .I1(n600_adj_4609), 
            .CO(n39506));
    SB_LUT4 add_5771_18_lut (.I0(GND_net), .I1(n14885[15]), .I2(GND_net), 
            .I3(n39953), .O(n14164[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5944_2_lut (.I0(GND_net), .I1(n35_adj_4608), .I2(n104_adj_4607), 
            .I3(GND_net), .O(n17265[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5944_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5957_5 (.CI(n39833), .I0(n17797[2]), .I1(n323), .CO(n39834));
    SB_CARRY add_12_21 (.CI(n39131), .I0(n106[19]), .I1(n155[19]), .CO(n39132));
    SB_CARRY add_5944_2 (.CI(GND_net), .I0(n35_adj_4608), .I1(n104_adj_4607), 
            .CO(n39397));
    SB_LUT4 add_12_20_lut (.I0(GND_net), .I1(n106[18]), .I2(n155[18]), 
            .I3(n39130), .O(duty_23__N_3672[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i645_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n959_adj_4431));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i645_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_add_1225_13_lut (.I0(GND_net), .I1(n9339[10]), .I2(n877_adj_4606), 
            .I3(n39619), .O(n155[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6003_4_lut (.I0(GND_net), .I1(n18325[1]), .I2(n256_adj_4605), 
            .I3(n39726), .O(n18084[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6003_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5789_8_lut (.I0(GND_net), .I1(n15209[5]), .I2(n527_adj_4604), 
            .I3(n39504), .O(n14525[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5789_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_13 (.CI(n39619), .I0(n9339[10]), .I1(n877_adj_4606), 
            .CO(n39620));
    SB_LUT4 mult_11_i694_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1032_adj_4427));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i694_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5789_8 (.CI(n39504), .I0(n15209[5]), .I1(n527_adj_4604), 
            .CO(n39505));
    SB_CARRY add_12_20 (.CI(n39130), .I0(n106[18]), .I1(n155[18]), .CO(n39131));
    SB_LUT4 add_5969_13_lut (.I0(GND_net), .I1(n17941[10]), .I2(n910_adj_4603), 
            .I3(n39396), .O(n17629[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5969_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6003_4 (.CI(n39726), .I0(n18325[1]), .I1(n256_adj_4605), 
            .CO(n39727));
    SB_LUT4 add_5789_7_lut (.I0(GND_net), .I1(n15209[4]), .I2(n454_adj_4602), 
            .I3(n39503), .O(n14525[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5789_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5789_7 (.CI(n39503), .I0(n15209[4]), .I1(n454_adj_4602), 
            .CO(n39504));
    SB_LUT4 add_5969_12_lut (.I0(GND_net), .I1(n17941[9]), .I2(n837_adj_4601), 
            .I3(n39395), .O(n17629[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5969_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5969_12 (.CI(n39395), .I0(n17941[9]), .I1(n837_adj_4601), 
            .CO(n39396));
    SB_LUT4 add_12_19_lut (.I0(GND_net), .I1(n106[17]), .I2(n155[17]), 
            .I3(n39129), .O(duty_23__N_3672[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i704_2_lut (.I0(\Ki[14] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1047));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i704_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6003_3_lut (.I0(GND_net), .I1(n18325[0]), .I2(n183), .I3(n39725), 
            .O(n18084[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6003_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_12_lut (.I0(GND_net), .I1(n9339[9]), .I2(n804_adj_4600), 
            .I3(n39618), .O(n155[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_19 (.CI(n39129), .I0(n106[17]), .I1(n155[17]), .CO(n39130));
    SB_LUT4 add_5957_4_lut (.I0(GND_net), .I1(n17797[1]), .I2(n250), .I3(n39832), 
            .O(n17460[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6003_3 (.CI(n39725), .I0(n18325[0]), .I1(n183), .CO(n39726));
    SB_LUT4 add_5789_6_lut (.I0(GND_net), .I1(n15209[3]), .I2(n381_adj_4599), 
            .I3(n39502), .O(n14525[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5789_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_12 (.CI(n39618), .I0(n9339[9]), .I1(n804_adj_4600), 
            .CO(n39619));
    SB_LUT4 add_6003_2_lut (.I0(GND_net), .I1(n41_adj_4598), .I2(n110), 
            .I3(GND_net), .O(n18084[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6003_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5771_18 (.CI(n39953), .I0(n14885[15]), .I1(GND_net), 
            .CO(n39954));
    SB_LUT4 mult_11_add_1225_11_lut (.I0(GND_net), .I1(n9339[8]), .I2(n731_adj_4597), 
            .I3(n39617), .O(n155[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_11 (.CI(n39617), .I0(n9339[8]), .I1(n731_adj_4597), 
            .CO(n39618));
    SB_LUT4 add_5771_17_lut (.I0(GND_net), .I1(n14885[14]), .I2(GND_net), 
            .I3(n39952), .O(n14164[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5789_6 (.CI(n39502), .I0(n15209[3]), .I1(n381_adj_4599), 
            .CO(n39503));
    SB_LUT4 add_5789_5_lut (.I0(GND_net), .I1(n15209[2]), .I2(n308_adj_4596), 
            .I3(n39501), .O(n14525[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5789_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6003_2 (.CI(GND_net), .I0(n41_adj_4598), .I1(n110), .CO(n39725));
    SB_CARRY add_5957_4 (.CI(n39832), .I0(n17797[1]), .I1(n250), .CO(n39833));
    SB_CARRY add_5789_5 (.CI(n39501), .I0(n15209[2]), .I1(n308_adj_4596), 
            .CO(n39502));
    SB_LUT4 add_5789_4_lut (.I0(GND_net), .I1(n15209[1]), .I2(n235_adj_4595), 
            .I3(n39500), .O(n14525[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5789_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_10_lut (.I0(GND_net), .I1(n9339[7]), .I2(n658_adj_4594), 
            .I3(n39616), .O(n155[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_10 (.CI(n39616), .I0(n9339[7]), .I1(n658_adj_4594), 
            .CO(n39617));
    SB_LUT4 mult_10_i359_2_lut (.I0(\Kp[7] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n533));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i359_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5789_4 (.CI(n39500), .I0(n15209[1]), .I1(n235_adj_4595), 
            .CO(n39501));
    SB_LUT4 mult_11_add_1225_9_lut (.I0(GND_net), .I1(n9339[6]), .I2(n585_adj_4593), 
            .I3(n39615), .O(n155[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_18_lut (.I0(GND_net), .I1(n106[16]), .I2(n155[16]), 
            .I3(n39128), .O(duty_23__N_3672[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5969_11_lut (.I0(GND_net), .I1(n17941[8]), .I2(n764_adj_4592), 
            .I3(n39394), .O(n17629[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5969_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5789_3_lut (.I0(GND_net), .I1(n15209[0]), .I2(n162_adj_4591), 
            .I3(n39499), .O(n14525[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5789_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5969_11 (.CI(n39394), .I0(n17941[8]), .I1(n764_adj_4592), 
            .CO(n39395));
    SB_LUT4 add_5969_10_lut (.I0(GND_net), .I1(n17941[7]), .I2(n691_adj_4590), 
            .I3(n39393), .O(n17629[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5969_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_inv_0_i6_1_lut (.I0(PWMLimit[5]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[5]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i6_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i743_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n1105_adj_4423));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i743_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5789_3 (.CI(n39499), .I0(n15209[0]), .I1(n162_adj_4591), 
            .CO(n39500));
    SB_CARRY add_5969_10 (.CI(n39393), .I0(n17941[7]), .I1(n691_adj_4590), 
            .CO(n39394));
    SB_LUT4 add_5957_3_lut (.I0(GND_net), .I1(n17797[0]), .I2(n177), .I3(n39831), 
            .O(n17460[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5771_17 (.CI(n39952), .I0(n14885[14]), .I1(GND_net), 
            .CO(n39953));
    SB_CARRY mult_11_add_1225_9 (.CI(n39615), .I0(n9339[6]), .I1(n585_adj_4593), 
            .CO(n39616));
    SB_CARRY add_5957_3 (.CI(n39831), .I0(n17797[0]), .I1(n177), .CO(n39832));
    SB_LUT4 add_5771_16_lut (.I0(GND_net), .I1(n14885[13]), .I2(n1108_adj_4589), 
            .I3(n39951), .O(n14164[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5969_9_lut (.I0(GND_net), .I1(n17941[6]), .I2(n618_adj_4588), 
            .I3(n39392), .O(n17629[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5969_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5957_2_lut (.I0(GND_net), .I1(n35_adj_4587), .I2(n104), 
            .I3(GND_net), .O(n17460[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5957_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5789_2_lut (.I0(GND_net), .I1(n20_adj_4586), .I2(n89_adj_4585), 
            .I3(GND_net), .O(n14525[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5789_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_18 (.CI(n39128), .I0(n106[16]), .I1(n155[16]), .CO(n39129));
    SB_LUT4 mult_11_add_1225_8_lut (.I0(GND_net), .I1(n9339[5]), .I2(n512_adj_4584), 
            .I3(n39614), .O(n155[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5789_2 (.CI(GND_net), .I0(n20_adj_4586), .I1(n89_adj_4585), 
            .CO(n39499));
    SB_CARRY mult_11_add_1225_8 (.CI(n39614), .I0(n9339[5]), .I1(n512_adj_4584), 
            .CO(n39615));
    SB_LUT4 add_6041_10_lut (.I0(GND_net), .I1(n18685[7]), .I2(n700_adj_4583), 
            .I3(n39498), .O(n18524[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_7_lut (.I0(GND_net), .I1(n9339[4]), .I2(n439_adj_4582), 
            .I3(n39613), .O(n155[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i322_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n478));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i322_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i7_1_lut (.I0(PWMLimit[6]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[6]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i7_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5771_16 (.CI(n39951), .I0(n14885[13]), .I1(n1108_adj_4589), 
            .CO(n39952));
    SB_LUT4 add_5771_15_lut (.I0(GND_net), .I1(n14885[12]), .I2(n1035_adj_4581), 
            .I3(n39950), .O(n14164[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_17_lut (.I0(GND_net), .I1(n106[15]), .I2(n155[15]), 
            .I3(n39127), .O(duty_23__N_3672[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_7 (.CI(n39613), .I0(n9339[4]), .I1(n439_adj_4582), 
            .CO(n39614));
    SB_CARRY add_5969_9 (.CI(n39392), .I0(n17941[6]), .I1(n618_adj_4588), 
            .CO(n39393));
    SB_LUT4 add_5969_8_lut (.I0(GND_net), .I1(n17941[5]), .I2(n545_adj_4580), 
            .I3(n39391), .O(n17629[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5969_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6041_9_lut (.I0(GND_net), .I1(n18685[6]), .I2(n627_adj_4579), 
            .I3(n39497), .O(n18524[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5969_8 (.CI(n39391), .I0(n17941[5]), .I1(n545_adj_4580), 
            .CO(n39392));
    SB_LUT4 mult_11_add_1225_6_lut (.I0(GND_net), .I1(n9339[3]), .I2(n366_adj_4578), 
            .I3(n39612), .O(n155[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5957_2 (.CI(GND_net), .I0(n35_adj_4587), .I1(n104), .CO(n39831));
    SB_CARRY mult_11_add_1225_6 (.CI(n39612), .I0(n9339[3]), .I1(n366_adj_4578), 
            .CO(n39613));
    SB_LUT4 add_5969_7_lut (.I0(GND_net), .I1(n17941[4]), .I2(n472_adj_4577), 
            .I3(n39390), .O(n17629[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5969_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_5_lut (.I0(GND_net), .I1(n9339[2]), .I2(n293_adj_4576), 
            .I3(n39611), .O(n155[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5771_15 (.CI(n39950), .I0(n14885[12]), .I1(n1035_adj_4581), 
            .CO(n39951));
    SB_CARRY mult_11_add_1225_5 (.CI(n39611), .I0(n9339[2]), .I1(n293_adj_4576), 
            .CO(n39612));
    SB_LUT4 add_5771_14_lut (.I0(GND_net), .I1(n14885[11]), .I2(n962_adj_4575), 
            .I3(n39949), .O(n14164[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5981_13_lut (.I0(GND_net), .I1(n18084[10]), .I2(n910), 
            .I3(n39830), .O(n17797[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5981_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5981_12_lut (.I0(GND_net), .I1(n18084[9]), .I2(n837), 
            .I3(n39829), .O(n17797[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5981_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6041_9 (.CI(n39497), .I0(n18685[6]), .I1(n627_adj_4579), 
            .CO(n39498));
    SB_CARRY add_5969_7 (.CI(n39390), .I0(n17941[4]), .I1(n472_adj_4577), 
            .CO(n39391));
    SB_CARRY add_5771_14 (.CI(n39949), .I0(n14885[11]), .I1(n962_adj_4575), 
            .CO(n39950));
    SB_LUT4 add_5969_6_lut (.I0(GND_net), .I1(n17941[3]), .I2(n399_adj_4574), 
            .I3(n39389), .O(n17629[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5969_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5981_12 (.CI(n39829), .I0(n18084[9]), .I1(n837), .CO(n39830));
    SB_CARRY add_5969_6 (.CI(n39389), .I0(n17941[3]), .I1(n399_adj_4574), 
            .CO(n39390));
    SB_LUT4 add_5981_11_lut (.I0(GND_net), .I1(n18084[8]), .I2(n764), 
            .I3(n39828), .O(n17797[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5981_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5771_13_lut (.I0(GND_net), .I1(n14885[10]), .I2(n889_adj_4573), 
            .I3(n39948), .O(n14164[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5771_13 (.CI(n39948), .I0(n14885[10]), .I1(n889_adj_4573), 
            .CO(n39949));
    SB_CARRY add_5981_11 (.CI(n39828), .I0(n18084[8]), .I1(n764), .CO(n39829));
    SB_LUT4 add_5771_12_lut (.I0(GND_net), .I1(n14885[9]), .I2(n816_adj_4572), 
            .I3(n39947), .O(n14164[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5771_12 (.CI(n39947), .I0(n14885[9]), .I1(n816_adj_4572), 
            .CO(n39948));
    SB_LUT4 add_6041_8_lut (.I0(GND_net), .I1(n18685[5]), .I2(n554_adj_4571), 
            .I3(n39496), .O(n18524[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5981_10_lut (.I0(GND_net), .I1(n18084[7]), .I2(n691), 
            .I3(n39827), .O(n17797[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5981_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5771_11_lut (.I0(GND_net), .I1(n14885[8]), .I2(n743_adj_4570), 
            .I3(n39946), .O(n14164[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5981_10 (.CI(n39827), .I0(n18084[7]), .I1(n691), .CO(n39828));
    SB_CARRY add_5771_11 (.CI(n39946), .I0(n14885[8]), .I1(n743_adj_4570), 
            .CO(n39947));
    SB_LUT4 mult_10_i408_2_lut (.I0(\Kp[8] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n606));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i753_2_lut (.I0(\Ki[15] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n1120));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i753_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_17 (.CI(n39127), .I0(n106[15]), .I1(n155[15]), .CO(n39128));
    SB_LUT4 add_5981_9_lut (.I0(GND_net), .I1(n18084[6]), .I2(n618), .I3(n39826), 
            .O(n17797[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5981_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5771_10_lut (.I0(GND_net), .I1(n14885[7]), .I2(n670), 
            .I3(n39945), .O(n14164[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5771_10 (.CI(n39945), .I0(n14885[7]), .I1(n670), .CO(n39946));
    SB_CARRY add_6041_8 (.CI(n39496), .I0(n18685[5]), .I1(n554_adj_4571), 
            .CO(n39497));
    SB_LUT4 add_12_16_lut (.I0(GND_net), .I1(n106[14]), .I2(n155[14]), 
            .I3(n39126), .O(duty_23__N_3672[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_4_lut (.I0(GND_net), .I1(n9339[1]), .I2(n220_adj_4569), 
            .I3(n39610), .O(n155[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_16 (.CI(n39126), .I0(n106[14]), .I1(n155[14]), .CO(n39127));
    SB_LUT4 add_5771_9_lut (.I0(GND_net), .I1(n14885[6]), .I2(n597), .I3(n39944), 
            .O(n14164[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_4 (.CI(n39610), .I0(n9339[1]), .I1(n220_adj_4569), 
            .CO(n39611));
    SB_CARRY add_5981_9 (.CI(n39826), .I0(n18084[6]), .I1(n618), .CO(n39827));
    SB_LUT4 unary_minus_16_inv_0_i8_1_lut (.I0(PWMLimit[7]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[7]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i8_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i371_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n551));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i371_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5771_9 (.CI(n39944), .I0(n14885[6]), .I1(n597), .CO(n39945));
    SB_LUT4 add_5981_8_lut (.I0(GND_net), .I1(n18084[5]), .I2(n545), .I3(n39825), 
            .O(n17797[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5981_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6041_7_lut (.I0(GND_net), .I1(n18685[4]), .I2(n481_adj_4568), 
            .I3(n39495), .O(n18524[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_add_1225_3_lut (.I0(GND_net), .I1(n9339[0]), .I2(n147), 
            .I3(n39609), .O(n155[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6041_7 (.CI(n39495), .I0(n18685[4]), .I1(n481_adj_4568), 
            .CO(n39496));
    SB_LUT4 mult_10_i81_2_lut (.I0(\Kp[1] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n119));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i81_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i34_2_lut (.I0(\Kp[0] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n50));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i34_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i53_2_lut (.I0(\Kp[1] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n77_adj_4380));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i53_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i6_2_lut (.I0(\Kp[0] ), .I1(n1[2]), .I2(GND_net), 
            .I3(GND_net), .O(n8_adj_4379));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i6_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i420_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n624));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i420_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5771_8_lut (.I0(GND_net), .I1(n14885[5]), .I2(n524), .I3(n39943), 
            .O(n14164[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_3 (.CI(n39609), .I0(n9339[0]), .I1(n147), 
            .CO(n39610));
    SB_CARRY add_5771_8 (.CI(n39943), .I0(n14885[5]), .I1(n524), .CO(n39944));
    SB_CARRY add_5981_8 (.CI(n39825), .I0(n18084[5]), .I1(n545), .CO(n39826));
    SB_LUT4 mult_11_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4567), .I2(n74), 
            .I3(GND_net), .O(n155[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_11_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i130_2_lut (.I0(\Kp[2] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n192));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i130_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i469_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n697));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i469_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6041_6_lut (.I0(GND_net), .I1(n18685[3]), .I2(n408_adj_4566), 
            .I3(n39494), .O(n18524[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_11_add_1225_2 (.CI(GND_net), .I0(n5_adj_4567), .I1(n74), 
            .CO(n39609));
    SB_LUT4 add_5969_5_lut (.I0(GND_net), .I1(n17941[2]), .I2(n326_adj_4565), 
            .I3(n39388), .O(n17629[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5969_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5771_7_lut (.I0(GND_net), .I1(n14885[4]), .I2(n451), .I3(n39942), 
            .O(n14164[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5981_7_lut (.I0(GND_net), .I1(n18084[4]), .I2(n472), .I3(n39824), 
            .O(n17797[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5981_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_15_lut (.I0(GND_net), .I1(n106[13]), .I2(n155[13]), 
            .I3(n39125), .O(duty_23__N_3672[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4054_23_lut (.I0(GND_net), .I1(n11628[20]), .I2(GND_net), 
            .I3(n39608), .O(n9339[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6041_6 (.CI(n39494), .I0(n18685[3]), .I1(n408_adj_4566), 
            .CO(n39495));
    SB_CARRY add_5771_7 (.CI(n39942), .I0(n14885[4]), .I1(n451), .CO(n39943));
    SB_LUT4 add_5771_6_lut (.I0(GND_net), .I1(n14885[3]), .I2(n378), .I3(n39941), 
            .O(n14164[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5981_7 (.CI(n39824), .I0(n18084[4]), .I1(n472), .CO(n39825));
    SB_LUT4 mult_10_i457_2_lut (.I0(\Kp[9] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n679_adj_4374));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i457_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i518_2_lut (.I0(\Ki[10] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n770));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i518_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i9_1_lut (.I0(PWMLimit[8]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[8]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i9_1_lut.LUT_INIT = 16'h5555;
    SB_CARRY add_5771_6 (.CI(n39941), .I0(n14885[3]), .I1(n378), .CO(n39942));
    SB_LUT4 add_4054_22_lut (.I0(GND_net), .I1(n11628[19]), .I2(GND_net), 
            .I3(n39607), .O(n9339[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5771_5_lut (.I0(GND_net), .I1(n14885[2]), .I2(n305), .I3(n39940), 
            .O(n14164[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_i179_2_lut (.I0(\Kp[3] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n265));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i179_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_6041_5_lut (.I0(GND_net), .I1(n18685[2]), .I2(n335_adj_4564), 
            .I3(n39493), .O(n18524[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5771_5 (.CI(n39940), .I0(n14885[2]), .I1(n305), .CO(n39941));
    SB_LUT4 add_5771_4_lut (.I0(GND_net), .I1(n14885[1]), .I2(n232), .I3(n39939), 
            .O(n14164[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5771_4 (.CI(n39939), .I0(n14885[1]), .I1(n232), .CO(n39940));
    SB_LUT4 add_5771_3_lut (.I0(GND_net), .I1(n14885[0]), .I2(n159), .I3(n39938), 
            .O(n14164[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5981_6_lut (.I0(GND_net), .I1(n18084[3]), .I2(n399), .I3(n39823), 
            .O(n17797[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5981_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4054_22 (.CI(n39607), .I0(n11628[19]), .I1(GND_net), 
            .CO(n39608));
    SB_LUT4 add_4054_21_lut (.I0(GND_net), .I1(n11628[18]), .I2(GND_net), 
            .I3(n39606), .O(n9339[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5771_3 (.CI(n39938), .I0(n14885[0]), .I1(n159), .CO(n39939));
    SB_CARRY add_5981_6 (.CI(n39823), .I0(n18084[3]), .I1(n399), .CO(n39824));
    SB_LUT4 mult_10_i228_2_lut (.I0(\Kp[4] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n338));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i228_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i751_2_lut (.I0(\Kp[15] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n1117));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i751_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5981_5_lut (.I0(GND_net), .I1(n18084[2]), .I2(n326), .I3(n39822), 
            .O(n17797[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5981_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5981_5 (.CI(n39822), .I0(n18084[2]), .I1(n326), .CO(n39823));
    SB_CARRY add_5969_5 (.CI(n39388), .I0(n17941[2]), .I1(n326_adj_4565), 
            .CO(n39389));
    SB_LUT4 add_5771_2_lut (.I0(GND_net), .I1(n17_adj_4563), .I2(n86), 
            .I3(GND_net), .O(n14164[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5771_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5981_4_lut (.I0(GND_net), .I1(n18084[1]), .I2(n253_adj_4561), 
            .I3(n39821), .O(n17797[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5981_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5771_2 (.CI(GND_net), .I0(n17_adj_4563), .I1(n86), .CO(n39938));
    SB_LUT4 mult_11_i104_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n153));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i104_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i298_2_lut (.I0(\Kp[6] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n442));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i298_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_4054_21 (.CI(n39606), .I0(n11628[18]), .I1(GND_net), 
            .CO(n39607));
    SB_LUT4 add_5969_4_lut (.I0(GND_net), .I1(n17941[1]), .I2(n253), .I3(n39387), 
            .O(n17629[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5969_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6041_5 (.CI(n39493), .I0(n18685[2]), .I1(n335_adj_4564), 
            .CO(n39494));
    SB_LUT4 add_4054_20_lut (.I0(GND_net), .I1(n11628[17]), .I2(GND_net), 
            .I3(n39605), .O(n9339[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5981_4 (.CI(n39821), .I0(n18084[1]), .I1(n253_adj_4561), 
            .CO(n39822));
    SB_LUT4 add_5807_19_lut (.I0(GND_net), .I1(n15532[16]), .I2(GND_net), 
            .I3(n39937), .O(n14885[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5807_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6041_4_lut (.I0(GND_net), .I1(n18685[1]), .I2(n262_adj_4560), 
            .I3(n39492), .O(n18524[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_15 (.CI(n39125), .I0(n106[13]), .I1(n155[13]), .CO(n39126));
    SB_CARRY add_4054_20 (.CI(n39605), .I0(n11628[17]), .I1(GND_net), 
            .CO(n39606));
    SB_LUT4 add_5807_18_lut (.I0(GND_net), .I1(n15532[15]), .I2(GND_net), 
            .I3(n39936), .O(n14885[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5807_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5807_18 (.CI(n39936), .I0(n15532[15]), .I1(GND_net), 
            .CO(n39937));
    SB_CARRY add_5969_4 (.CI(n39387), .I0(n17941[1]), .I1(n253), .CO(n39388));
    SB_CARRY add_6041_4 (.CI(n39492), .I0(n18685[1]), .I1(n262_adj_4560), 
            .CO(n39493));
    SB_LUT4 add_12_14_lut (.I0(GND_net), .I1(n106[12]), .I2(n155[12]), 
            .I3(n39124), .O(duty_23__N_3672[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5807_17_lut (.I0(GND_net), .I1(n15532[14]), .I2(GND_net), 
            .I3(n39935), .O(n14885[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5807_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4054_19_lut (.I0(GND_net), .I1(n11628[16]), .I2(GND_net), 
            .I3(n39604), .O(n9339[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_19_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5981_3_lut (.I0(GND_net), .I1(n18084[0]), .I2(n180_adj_4559), 
            .I3(n39820), .O(n17797[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5981_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4054_19 (.CI(n39604), .I0(n11628[16]), .I1(GND_net), 
            .CO(n39605));
    SB_LUT4 add_5969_3_lut (.I0(GND_net), .I1(n17941[0]), .I2(n180), .I3(n39386), 
            .O(n17629[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5969_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6041_3_lut (.I0(GND_net), .I1(n18685[0]), .I2(n189_adj_4558), 
            .I3(n39491), .O(n18524[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_14 (.CI(n39124), .I0(n106[12]), .I1(n155[12]), .CO(n39125));
    SB_CARRY add_6041_3 (.CI(n39491), .I0(n18685[0]), .I1(n189_adj_4558), 
            .CO(n39492));
    SB_CARRY add_5807_17 (.CI(n39935), .I0(n15532[14]), .I1(GND_net), 
            .CO(n39936));
    SB_LUT4 add_4054_18_lut (.I0(GND_net), .I1(n11628[15]), .I2(GND_net), 
            .I3(n39603), .O(n9339[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6041_2_lut (.I0(GND_net), .I1(n47_adj_4557), .I2(n116_adj_4556), 
            .I3(GND_net), .O(n18524[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6041_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5981_3 (.CI(n39820), .I0(n18084[0]), .I1(n180_adj_4559), 
            .CO(n39821));
    SB_LUT4 i35123_2_lut_4_lut (.I0(duty_23__N_3672[21]), .I1(n257[21]), 
            .I2(duty_23__N_3672[9]), .I3(n257[9]), .O(n50075));
    defparam i35123_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 i35134_2_lut_4_lut (.I0(duty_23__N_3672[16]), .I1(n257[16]), 
            .I2(duty_23__N_3672[7]), .I3(n257[7]), .O(n50086));
    defparam i35134_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_5807_16_lut (.I0(GND_net), .I1(n15532[13]), .I2(n1111), 
            .I3(n39934), .O(n14885[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5807_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4054_18 (.CI(n39603), .I0(n11628[15]), .I1(GND_net), 
            .CO(n39604));
    SB_CARRY add_5807_16 (.CI(n39934), .I0(n15532[13]), .I1(n1111), .CO(n39935));
    SB_LUT4 i35161_2_lut_4_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3672[21]), 
            .I2(PWMLimit[9]), .I3(duty_23__N_3672[9]), .O(n50113));
    defparam i35161_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_5807_15_lut (.I0(GND_net), .I1(n15532[12]), .I2(n1038), 
            .I3(n39933), .O(n14885[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5807_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6041_2 (.CI(GND_net), .I0(n47_adj_4557), .I1(n116_adj_4556), 
            .CO(n39491));
    SB_CARRY add_5969_3 (.CI(n39386), .I0(n17941[0]), .I1(n180), .CO(n39387));
    SB_LUT4 add_5981_2_lut (.I0(GND_net), .I1(n38_adj_4551), .I2(n107_adj_4549), 
            .I3(GND_net), .O(n17797[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5981_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4054_17_lut (.I0(GND_net), .I1(n11628[14]), .I2(GND_net), 
            .I3(n39602), .O(n9339[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5824_18_lut (.I0(GND_net), .I1(n15821[15]), .I2(GND_net), 
            .I3(n39490), .O(n15209[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5824_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5807_15 (.CI(n39933), .I0(n15532[12]), .I1(n1038), .CO(n39934));
    SB_LUT4 add_5969_2_lut (.I0(GND_net), .I1(n38), .I2(n107), .I3(GND_net), 
            .O(n17629[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5969_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5824_17_lut (.I0(GND_net), .I1(n15821[14]), .I2(GND_net), 
            .I3(n39489), .O(n15209[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5824_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5824_17 (.CI(n39489), .I0(n15821[14]), .I1(GND_net), 
            .CO(n39490));
    SB_CARRY add_4054_17 (.CI(n39602), .I0(n11628[14]), .I1(GND_net), 
            .CO(n39603));
    SB_LUT4 add_5824_16_lut (.I0(GND_net), .I1(n15821[13]), .I2(n1114_adj_4547), 
            .I3(n39488), .O(n15209[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5824_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5981_2 (.CI(GND_net), .I0(n38_adj_4551), .I1(n107_adj_4549), 
            .CO(n39820));
    SB_LUT4 add_12_13_lut (.I0(GND_net), .I1(n106[11]), .I2(n155[11]), 
            .I3(n39123), .O(duty_23__N_3672[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5969_2 (.CI(GND_net), .I0(n38), .I1(n107), .CO(n39386));
    SB_LUT4 add_4054_16_lut (.I0(GND_net), .I1(n11628[13]), .I2(n1099), 
            .I3(n39601), .O(n9339[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5807_14_lut (.I0(GND_net), .I1(n15532[11]), .I2(n965), 
            .I3(n39932), .O(n14885[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5807_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4054_16 (.CI(n39601), .I0(n11628[13]), .I1(n1099), .CO(n39602));
    SB_LUT4 add_6083_7_lut (.I0(GND_net), .I1(n46504), .I2(n490_adj_4525), 
            .I3(n39385), .O(n18909[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6083_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_13 (.CI(n39123), .I0(n106[11]), .I1(n155[11]), .CO(n39124));
    SB_LUT4 add_6083_6_lut (.I0(GND_net), .I1(n18980[3]), .I2(n417_adj_4513), 
            .I3(n39384), .O(n18909[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6083_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_12_lut (.I0(GND_net), .I1(n106[10]), .I2(n155[10]), 
            .I3(n39122), .O(duty_23__N_3672[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4054_15_lut (.I0(GND_net), .I1(n11628[12]), .I2(n1026), 
            .I3(n39600), .O(n9339[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4054_15 (.CI(n39600), .I0(n11628[12]), .I1(n1026), .CO(n39601));
    SB_CARRY add_12_12 (.CI(n39122), .I0(n106[10]), .I1(n155[10]), .CO(n39123));
    SB_CARRY add_5807_14 (.CI(n39932), .I0(n15532[11]), .I1(n965), .CO(n39933));
    SB_LUT4 i35171_2_lut_4_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3672[16]), 
            .I2(PWMLimit[7]), .I3(duty_23__N_3672[7]), .O(n50123));
    defparam i35171_2_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 add_5807_13_lut (.I0(GND_net), .I1(n15532[10]), .I2(n892), 
            .I3(n39931), .O(n14885[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5807_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5807_13 (.CI(n39931), .I0(n15532[10]), .I1(n892), .CO(n39932));
    SB_LUT4 add_5807_12_lut (.I0(GND_net), .I1(n15532[9]), .I2(n819), 
            .I3(n39930), .O(n14885[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5807_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_11_lut (.I0(GND_net), .I1(n106[9]), .I2(n155[9]), .I3(n39121), 
            .O(duty_23__N_3672[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5807_12 (.CI(n39930), .I0(n15532[9]), .I1(n819), .CO(n39931));
    SB_CARRY add_12_11 (.CI(n39121), .I0(n106[9]), .I1(n155[9]), .CO(n39122));
    SB_LUT4 add_5807_11_lut (.I0(GND_net), .I1(n15532[8]), .I2(n746), 
            .I3(n39929), .O(n14885[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5807_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5807_11 (.CI(n39929), .I0(n15532[8]), .I1(n746), .CO(n39930));
    SB_CARRY add_6083_6 (.CI(n39384), .I0(n18980[3]), .I1(n417_adj_4513), 
            .CO(n39385));
    SB_LUT4 add_4054_14_lut (.I0(GND_net), .I1(n11628[11]), .I2(n953), 
            .I3(n39599), .O(n9339[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4054_14 (.CI(n39599), .I0(n11628[11]), .I1(n953), .CO(n39600));
    SB_LUT4 add_4054_13_lut (.I0(GND_net), .I1(n11628[10]), .I2(n880), 
            .I3(n39598), .O(n9339[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5824_16 (.CI(n39488), .I0(n15821[13]), .I1(n1114_adj_4547), 
            .CO(n39489));
    SB_LUT4 add_5824_15_lut (.I0(GND_net), .I1(n15821[12]), .I2(n1041_adj_4509), 
            .I3(n39487), .O(n15209[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5824_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5824_15 (.CI(n39487), .I0(n15821[12]), .I1(n1041_adj_4509), 
            .CO(n39488));
    SB_LUT4 add_5824_14_lut (.I0(GND_net), .I1(n15821[11]), .I2(n968_adj_4508), 
            .I3(n39486), .O(n15209[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5824_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6083_5_lut (.I0(GND_net), .I1(n18980[2]), .I2(n344_adj_4505), 
            .I3(n39383), .O(n18909[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6083_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6083_5 (.CI(n39383), .I0(n18980[2]), .I1(n344_adj_4505), 
            .CO(n39384));
    SB_LUT4 add_12_10_lut (.I0(GND_net), .I1(n106[8]), .I2(n155[8]), .I3(n39120), 
            .O(duty_23__N_3672[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_10 (.CI(n39120), .I0(n106[8]), .I1(n155[8]), .CO(n39121));
    SB_LUT4 unary_minus_16_inv_0_i15_1_lut (.I0(PWMLimit[14]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[14]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i15_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i347_2_lut (.I0(\Kp[7] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n515));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i347_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35159_3_lut_4_lut (.I0(duty_23__N_3672[3]), .I1(n257[3]), .I2(n257[2]), 
            .I3(duty_23__N_3672[2]), .O(n50111));   // verilog/motorControl.v(38[19:35])
    defparam i35159_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 LessThan_15_i6_3_lut_3_lut (.I0(duty_23__N_3672[3]), .I1(n257[3]), 
            .I2(n257[2]), .I3(GND_net), .O(n6_adj_4670));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 i34888_3_lut_4_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3672[3]), 
            .I2(duty_23__N_3672[2]), .I3(PWMLimit[2]), .O(n49840));   // verilog/motorControl.v(36[10:25])
    defparam i34888_3_lut_4_lut.LUT_INIT = 16'h6ff6;
    SB_LUT4 duty_23__I_832_i6_3_lut_3_lut (.I0(PWMLimit[3]), .I1(duty_23__N_3672[3]), 
            .I2(duty_23__N_3672[2]), .I3(GND_net), .O(n6_adj_4671));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i6_3_lut_3_lut.LUT_INIT = 16'hd4d4;
    SB_LUT4 mult_10_i155_2_lut (.I0(\Kp[3] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n229_adj_4656));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i155_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20701_2_lut (.I0(n1[6]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[6]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20701_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 add_5807_10_lut (.I0(GND_net), .I1(n15532[7]), .I2(n673), 
            .I3(n39928), .O(n14885[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5807_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_9_lut (.I0(GND_net), .I1(n106[7]), .I2(n155[7]), .I3(n39119), 
            .O(duty_23__N_3672[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4054_13 (.CI(n39598), .I0(n11628[10]), .I1(n880), .CO(n39599));
    SB_CARRY add_5824_14 (.CI(n39486), .I0(n15821[11]), .I1(n968_adj_4508), 
            .CO(n39487));
    SB_LUT4 add_4054_12_lut (.I0(GND_net), .I1(n11628[9]), .I2(n807), 
            .I3(n39597), .O(n9339[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5824_13_lut (.I0(GND_net), .I1(n15821[10]), .I2(n895), 
            .I3(n39485), .O(n15209[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5824_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_9 (.CI(n39119), .I0(n106[7]), .I1(n155[7]), .CO(n39120));
    SB_CARRY add_4054_12 (.CI(n39597), .I0(n11628[9]), .I1(n807), .CO(n39598));
    SB_CARRY add_5807_10 (.CI(n39928), .I0(n15532[7]), .I1(n673), .CO(n39929));
    SB_CARRY add_5824_13 (.CI(n39485), .I0(n15821[10]), .I1(n895), .CO(n39486));
    SB_LUT4 add_6083_4_lut (.I0(GND_net), .I1(n18980[1]), .I2(n271_adj_4428), 
            .I3(n39382), .O(n18909[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6083_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6083_4 (.CI(n39382), .I0(n18980[1]), .I1(n271_adj_4428), 
            .CO(n39383));
    SB_LUT4 add_5824_12_lut (.I0(GND_net), .I1(n15821[9]), .I2(n822), 
            .I3(n39484), .O(n15209[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5824_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5807_9_lut (.I0(GND_net), .I1(n15532[6]), .I2(n600), .I3(n39927), 
            .O(n14885[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5807_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_6083_3_lut (.I0(GND_net), .I1(n18980[0]), .I2(n198_adj_4425), 
            .I3(n39381), .O(n18909[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6083_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5807_9 (.CI(n39927), .I0(n15532[6]), .I1(n600), .CO(n39928));
    SB_LUT4 add_5807_8_lut (.I0(GND_net), .I1(n15532[5]), .I2(n527), .I3(n39926), 
            .O(n14885[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5807_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_8_lut (.I0(GND_net), .I1(n106[6]), .I2(n155[6]), .I3(n39118), 
            .O(duty_23__N_3672[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5824_12 (.CI(n39484), .I0(n15821[9]), .I1(n822), .CO(n39485));
    SB_CARRY add_5807_8 (.CI(n39926), .I0(n15532[5]), .I1(n527), .CO(n39927));
    SB_LUT4 add_5807_7_lut (.I0(GND_net), .I1(n15532[4]), .I2(n454), .I3(n39925), 
            .O(n14885[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5807_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5807_7 (.CI(n39925), .I0(n15532[4]), .I1(n454), .CO(n39926));
    SB_LUT4 add_5807_6_lut (.I0(GND_net), .I1(n15532[3]), .I2(n381), .I3(n39924), 
            .O(n14885[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5807_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4054_11_lut (.I0(GND_net), .I1(n11628[8]), .I2(n734), 
            .I3(n39596), .O(n9339[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4054_11 (.CI(n39596), .I0(n11628[8]), .I1(n734), .CO(n39597));
    SB_LUT4 add_5824_11_lut (.I0(GND_net), .I1(n15821[8]), .I2(n749), 
            .I3(n39483), .O(n15209[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5824_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5824_11 (.CI(n39483), .I0(n15821[8]), .I1(n749), .CO(n39484));
    SB_CARRY add_5807_6 (.CI(n39924), .I0(n15532[3]), .I1(n381), .CO(n39925));
    SB_LUT4 add_5807_5_lut (.I0(GND_net), .I1(n15532[2]), .I2(n308), .I3(n39923), 
            .O(n14885[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5807_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_6083_3 (.CI(n39381), .I0(n18980[0]), .I1(n198_adj_4425), 
            .CO(n39382));
    SB_LUT4 add_6083_2_lut (.I0(GND_net), .I1(n56_adj_4421), .I2(n125_adj_4420), 
            .I3(GND_net), .O(n18909[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_6083_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4054_10_lut (.I0(GND_net), .I1(n11628[7]), .I2(n661), 
            .I3(n39595), .O(n9339[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5824_10_lut (.I0(GND_net), .I1(n15821[7]), .I2(n676), 
            .I3(n39482), .O(n15209[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5824_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5807_5 (.CI(n39923), .I0(n15532[2]), .I1(n308), .CO(n39924));
    SB_CARRY add_4054_10 (.CI(n39595), .I0(n11628[7]), .I1(n661), .CO(n39596));
    SB_CARRY add_6083_2 (.CI(GND_net), .I0(n56_adj_4421), .I1(n125_adj_4420), 
            .CO(n39381));
    SB_LUT4 add_4054_9_lut (.I0(GND_net), .I1(n11628[6]), .I2(n588), .I3(n39594), 
            .O(n9339[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5824_10 (.CI(n39482), .I0(n15821[7]), .I1(n676), .CO(n39483));
    SB_LUT4 add_5807_4_lut (.I0(GND_net), .I1(n15532[1]), .I2(n235), .I3(n39922), 
            .O(n14885[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5807_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i610_2_lut (.I0(\Ki[12] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n907_adj_4655));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i610_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_12_8 (.CI(n39118), .I0(n106[6]), .I1(n155[6]), .CO(n39119));
    SB_CARRY add_4054_9 (.CI(n39594), .I0(n11628[6]), .I1(n588), .CO(n39595));
    SB_LUT4 add_5824_9_lut (.I0(GND_net), .I1(n15821[6]), .I2(n603), .I3(n39481), 
            .O(n15209[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5824_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5807_4 (.CI(n39922), .I0(n15532[1]), .I1(n235), .CO(n39923));
    SB_LUT4 add_4054_8_lut (.I0(GND_net), .I1(n11628[5]), .I2(n515_adj_4403), 
            .I3(n39593), .O(n9339[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5807_3_lut (.I0(GND_net), .I1(n15532[0]), .I2(n162), .I3(n39921), 
            .O(n14885[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5807_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5824_9 (.CI(n39481), .I0(n15821[6]), .I1(n603), .CO(n39482));
    SB_LUT4 add_12_7_lut (.I0(GND_net), .I1(n106[5]), .I2(n155[5]), .I3(n39117), 
            .O(duty_23__N_3672[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_7 (.CI(n39117), .I0(n106[5]), .I1(n155[5]), .CO(n39118));
    SB_CARRY add_5807_3 (.CI(n39921), .I0(n15532[0]), .I1(n162), .CO(n39922));
    SB_LUT4 add_12_6_lut (.I0(GND_net), .I1(n106[4]), .I2(n155[4]), .I3(n39116), 
            .O(duty_23__N_3672[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_6 (.CI(n39116), .I0(n106[4]), .I1(n155[4]), .CO(n39117));
    SB_LUT4 add_5807_2_lut (.I0(GND_net), .I1(n20_adj_4398), .I2(n89), 
            .I3(GND_net), .O(n14885[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5807_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5807_2 (.CI(GND_net), .I0(n20_adj_4398), .I1(n89), .CO(n39921));
    SB_LUT4 add_5824_8_lut (.I0(GND_net), .I1(n15821[5]), .I2(n530), .I3(n39480), 
            .O(n15209[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5824_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_5_lut (.I0(GND_net), .I1(n106[3]), .I2(n155[3]), .I3(n39115), 
            .O(duty_23__N_3672[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5824_8 (.CI(n39480), .I0(n15821[5]), .I1(n530), .CO(n39481));
    SB_LUT4 add_5824_7_lut (.I0(GND_net), .I1(n15821[4]), .I2(n457), .I3(n39479), 
            .O(n15209[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5824_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_25_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[23]), 
            .I3(n39278), .O(n257[23])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_25_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_24_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[22]), 
            .I3(n39277), .O(n257[22])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4054_8 (.CI(n39593), .I0(n11628[5]), .I1(n515_adj_4403), 
            .CO(n39594));
    SB_CARRY unary_minus_16_add_3_24 (.CI(n39277), .I0(GND_net), .I1(n1_adj_4767[22]), 
            .CO(n39278));
    SB_CARRY add_5824_7 (.CI(n39479), .I0(n15821[4]), .I1(n457), .CO(n39480));
    SB_CARRY add_12_5 (.CI(n39115), .I0(n106[3]), .I1(n155[3]), .CO(n39116));
    SB_LUT4 add_4054_7_lut (.I0(GND_net), .I1(n11628[4]), .I2(n442_adj_4375), 
            .I3(n39592), .O(n9339[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_4_lut (.I0(GND_net), .I1(n106[2]), .I2(n155[2]), .I3(n39114), 
            .O(duty_23__N_3672[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_4 (.CI(n39114), .I0(n106[2]), .I1(n155[2]), .CO(n39115));
    SB_LUT4 add_5824_6_lut (.I0(GND_net), .I1(n15821[3]), .I2(n384), .I3(n39478), 
            .O(n15209[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5824_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4054_7 (.CI(n39592), .I0(n11628[4]), .I1(n442_adj_4375), 
            .CO(n39593));
    SB_CARRY add_5824_6 (.CI(n39478), .I0(n15821[3]), .I1(n384), .CO(n39479));
    SB_LUT4 add_4054_6_lut (.I0(GND_net), .I1(n11628[3]), .I2(n369_adj_4356), 
            .I3(n39591), .O(n9339[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5824_5_lut (.I0(GND_net), .I1(n15821[2]), .I2(n311), .I3(n39477), 
            .O(n15209[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5824_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_23_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[21]), 
            .I3(n39276), .O(n257[21])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_11_i659_2_lut (.I0(\Ki[13] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [10]), 
            .I2(GND_net), .I3(GND_net), .O(n980_adj_4654));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i659_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY add_5824_5 (.CI(n39477), .I0(n15821[2]), .I1(n311), .CO(n39478));
    SB_CARRY add_4054_6 (.CI(n39591), .I0(n11628[3]), .I1(n369_adj_4356), 
            .CO(n39592));
    SB_LUT4 add_4054_5_lut (.I0(GND_net), .I1(n11628[2]), .I2(n296_adj_4352), 
            .I3(n39590), .O(n9339[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4054_5 (.CI(n39590), .I0(n11628[2]), .I1(n296_adj_4352), 
            .CO(n39591));
    SB_LUT4 add_12_3_lut (.I0(GND_net), .I1(n106[1]), .I2(n155[1]), .I3(n39113), 
            .O(duty_23__N_3672[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4054_4_lut (.I0(GND_net), .I1(n11628[1]), .I2(n223), .I3(n39589), 
            .O(n9339[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5824_4_lut (.I0(GND_net), .I1(n15821[1]), .I2(n238), .I3(n39476), 
            .O(n15209[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5824_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_23 (.CI(n39276), .I0(GND_net), .I1(n1_adj_4767[21]), 
            .CO(n39277));
    SB_CARRY add_4054_4 (.CI(n39589), .I0(n11628[1]), .I1(n223), .CO(n39590));
    SB_LUT4 add_4054_3_lut (.I0(GND_net), .I1(n11628[0]), .I2(n150), .I3(n39588), 
            .O(n9339[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5992_12_lut (.I0(GND_net), .I1(n18205[9]), .I2(n840), 
            .I3(n39375), .O(n17941[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4054_3 (.CI(n39588), .I0(n11628[0]), .I1(n150), .CO(n39589));
    SB_LUT4 add_4054_2_lut (.I0(GND_net), .I1(n8_adj_4351), .I2(n77), 
            .I3(GND_net), .O(n9339[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4054_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4054_2 (.CI(GND_net), .I0(n8_adj_4351), .I1(n77), .CO(n39588));
    SB_LUT4 add_5299_22_lut (.I0(GND_net), .I1(n12924[19]), .I2(GND_net), 
            .I3(n39587), .O(n11628[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5299_21_lut (.I0(GND_net), .I1(n12924[18]), .I2(GND_net), 
            .I3(n39586), .O(n11628[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_21_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_22_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[20]), 
            .I3(n39275), .O(n257[20])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5824_4 (.CI(n39476), .I0(n15821[1]), .I1(n238), .CO(n39477));
    SB_CARRY add_5299_21 (.CI(n39586), .I0(n12924[18]), .I1(GND_net), 
            .CO(n39587));
    SB_LUT4 add_5299_20_lut (.I0(GND_net), .I1(n12924[17]), .I2(GND_net), 
            .I3(n39585), .O(n11628[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_20_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5824_3_lut (.I0(GND_net), .I1(n15821[0]), .I2(n165), .I3(n39475), 
            .O(n15209[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5824_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5299_20 (.CI(n39585), .I0(n12924[17]), .I1(GND_net), 
            .CO(n39586));
    SB_LUT4 add_5992_11_lut (.I0(GND_net), .I1(n18205[8]), .I2(n767), 
            .I3(n39374), .O(n17941[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5824_3 (.CI(n39475), .I0(n15821[0]), .I1(n165), .CO(n39476));
    SB_LUT4 add_5824_2_lut (.I0(GND_net), .I1(n23_adj_4348), .I2(n92), 
            .I3(GND_net), .O(n15209[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5824_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5299_19_lut (.I0(GND_net), .I1(n12924[16]), .I2(GND_net), 
            .I3(n39584), .O(n11628[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_3 (.CI(n39113), .I0(n106[1]), .I1(n155[1]), .CO(n39114));
    SB_CARRY add_5299_19 (.CI(n39584), .I0(n12924[16]), .I1(GND_net), 
            .CO(n39585));
    SB_CARRY add_5824_2 (.CI(GND_net), .I0(n23_adj_4348), .I1(n92), .CO(n39475));
    SB_LUT4 add_5299_18_lut (.I0(GND_net), .I1(n12924[15]), .I2(GND_net), 
            .I3(n39583), .O(n11628[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5299_18 (.CI(n39583), .I0(n12924[15]), .I1(GND_net), 
            .CO(n39584));
    SB_LUT4 add_5857_17_lut (.I0(GND_net), .I1(n16365[14]), .I2(GND_net), 
            .I3(n39474), .O(n15821[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5857_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5857_16_lut (.I0(GND_net), .I1(n16365[13]), .I2(n1117_adj_4347), 
            .I3(n39473), .O(n15821[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5857_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5857_16 (.CI(n39473), .I0(n16365[13]), .I1(n1117_adj_4347), 
            .CO(n39474));
    SB_LUT4 add_5299_17_lut (.I0(GND_net), .I1(n12924[14]), .I2(GND_net), 
            .I3(n39582), .O(n11628[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5299_17 (.CI(n39582), .I0(n12924[14]), .I1(GND_net), 
            .CO(n39583));
    SB_LUT4 add_5299_16_lut (.I0(GND_net), .I1(n12924[13]), .I2(n1102), 
            .I3(n39581), .O(n11628[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5299_16 (.CI(n39581), .I0(n12924[13]), .I1(n1102), .CO(n39582));
    SB_LUT4 add_5857_15_lut (.I0(GND_net), .I1(n16365[12]), .I2(n1044), 
            .I3(n39472), .O(n15821[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5857_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5992_11 (.CI(n39374), .I0(n18205[8]), .I1(n767), .CO(n39375));
    SB_LUT4 add_5299_15_lut (.I0(GND_net), .I1(n12924[12]), .I2(n1029), 
            .I3(n39580), .O(n11628[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_24_lut (.I0(n1[23]), .I1(n9870[21]), .I2(GND_net), 
            .I3(n40037), .O(n9363[0])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_24_lut.LUT_INIT = 16'h6996;
    SB_LUT4 mult_10_add_1225_23_lut (.I0(GND_net), .I1(n9870[20]), .I2(GND_net), 
            .I3(n40036), .O(n106[22])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5857_15 (.CI(n39472), .I0(n16365[12]), .I1(n1044), .CO(n39473));
    SB_CARRY mult_10_add_1225_23 (.CI(n40036), .I0(n9870[20]), .I1(GND_net), 
            .CO(n40037));
    SB_LUT4 add_5992_10_lut (.I0(GND_net), .I1(n18205[7]), .I2(n694), 
            .I3(n39373), .O(n17941[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_22_lut (.I0(GND_net), .I1(n9870[19]), .I2(GND_net), 
            .I3(n40035), .O(n106[21])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_22_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5857_14_lut (.I0(GND_net), .I1(n16365[11]), .I2(n971_adj_4346), 
            .I3(n39471), .O(n15821[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5857_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_22 (.CI(n40035), .I0(n9870[19]), .I1(GND_net), 
            .CO(n40036));
    SB_LUT4 mult_10_add_1225_21_lut (.I0(GND_net), .I1(n9870[18]), .I2(GND_net), 
            .I3(n40034), .O(n106[20])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5857_14 (.CI(n39471), .I0(n16365[11]), .I1(n971_adj_4346), 
            .CO(n39472));
    SB_CARRY mult_10_add_1225_21 (.CI(n40034), .I0(n9870[18]), .I1(GND_net), 
            .CO(n40035));
    SB_LUT4 mult_10_add_1225_20_lut (.I0(GND_net), .I1(n9870[17]), .I2(GND_net), 
            .I3(n40033), .O(n106[19])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5299_15 (.CI(n39580), .I0(n12924[12]), .I1(n1029), .CO(n39581));
    SB_CARRY mult_10_add_1225_20 (.CI(n40033), .I0(n9870[17]), .I1(GND_net), 
            .CO(n40034));
    SB_LUT4 mult_10_add_1225_19_lut (.I0(GND_net), .I1(n9870[16]), .I2(GND_net), 
            .I3(n40032), .O(n106[18])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_19 (.CI(n40032), .I0(n9870[16]), .I1(GND_net), 
            .CO(n40033));
    SB_LUT4 mult_10_add_1225_18_lut (.I0(GND_net), .I1(n9870[15]), .I2(GND_net), 
            .I3(n40031), .O(n106[17])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_18_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5857_13_lut (.I0(GND_net), .I1(n16365[10]), .I2(n898), 
            .I3(n39470), .O(n15821[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5857_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_18 (.CI(n40031), .I0(n9870[15]), .I1(GND_net), 
            .CO(n40032));
    SB_LUT4 mult_10_add_1225_17_lut (.I0(GND_net), .I1(n9870[14]), .I2(GND_net), 
            .I3(n40030), .O(n106[16])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_17 (.CI(n40030), .I0(n9870[14]), .I1(GND_net), 
            .CO(n40031));
    SB_LUT4 mult_10_add_1225_16_lut (.I0(GND_net), .I1(n9870[13]), .I2(n1096), 
            .I3(n40029), .O(n106[15])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_16 (.CI(n40029), .I0(n9870[13]), .I1(n1096), 
            .CO(n40030));
    SB_CARRY add_5992_10 (.CI(n39373), .I0(n18205[7]), .I1(n694), .CO(n39374));
    SB_LUT4 mult_10_add_1225_15_lut (.I0(GND_net), .I1(n9870[12]), .I2(n1023), 
            .I3(n40028), .O(n106[14])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5992_9_lut (.I0(GND_net), .I1(n18205[6]), .I2(n621), .I3(n39372), 
            .O(n17941[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_15 (.CI(n40028), .I0(n9870[12]), .I1(n1023), 
            .CO(n40029));
    SB_LUT4 mult_10_add_1225_14_lut (.I0(GND_net), .I1(n9870[11]), .I2(n950), 
            .I3(n40027), .O(n106[13])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5857_13 (.CI(n39470), .I0(n16365[10]), .I1(n898), .CO(n39471));
    SB_CARRY add_5992_9 (.CI(n39372), .I0(n18205[6]), .I1(n621), .CO(n39373));
    SB_LUT4 add_5299_14_lut (.I0(GND_net), .I1(n12924[11]), .I2(n956), 
            .I3(n39579), .O(n11628[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5992_8_lut (.I0(GND_net), .I1(n18205[5]), .I2(n548), .I3(n39371), 
            .O(n17941[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_14 (.CI(n40027), .I0(n9870[11]), .I1(n950), 
            .CO(n40028));
    SB_CARRY unary_minus_16_add_3_22 (.CI(n39275), .I0(GND_net), .I1(n1_adj_4767[20]), 
            .CO(n39276));
    SB_CARRY add_5299_14 (.CI(n39579), .I0(n12924[11]), .I1(n956), .CO(n39580));
    SB_LUT4 mult_10_add_1225_13_lut (.I0(GND_net), .I1(n9870[10]), .I2(n877), 
            .I3(n40026), .O(n106[12])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5299_13_lut (.I0(GND_net), .I1(n12924[10]), .I2(n883), 
            .I3(n39578), .O(n11628[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5992_8 (.CI(n39371), .I0(n18205[5]), .I1(n548), .CO(n39372));
    SB_LUT4 add_5992_7_lut (.I0(GND_net), .I1(n18205[4]), .I2(n475), .I3(n39370), 
            .O(n17941[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_21_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[19]), 
            .I3(n39274), .O(n257[19])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_13 (.CI(n40026), .I0(n9870[10]), .I1(n877), 
            .CO(n40027));
    SB_LUT4 mult_10_add_1225_12_lut (.I0(GND_net), .I1(n9870[9]), .I2(n804), 
            .I3(n40025), .O(n106[11])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5992_7 (.CI(n39370), .I0(n18205[4]), .I1(n475), .CO(n39371));
    SB_LUT4 add_12_2_lut (.I0(GND_net), .I1(n106[0]), .I2(n155[0]), .I3(GND_net), 
            .O(duty_23__N_3672[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_21 (.CI(n39274), .I0(GND_net), .I1(n1_adj_4767[19]), 
            .CO(n39275));
    SB_CARRY mult_10_add_1225_12 (.CI(n40025), .I0(n9870[9]), .I1(n804), 
            .CO(n40026));
    SB_LUT4 add_5857_12_lut (.I0(GND_net), .I1(n16365[9]), .I2(n825), 
            .I3(n39469), .O(n15821[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5857_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5992_6_lut (.I0(GND_net), .I1(n18205[3]), .I2(n402), .I3(n39369), 
            .O(n17941[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5992_6 (.CI(n39369), .I0(n18205[3]), .I1(n402), .CO(n39370));
    SB_LUT4 add_5992_5_lut (.I0(GND_net), .I1(n18205[2]), .I2(n329), .I3(n39368), 
            .O(n17941[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5299_13 (.CI(n39578), .I0(n12924[10]), .I1(n883), .CO(n39579));
    SB_CARRY add_5857_12 (.CI(n39469), .I0(n16365[9]), .I1(n825), .CO(n39470));
    SB_LUT4 unary_minus_16_add_3_20_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[18]), 
            .I3(n39273), .O(n257[18])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_20 (.CI(n39273), .I0(GND_net), .I1(n1_adj_4767[18]), 
            .CO(n39274));
    SB_CARRY add_12_2 (.CI(GND_net), .I0(n106[0]), .I1(n155[0]), .CO(n39113));
    SB_LUT4 mult_10_add_1225_11_lut (.I0(GND_net), .I1(n9870[8]), .I2(n731), 
            .I3(n40024), .O(n106[10])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_11 (.CI(n40024), .I0(n9870[8]), .I1(n731), 
            .CO(n40025));
    SB_LUT4 add_5299_12_lut (.I0(GND_net), .I1(n12924[9]), .I2(n810), 
            .I3(n39577), .O(n11628[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_12_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_10_lut (.I0(GND_net), .I1(n9870[7]), .I2(n658), 
            .I3(n40023), .O(n106[9])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_10 (.CI(n40023), .I0(n9870[7]), .I1(n658), 
            .CO(n40024));
    SB_CARRY add_5992_5 (.CI(n39368), .I0(n18205[2]), .I1(n329), .CO(n39369));
    SB_LUT4 mult_10_add_1225_9_lut (.I0(GND_net), .I1(n9870[6]), .I2(n585), 
            .I3(n40022), .O(n106[8])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5841_18_lut (.I0(GND_net), .I1(n16109[15]), .I2(GND_net), 
            .I3(n39900), .O(n15532[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_9 (.CI(n40022), .I0(n9870[6]), .I1(n585), 
            .CO(n40023));
    SB_LUT4 add_5841_17_lut (.I0(GND_net), .I1(n16109[14]), .I2(GND_net), 
            .I3(n39899), .O(n15532[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_8_lut (.I0(GND_net), .I1(n9870[5]), .I2(n512), 
            .I3(n40021), .O(n106[7])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5299_12 (.CI(n39577), .I0(n12924[9]), .I1(n810), .CO(n39578));
    SB_CARRY add_5841_17 (.CI(n39899), .I0(n16109[14]), .I1(GND_net), 
            .CO(n39900));
    SB_CARRY mult_10_add_1225_8 (.CI(n40021), .I0(n9870[5]), .I1(n512), 
            .CO(n40022));
    SB_LUT4 mult_10_add_1225_7_lut (.I0(GND_net), .I1(n9870[4]), .I2(n439), 
            .I3(n40020), .O(n106[6])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5299_11_lut (.I0(GND_net), .I1(n12924[8]), .I2(n737), 
            .I3(n39576), .O(n11628[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5857_11_lut (.I0(GND_net), .I1(n16365[8]), .I2(n752), 
            .I3(n39468), .O(n15821[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5857_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5841_16_lut (.I0(GND_net), .I1(n16109[13]), .I2(n1114), 
            .I3(n39898), .O(n15532[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5992_4_lut (.I0(GND_net), .I1(n18205[1]), .I2(n256), .I3(n39367), 
            .O(n17941[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_7 (.CI(n40020), .I0(n9870[4]), .I1(n439), 
            .CO(n40021));
    SB_CARRY add_5841_16 (.CI(n39898), .I0(n16109[13]), .I1(n1114), .CO(n39899));
    SB_CARRY add_5299_11 (.CI(n39576), .I0(n12924[8]), .I1(n737), .CO(n39577));
    SB_LUT4 unary_minus_16_add_3_19_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[17]), 
            .I3(n39272), .O(n257[17])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5857_11 (.CI(n39468), .I0(n16365[8]), .I1(n752), .CO(n39469));
    SB_CARRY unary_minus_16_add_3_19 (.CI(n39272), .I0(GND_net), .I1(n1_adj_4767[17]), 
            .CO(n39273));
    SB_LUT4 mult_10_add_1225_6_lut (.I0(GND_net), .I1(n9870[3]), .I2(n366), 
            .I3(n40019), .O(n106[5])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5299_10_lut (.I0(GND_net), .I1(n12924[7]), .I2(n664), 
            .I3(n39575), .O(n11628[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5857_10_lut (.I0(GND_net), .I1(n16365[7]), .I2(n679), 
            .I3(n39467), .O(n15821[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5857_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_6 (.CI(n40019), .I0(n9870[3]), .I1(n366), 
            .CO(n40020));
    SB_LUT4 add_5841_15_lut (.I0(GND_net), .I1(n16109[12]), .I2(n1041), 
            .I3(n39897), .O(n15532[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_15_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_5_lut (.I0(GND_net), .I1(n9870[2]), .I2(n293), 
            .I3(n40018), .O(n106[4])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_15 (.CI(n39897), .I0(n16109[12]), .I1(n1041), .CO(n39898));
    SB_CARRY add_5299_10 (.CI(n39575), .I0(n12924[7]), .I1(n664), .CO(n39576));
    SB_LUT4 add_5841_14_lut (.I0(GND_net), .I1(n16109[11]), .I2(n968), 
            .I3(n39896), .O(n15532[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_14 (.CI(n39896), .I0(n16109[11]), .I1(n968), .CO(n39897));
    SB_CARRY mult_10_add_1225_5 (.CI(n40018), .I0(n9870[2]), .I1(n293), 
            .CO(n40019));
    SB_CARRY add_5992_4 (.CI(n39367), .I0(n18205[1]), .I1(n256), .CO(n39368));
    SB_LUT4 add_5299_9_lut (.I0(GND_net), .I1(n12924[6]), .I2(n591), .I3(n39574), 
            .O(n11628[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_4_lut (.I0(GND_net), .I1(n9870[1]), .I2(n220), 
            .I3(n40017), .O(n106[3])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_4 (.CI(n40017), .I0(n9870[1]), .I1(n220), 
            .CO(n40018));
    SB_LUT4 add_5841_13_lut (.I0(GND_net), .I1(n16109[10]), .I2(n895_adj_4675), 
            .I3(n39895), .O(n15532[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mult_10_add_1225_3_lut (.I0(GND_net), .I1(n9870[0]), .I2(n147_adj_4676), 
            .I3(n40016), .O(n106[2])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY mult_10_add_1225_3 (.CI(n40016), .I0(n9870[0]), .I1(n147_adj_4676), 
            .CO(n40017));
    SB_CARRY add_5841_13 (.CI(n39895), .I0(n16109[10]), .I1(n895_adj_4675), 
            .CO(n39896));
    SB_LUT4 mult_10_add_1225_2_lut (.I0(GND_net), .I1(n5_adj_4677), .I2(n74_adj_4678), 
            .I3(GND_net), .O(n106[1])) /* synthesis syn_instantiated=1 */ ;
    defparam mult_10_add_1225_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5841_12_lut (.I0(GND_net), .I1(n16109[9]), .I2(n822_adj_4679), 
            .I3(n39894), .O(n15532[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_12 (.CI(n39894), .I0(n16109[9]), .I1(n822_adj_4679), 
            .CO(n39895));
    SB_CARRY add_5299_9 (.CI(n39574), .I0(n12924[6]), .I1(n591), .CO(n39575));
    SB_LUT4 add_5841_11_lut (.I0(GND_net), .I1(n16109[8]), .I2(n749_adj_4680), 
            .I3(n39893), .O(n15532[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5299_8_lut (.I0(GND_net), .I1(n12924[5]), .I2(n518_adj_4681), 
            .I3(n39573), .O(n11628[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5992_3_lut (.I0(GND_net), .I1(n18205[0]), .I2(n183_adj_4682), 
            .I3(n39366), .O(n17941[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 unary_minus_16_add_3_18_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[16]), 
            .I3(n39271), .O(n257[16])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5857_10 (.CI(n39467), .I0(n16365[7]), .I1(n679), .CO(n39468));
    SB_LUT4 add_5857_9_lut (.I0(GND_net), .I1(n16365[6]), .I2(n606_adj_4684), 
            .I3(n39466), .O(n15821[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5857_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5299_8 (.CI(n39573), .I0(n12924[5]), .I1(n518_adj_4681), 
            .CO(n39574));
    SB_CARRY add_5841_11 (.CI(n39893), .I0(n16109[8]), .I1(n749_adj_4680), 
            .CO(n39894));
    SB_CARRY mult_10_add_1225_2 (.CI(GND_net), .I0(n5_adj_4677), .I1(n74_adj_4678), 
            .CO(n40016));
    SB_LUT4 add_5841_10_lut (.I0(GND_net), .I1(n16109[7]), .I2(n676_adj_4685), 
            .I3(n39892), .O(n15532[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_10 (.CI(n39892), .I0(n16109[7]), .I1(n676_adj_4685), 
            .CO(n39893));
    SB_LUT4 add_4077_23_lut (.I0(GND_net), .I1(n12113[20]), .I2(GND_net), 
            .I3(n40015), .O(n9870[21])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_23_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5841_9_lut (.I0(GND_net), .I1(n16109[6]), .I2(n603_adj_4686), 
            .I3(n39891), .O(n15532[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5857_9 (.CI(n39466), .I0(n16365[6]), .I1(n606_adj_4684), 
            .CO(n39467));
    SB_LUT4 add_5857_8_lut (.I0(GND_net), .I1(n16365[5]), .I2(n533_adj_4687), 
            .I3(n39465), .O(n15821[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5857_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_18 (.CI(n39271), .I0(GND_net), .I1(n1_adj_4767[16]), 
            .CO(n39272));
    SB_LUT4 add_5299_7_lut (.I0(GND_net), .I1(n12924[4]), .I2(n445_adj_4688), 
            .I3(n39572), .O(n11628[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_9 (.CI(n39891), .I0(n16109[6]), .I1(n603_adj_4686), 
            .CO(n39892));
    SB_LUT4 unary_minus_16_add_3_17_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[15]), 
            .I3(n39270), .O(n257[15])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5992_3 (.CI(n39366), .I0(n18205[0]), .I1(n183_adj_4682), 
            .CO(n39367));
    SB_LUT4 add_5841_8_lut (.I0(GND_net), .I1(n16109[5]), .I2(n530_adj_4690), 
            .I3(n39890), .O(n15532[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5857_8 (.CI(n39465), .I0(n16365[5]), .I1(n533_adj_4687), 
            .CO(n39466));
    SB_LUT4 add_5857_7_lut (.I0(GND_net), .I1(n16365[4]), .I2(n460_adj_4691), 
            .I3(n39464), .O(n15821[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5857_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5992_2_lut (.I0(GND_net), .I1(n41_adj_4692), .I2(n110_adj_4693), 
            .I3(GND_net), .O(n17941[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5992_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5299_7 (.CI(n39572), .I0(n12924[4]), .I1(n445_adj_4688), 
            .CO(n39573));
    SB_LUT4 add_4077_22_lut (.I0(GND_net), .I1(n12113[19]), .I2(GND_net), 
            .I3(n40014), .O(n9870[20])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY unary_minus_16_add_3_17 (.CI(n39270), .I0(GND_net), .I1(n1_adj_4767[15]), 
            .CO(n39271));
    SB_CARRY add_5992_2 (.CI(GND_net), .I0(n41_adj_4692), .I1(n110_adj_4693), 
            .CO(n39366));
    SB_CARRY add_5841_8 (.CI(n39890), .I0(n16109[5]), .I1(n530_adj_4690), 
            .CO(n39891));
    SB_CARRY add_5857_7 (.CI(n39464), .I0(n16365[4]), .I1(n460_adj_4691), 
            .CO(n39465));
    SB_LUT4 add_5841_7_lut (.I0(GND_net), .I1(n16109[4]), .I2(n457_adj_4694), 
            .I3(n39889), .O(n15532[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4077_22 (.CI(n40014), .I0(n12113[19]), .I1(GND_net), 
            .CO(n40015));
    SB_LUT4 add_5299_6_lut (.I0(GND_net), .I1(n12924[3]), .I2(n372_adj_4695), 
            .I3(n39571), .O(n11628[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_7 (.CI(n39889), .I0(n16109[4]), .I1(n457_adj_4694), 
            .CO(n39890));
    SB_CARRY add_5299_6 (.CI(n39571), .I0(n12924[3]), .I1(n372_adj_4695), 
            .CO(n39572));
    SB_LUT4 add_5841_6_lut (.I0(GND_net), .I1(n16109[3]), .I2(n384_adj_4696), 
            .I3(n39888), .O(n15532[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_6 (.CI(n39888), .I0(n16109[3]), .I1(n384_adj_4696), 
            .CO(n39889));
    SB_LUT4 add_4077_21_lut (.I0(GND_net), .I1(n12113[18]), .I2(GND_net), 
            .I3(n40013), .O(n9870[19])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4077_21 (.CI(n40013), .I0(n12113[18]), .I1(GND_net), 
            .CO(n40014));
    SB_LUT4 add_5841_5_lut (.I0(GND_net), .I1(n16109[2]), .I2(n311_adj_4697), 
            .I3(n39887), .O(n15532[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_5 (.CI(n39887), .I0(n16109[2]), .I1(n311_adj_4697), 
            .CO(n39888));
    SB_LUT4 add_5299_5_lut (.I0(GND_net), .I1(n12924[2]), .I2(n299_adj_4698), 
            .I3(n39570), .O(n11628[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5299_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5841_4_lut (.I0(GND_net), .I1(n16109[1]), .I2(n238_adj_4699), 
            .I3(n39886), .O(n15532[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5857_6_lut (.I0(GND_net), .I1(n16365[3]), .I2(n387_adj_4700), 
            .I3(n39463), .O(n15821[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5857_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4077_20_lut (.I0(GND_net), .I1(n12113[17]), .I2(GND_net), 
            .I3(n40012), .O(n9870[18])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4077_20 (.CI(n40012), .I0(n12113[17]), .I1(GND_net), 
            .CO(n40013));
    SB_LUT4 add_4077_19_lut (.I0(GND_net), .I1(n12113[16]), .I2(GND_net), 
            .I3(n40011), .O(n9870[17])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4077_19 (.CI(n40011), .I0(n12113[16]), .I1(GND_net), 
            .CO(n40012));
    SB_LUT4 add_4077_18_lut (.I0(GND_net), .I1(n12113[15]), .I2(GND_net), 
            .I3(n40010), .O(n9870[16])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4077_18 (.CI(n40010), .I0(n12113[15]), .I1(GND_net), 
            .CO(n40011));
    SB_LUT4 add_4077_17_lut (.I0(GND_net), .I1(n12113[14]), .I2(GND_net), 
            .I3(n40009), .O(n9870[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4077_17 (.CI(n40009), .I0(n12113[14]), .I1(GND_net), 
            .CO(n40010));
    SB_CARRY add_5857_6 (.CI(n39463), .I0(n16365[3]), .I1(n387_adj_4700), 
            .CO(n39464));
    SB_LUT4 add_4077_16_lut (.I0(GND_net), .I1(n12113[13]), .I2(n1099_adj_4701), 
            .I3(n40008), .O(n9870[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_4 (.CI(n39886), .I0(n16109[1]), .I1(n238_adj_4699), 
            .CO(n39887));
    SB_LUT4 add_5841_3_lut (.I0(GND_net), .I1(n16109[0]), .I2(n165_adj_4702), 
            .I3(n39885), .O(n15532[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4077_16 (.CI(n40008), .I0(n12113[13]), .I1(n1099_adj_4701), 
            .CO(n40009));
    SB_LUT4 unary_minus_16_add_3_16_lut (.I0(GND_net), .I1(GND_net), .I2(n1_adj_4767[14]), 
            .I3(n39269), .O(n257[14])) /* synthesis syn_instantiated=1 */ ;
    defparam unary_minus_16_add_3_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_4077_15_lut (.I0(GND_net), .I1(n12113[12]), .I2(n1026_adj_4703), 
            .I3(n40007), .O(n9870[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_3 (.CI(n39885), .I0(n16109[0]), .I1(n165_adj_4702), 
            .CO(n39886));
    SB_CARRY add_4077_15 (.CI(n40007), .I0(n12113[12]), .I1(n1026_adj_4703), 
            .CO(n40008));
    SB_LUT4 add_4077_14_lut (.I0(GND_net), .I1(n12113[11]), .I2(n953_adj_4704), 
            .I3(n40006), .O(n9870[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4077_14 (.CI(n40006), .I0(n12113[11]), .I1(n953_adj_4704), 
            .CO(n40007));
    SB_LUT4 add_4077_13_lut (.I0(GND_net), .I1(n12113[10]), .I2(n880_adj_4705), 
            .I3(n40005), .O(n9870[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4077_13 (.CI(n40005), .I0(n12113[10]), .I1(n880_adj_4705), 
            .CO(n40006));
    SB_LUT4 add_4077_12_lut (.I0(GND_net), .I1(n12113[9]), .I2(n807_adj_4706), 
            .I3(n40004), .O(n9870[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4077_12 (.CI(n40004), .I0(n12113[9]), .I1(n807_adj_4706), 
            .CO(n40005));
    SB_LUT4 add_5841_2_lut (.I0(GND_net), .I1(n23_adj_4707), .I2(n92_adj_4708), 
            .I3(GND_net), .O(n15532[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5841_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5299_5 (.CI(n39570), .I0(n12924[2]), .I1(n299_adj_4698), 
            .CO(n39571));
    SB_LUT4 add_4077_11_lut (.I0(GND_net), .I1(n12113[8]), .I2(n734_adj_4709), 
            .I3(n40003), .O(n9870[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5857_5_lut (.I0(GND_net), .I1(n16365[2]), .I2(n314_adj_4710), 
            .I3(n39462), .O(n15821[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5857_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_5841_2 (.CI(GND_net), .I0(n23_adj_4707), .I1(n92_adj_4708), 
            .CO(n39885));
    SB_CARRY add_4077_11 (.CI(n40003), .I0(n12113[8]), .I1(n734_adj_4709), 
            .CO(n40004));
    SB_LUT4 add_4077_10_lut (.I0(GND_net), .I1(n12113[7]), .I2(n661_adj_4711), 
            .I3(n40002), .O(n9870[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5873_17_lut (.I0(GND_net), .I1(n16620[14]), .I2(GND_net), 
            .I3(n39884), .O(n16109[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5873_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4077_10 (.CI(n40002), .I0(n12113[7]), .I1(n661_adj_4711), 
            .CO(n40003));
    SB_LUT4 add_4077_9_lut (.I0(GND_net), .I1(n12113[6]), .I2(n588_adj_4712), 
            .I3(n40001), .O(n9870[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_5873_16_lut (.I0(GND_net), .I1(n16620[13]), .I2(n1117), 
            .I3(n39883), .O(n16109[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_5873_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_4077_9 (.CI(n40001), .I0(n12113[6]), .I1(n588_adj_4712), 
            .CO(n40002));
    SB_CARRY add_5857_5 (.CI(n39462), .I0(n16365[2]), .I1(n314_adj_4710), 
            .CO(n39463));
    SB_LUT4 add_4077_8_lut (.I0(GND_net), .I1(n12113[5]), .I2(n515), .I3(n40000), 
            .O(n9870[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_4077_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 duty_23__I_832_i39_2_lut (.I0(PWMLimit[19]), .I1(duty_23__N_3672[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4713));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i41_2_lut (.I0(PWMLimit[20]), .I1(duty_23__N_3672[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4714));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i45_2_lut (.I0(PWMLimit[22]), .I1(duty_23__N_3672[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4715));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i37_2_lut (.I0(PWMLimit[18]), .I1(duty_23__N_3672[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4716));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i29_2_lut (.I0(PWMLimit[14]), .I1(duty_23__N_3672[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4717));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i31_2_lut (.I0(PWMLimit[15]), .I1(duty_23__N_3672[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4718));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i43_2_lut (.I0(PWMLimit[21]), .I1(duty_23__N_3672[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4719));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i35_2_lut (.I0(PWMLimit[17]), .I1(duty_23__N_3672[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4720));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i23_2_lut (.I0(PWMLimit[11]), .I1(duty_23__N_3672[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4721));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i25_2_lut (.I0(PWMLimit[12]), .I1(duty_23__N_3672[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4722));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i33_2_lut (.I0(PWMLimit[16]), .I1(duty_23__N_3672[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4723));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i9_2_lut (.I0(PWMLimit[4]), .I1(duty_23__N_3672[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4724));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i17_2_lut (.I0(PWMLimit[8]), .I1(duty_23__N_3672[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4725));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i19_2_lut (.I0(PWMLimit[9]), .I1(duty_23__N_3672[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4726));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i21_2_lut (.I0(PWMLimit[10]), .I1(duty_23__N_3672[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4727));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i11_2_lut (.I0(PWMLimit[5]), .I1(duty_23__N_3672[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4728));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i13_2_lut (.I0(PWMLimit[6]), .I1(duty_23__N_3672[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4729));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i15_2_lut (.I0(PWMLimit[7]), .I1(duty_23__N_3672[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4730));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 duty_23__I_832_i27_2_lut (.I0(PWMLimit[13]), .I1(duty_23__N_3672[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4731));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i34878_4_lut (.I0(n21_adj_4727), .I1(n19_adj_4726), .I2(n17_adj_4725), 
            .I3(n9_adj_4724), .O(n49830));
    defparam i34878_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i34871_4_lut (.I0(n27_adj_4731), .I1(n15_adj_4730), .I2(n13_adj_4729), 
            .I3(n11_adj_4728), .O(n49823));
    defparam i34871_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 duty_23__I_832_i12_3_lut (.I0(duty_23__N_3672[7]), .I1(duty_23__N_3672[16]), 
            .I2(n33_adj_4723), .I3(GND_net), .O(n12_adj_4732));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_832_i10_3_lut (.I0(duty_23__N_3672[5]), .I1(duty_23__N_3672[6]), 
            .I2(n13_adj_4729), .I3(GND_net), .O(n10_adj_4733));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_832_i30_3_lut (.I0(n12_adj_4732), .I1(duty_23__N_3672[17]), 
            .I2(n35_adj_4720), .I3(GND_net), .O(n30_adj_4734));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35196_4_lut (.I0(n13_adj_4729), .I1(n11_adj_4728), .I2(n9_adj_4724), 
            .I3(n49840), .O(n50148));
    defparam i35196_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35192_4_lut (.I0(n19_adj_4726), .I1(n17_adj_4725), .I2(n15_adj_4730), 
            .I3(n50148), .O(n50144));
    defparam i35192_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35576_4_lut (.I0(n25_adj_4722), .I1(n23_adj_4721), .I2(n21_adj_4727), 
            .I3(n50144), .O(n50529));
    defparam i35576_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35404_4_lut (.I0(n31_adj_4718), .I1(n29_adj_4717), .I2(n27_adj_4731), 
            .I3(n50529), .O(n50357));
    defparam i35404_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35650_4_lut (.I0(n37_adj_4716), .I1(n35_adj_4720), .I2(n33_adj_4723), 
            .I3(n50357), .O(n50603));
    defparam i35650_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 duty_23__I_832_i16_3_lut (.I0(duty_23__N_3672[9]), .I1(duty_23__N_3672[21]), 
            .I2(n43_adj_4719), .I3(GND_net), .O(n16_adj_4735));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35586_3_lut (.I0(n6_adj_4671), .I1(duty_23__N_3672[10]), .I2(n21_adj_4727), 
            .I3(GND_net), .O(n50539));   // verilog/motorControl.v(36[10:25])
    defparam i35586_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35587_3_lut (.I0(n50539), .I1(duty_23__N_3672[11]), .I2(n23_adj_4721), 
            .I3(GND_net), .O(n50540));   // verilog/motorControl.v(36[10:25])
    defparam i35587_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_832_i8_3_lut (.I0(duty_23__N_3672[4]), .I1(duty_23__N_3672[8]), 
            .I2(n17_adj_4725), .I3(GND_net), .O(n8_adj_4736));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_832_i24_3_lut (.I0(n16_adj_4735), .I1(duty_23__N_3672[22]), 
            .I2(n45_adj_4715), .I3(GND_net), .O(n24_adj_4737));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35163_4_lut (.I0(n43_adj_4719), .I1(n25_adj_4722), .I2(n23_adj_4721), 
            .I3(n49830), .O(n50115));
    defparam i35163_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35534_4_lut (.I0(n24_adj_4737), .I1(n8_adj_4736), .I2(n45_adj_4715), 
            .I3(n50113), .O(n50487));   // verilog/motorControl.v(36[10:25])
    defparam i35534_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35533_3_lut (.I0(n50540), .I1(duty_23__N_3672[12]), .I2(n25_adj_4722), 
            .I3(GND_net), .O(n50486));   // verilog/motorControl.v(36[10:25])
    defparam i35533_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_832_i4_4_lut (.I0(duty_23__N_3672[0]), .I1(duty_23__N_3672[1]), 
            .I2(PWMLimit[1]), .I3(PWMLimit[0]), .O(n4_adj_4738));   // verilog/motorControl.v(36[10:25])
    defparam duty_23__I_832_i4_4_lut.LUT_INIT = 16'h0c8e;
    SB_LUT4 i35548_3_lut (.I0(n4_adj_4738), .I1(duty_23__N_3672[13]), .I2(n27_adj_4731), 
            .I3(GND_net), .O(n50501));   // verilog/motorControl.v(36[10:25])
    defparam i35548_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35549_3_lut (.I0(n50501), .I1(duty_23__N_3672[14]), .I2(n29_adj_4717), 
            .I3(GND_net), .O(n50502));   // verilog/motorControl.v(36[10:25])
    defparam i35549_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35176_4_lut (.I0(n33_adj_4723), .I1(n31_adj_4718), .I2(n29_adj_4717), 
            .I3(n49823), .O(n50128));
    defparam i35176_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35632_4_lut (.I0(n30_adj_4734), .I1(n10_adj_4733), .I2(n35_adj_4720), 
            .I3(n50123), .O(n50585));   // verilog/motorControl.v(36[10:25])
    defparam i35632_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35280_3_lut (.I0(n50502), .I1(duty_23__N_3672[15]), .I2(n31_adj_4718), 
            .I3(GND_net), .O(n50232));   // verilog/motorControl.v(36[10:25])
    defparam i35280_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35694_4_lut (.I0(n50232), .I1(n50585), .I2(n35_adj_4720), 
            .I3(n50128), .O(n50647));   // verilog/motorControl.v(36[10:25])
    defparam i35694_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35695_3_lut (.I0(n50647), .I1(duty_23__N_3672[18]), .I2(n37_adj_4716), 
            .I3(GND_net), .O(n50648));   // verilog/motorControl.v(36[10:25])
    defparam i35695_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35691_3_lut (.I0(n50648), .I1(duty_23__N_3672[19]), .I2(n39_adj_4713), 
            .I3(GND_net), .O(n50644));   // verilog/motorControl.v(36[10:25])
    defparam i35691_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35165_4_lut (.I0(n43_adj_4719), .I1(n41_adj_4714), .I2(n39_adj_4713), 
            .I3(n50603), .O(n50117));
    defparam i35165_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35656_4_lut (.I0(n50486), .I1(n50487), .I2(n45_adj_4715), 
            .I3(n50115), .O(n50609));   // verilog/motorControl.v(36[10:25])
    defparam i35656_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35286_3_lut (.I0(n50644), .I1(duty_23__N_3672[20]), .I2(n41_adj_4714), 
            .I3(GND_net), .O(n50238));   // verilog/motorControl.v(36[10:25])
    defparam i35286_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i418_2_lut (.I0(\Kp[8] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n621_adj_4653));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i418_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i83_2_lut (.I0(\Kp[1] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n122_adj_4651));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i83_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i36_2_lut (.I0(\Kp[0] ), .I1(n1[17]), .I2(GND_net), 
            .I3(GND_net), .O(n53_adj_4650));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i36_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35658_4_lut (.I0(n50238), .I1(n50609), .I2(n45_adj_4715), 
            .I3(n50117), .O(n50611));   // verilog/motorControl.v(36[10:25])
    defparam i35658_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35659_3_lut (.I0(n50611), .I1(PWMLimit[23]), .I2(duty_23__N_3672[23]), 
            .I3(GND_net), .O(duty_23__N_3671));   // verilog/motorControl.v(36[10:25])
    defparam i35659_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 LessThan_15_i41_2_lut (.I0(duty_23__N_3672[20]), .I1(n257[20]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4739));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i41_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i39_2_lut (.I0(duty_23__N_3672[19]), .I1(n257[19]), 
            .I2(GND_net), .I3(GND_net), .O(n39_adj_4740));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i39_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i45_2_lut (.I0(duty_23__N_3672[22]), .I1(n257[22]), 
            .I2(GND_net), .I3(GND_net), .O(n45_adj_4741));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i45_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i43_2_lut (.I0(duty_23__N_3672[21]), .I1(n257[21]), 
            .I2(GND_net), .I3(GND_net), .O(n43_adj_4742));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i43_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i37_2_lut (.I0(duty_23__N_3672[18]), .I1(n257[18]), 
            .I2(GND_net), .I3(GND_net), .O(n37_adj_4743));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i37_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i29_2_lut (.I0(duty_23__N_3672[14]), .I1(n257[14]), 
            .I2(GND_net), .I3(GND_net), .O(n29_adj_4744));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i29_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i31_2_lut (.I0(duty_23__N_3672[15]), .I1(n257[15]), 
            .I2(GND_net), .I3(GND_net), .O(n31_adj_4745));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i31_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i21_2_lut (.I0(duty_23__N_3672[10]), .I1(n257[10]), 
            .I2(GND_net), .I3(GND_net), .O(n21_adj_4746));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i21_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i23_2_lut (.I0(duty_23__N_3672[11]), .I1(n257[11]), 
            .I2(GND_net), .I3(GND_net), .O(n23_adj_4747));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i23_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i25_2_lut (.I0(duty_23__N_3672[12]), .I1(n257[12]), 
            .I2(GND_net), .I3(GND_net), .O(n25_adj_4748));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i25_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i17_2_lut (.I0(duty_23__N_3672[8]), .I1(n257[8]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4749));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i17_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i19_2_lut (.I0(duty_23__N_3672[9]), .I1(n257[9]), 
            .I2(GND_net), .I3(GND_net), .O(n19_adj_4750));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i19_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i9_2_lut (.I0(duty_23__N_3672[4]), .I1(n257[4]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4751));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i9_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i35_2_lut (.I0(duty_23__N_3672[17]), .I1(n257[17]), 
            .I2(GND_net), .I3(GND_net), .O(n35_adj_4752));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i35_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i33_2_lut (.I0(duty_23__N_3672[16]), .I1(n257[16]), 
            .I2(GND_net), .I3(GND_net), .O(n33_adj_4753));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i33_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i11_2_lut (.I0(duty_23__N_3672[5]), .I1(n257[5]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4754));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i11_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 LessThan_15_i13_2_lut (.I0(duty_23__N_3672[6]), .I1(n257[6]), 
            .I2(GND_net), .I3(GND_net), .O(n13_adj_4755));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i13_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i25858_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[20]), .I2(n38876), 
            .I3(n19077[0]), .O(n4_adj_4546));   // verilog/motorControl.v(34[16:22])
    defparam i25858_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[20]), .I2(n19077[0]), 
            .I3(n38876), .O(n19060[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h8778;
    SB_LUT4 i25845_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n19060[0]));   // verilog/motorControl.v(34[16:22])
    defparam i25845_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i25847_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[21]), .I2(n1[20]), 
            .I3(\Kp[1] ), .O(n38876));   // verilog/motorControl.v(34[16:22])
    defparam i25847_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 LessThan_15_i15_2_lut (.I0(duty_23__N_3672[7]), .I1(n257[7]), 
            .I2(GND_net), .I3(GND_net), .O(n15_adj_4756));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i15_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i25881_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[19]), .I2(n38901), 
            .I3(n19060[0]), .O(n4_adj_4524));   // verilog/motorControl.v(34[16:22])
    defparam i25881_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1531 (.I0(\Kp[2] ), .I1(n1[19]), .I2(n19060[0]), 
            .I3(n38901), .O(n19029[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1531.LUT_INIT = 16'h8778;
    SB_LUT4 i25868_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(n1[19]), 
            .I3(\Kp[1] ), .O(n19029[0]));   // verilog/motorControl.v(34[16:22])
    defparam i25868_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i25870_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[20]), .I2(n1[19]), 
            .I3(\Kp[1] ), .O(n38901));   // verilog/motorControl.v(34[16:22])
    defparam i25870_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i25920_3_lut_4_lut (.I0(\Kp[3] ), .I1(n1[18]), .I2(n4_adj_4757), 
            .I3(n19029[1]), .O(n6_adj_4514));   // verilog/motorControl.v(34[16:22])
    defparam i25920_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1532 (.I0(\Kp[3] ), .I1(n1[18]), .I2(n19029[1]), 
            .I3(n4_adj_4757), .O(n18980[2]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1532.LUT_INIT = 16'h8778;
    SB_LUT4 LessThan_15_i27_2_lut (.I0(duty_23__N_3672[13]), .I1(n257[13]), 
            .I2(GND_net), .I3(GND_net), .O(n27_adj_4758));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i27_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35149_4_lut (.I0(n21_adj_4746), .I1(n19_adj_4750), .I2(n17_adj_4749), 
            .I3(n9_adj_4751), .O(n50101));
    defparam i35149_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i2_3_lut_4_lut_adj_1533 (.I0(\Kp[2] ), .I1(n1[18]), .I2(n19029[0]), 
            .I3(n38935), .O(n18980[1]));   // verilog/motorControl.v(34[16:22])
    defparam i2_3_lut_4_lut_adj_1533.LUT_INIT = 16'h8778;
    SB_LUT4 i35141_4_lut (.I0(n27_adj_4758), .I1(n15_adj_4756), .I2(n13_adj_4755), 
            .I3(n11_adj_4754), .O(n50093));
    defparam i35141_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 LessThan_15_i12_3_lut (.I0(n257[7]), .I1(n257[16]), .I2(n33_adj_4753), 
            .I3(GND_net), .O(n12_adj_4759));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i10_3_lut (.I0(n257[5]), .I1(n257[6]), .I2(n13_adj_4755), 
            .I3(GND_net), .O(n10_adj_4760));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i30_3_lut (.I0(n12_adj_4759), .I1(n257[17]), .I2(n35_adj_4752), 
            .I3(GND_net), .O(n30_adj_4761));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i30_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i25912_3_lut_4_lut (.I0(\Kp[2] ), .I1(n1[18]), .I2(n38935), 
            .I3(n19029[0]), .O(n4_adj_4757));   // verilog/motorControl.v(34[16:22])
    defparam i25912_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i25899_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n18980[0]));   // verilog/motorControl.v(34[16:22])
    defparam i25899_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i20700_2_lut (.I0(n1[7]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[7]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20700_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i25901_2_lut_3_lut_4_lut (.I0(\Kp[0] ), .I1(n1[19]), .I2(n1[18]), 
            .I3(\Kp[1] ), .O(n38935));   // verilog/motorControl.v(34[16:22])
    defparam i25901_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i35384_4_lut (.I0(n13_adj_4755), .I1(n11_adj_4754), .I2(n9_adj_4751), 
            .I3(n50111), .O(n50337));
    defparam i35384_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35380_4_lut (.I0(n19_adj_4750), .I1(n17_adj_4749), .I2(n15_adj_4756), 
            .I3(n50337), .O(n50333));
    defparam i35380_4_lut.LUT_INIT = 16'heeef;
    SB_LUT4 i35646_4_lut (.I0(n25_adj_4748), .I1(n23_adj_4747), .I2(n21_adj_4746), 
            .I3(n50333), .O(n50599));
    defparam i35646_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i35482_4_lut (.I0(n31_adj_4745), .I1(n29_adj_4744), .I2(n27_adj_4758), 
            .I3(n50599), .O(n50435));
    defparam i35482_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i35674_4_lut (.I0(n37_adj_4743), .I1(n35_adj_4752), .I2(n33_adj_4753), 
            .I3(n50435), .O(n50627));
    defparam i35674_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 LessThan_15_i16_3_lut (.I0(n257[9]), .I1(n257[21]), .I2(n43_adj_4742), 
            .I3(GND_net), .O(n16_adj_4762));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35542_3_lut (.I0(n6_adj_4670), .I1(n257[10]), .I2(n21_adj_4746), 
            .I3(GND_net), .O(n50495));   // verilog/motorControl.v(38[19:35])
    defparam i35542_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35543_3_lut (.I0(n50495), .I1(n257[11]), .I2(n23_adj_4747), 
            .I3(GND_net), .O(n50496));   // verilog/motorControl.v(38[19:35])
    defparam i35543_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i8_3_lut (.I0(n257[4]), .I1(n257[8]), .I2(n17_adj_4749), 
            .I3(GND_net), .O(n8_adj_4763));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i24_3_lut (.I0(n16_adj_4762), .I1(n257[22]), .I2(n45_adj_4741), 
            .I3(GND_net), .O(n24_adj_4764));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20699_2_lut (.I0(n1[8]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[8]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20699_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35125_4_lut (.I0(n43_adj_4742), .I1(n25_adj_4748), .I2(n23_adj_4747), 
            .I3(n50101), .O(n50077));
    defparam i35125_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35536_4_lut (.I0(n24_adj_4764), .I1(n8_adj_4763), .I2(n45_adj_4741), 
            .I3(n50075), .O(n50489));   // verilog/motorControl.v(38[19:35])
    defparam i35536_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35288_3_lut (.I0(n50496), .I1(n257[12]), .I2(n25_adj_4748), 
            .I3(GND_net), .O(n50240));   // verilog/motorControl.v(38[19:35])
    defparam i35288_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 LessThan_15_i4_4_lut (.I0(duty_23__N_3672[0]), .I1(n257[1]), 
            .I2(duty_23__N_3672[1]), .I3(n257[0]), .O(n4_adj_4765));   // verilog/motorControl.v(38[19:35])
    defparam LessThan_15_i4_4_lut.LUT_INIT = 16'h4d0c;
    SB_LUT4 i35540_3_lut (.I0(n4_adj_4765), .I1(n257[13]), .I2(n27_adj_4758), 
            .I3(GND_net), .O(n50493));   // verilog/motorControl.v(38[19:35])
    defparam i35540_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35541_3_lut (.I0(n50493), .I1(n257[14]), .I2(n29_adj_4744), 
            .I3(GND_net), .O(n50494));   // verilog/motorControl.v(38[19:35])
    defparam i35541_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35136_4_lut (.I0(n33_adj_4753), .I1(n31_adj_4745), .I2(n29_adj_4744), 
            .I3(n50093), .O(n50088));
    defparam i35136_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35634_4_lut (.I0(n30_adj_4761), .I1(n10_adj_4760), .I2(n35_adj_4752), 
            .I3(n50086), .O(n50587));   // verilog/motorControl.v(38[19:35])
    defparam i35634_4_lut.LUT_INIT = 16'haaac;
    SB_LUT4 i35290_3_lut (.I0(n50494), .I1(n257[15]), .I2(n31_adj_4745), 
            .I3(GND_net), .O(n50242));   // verilog/motorControl.v(38[19:35])
    defparam i35290_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35696_4_lut (.I0(n50242), .I1(n50587), .I2(n35_adj_4752), 
            .I3(n50088), .O(n50649));   // verilog/motorControl.v(38[19:35])
    defparam i35696_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35697_3_lut (.I0(n50649), .I1(n257[18]), .I2(n37_adj_4743), 
            .I3(GND_net), .O(n50650));   // verilog/motorControl.v(38[19:35])
    defparam i35697_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35687_3_lut (.I0(n50650), .I1(n257[19]), .I2(n39_adj_4740), 
            .I3(GND_net), .O(n50640));   // verilog/motorControl.v(38[19:35])
    defparam i35687_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35127_4_lut (.I0(n43_adj_4742), .I1(n41_adj_4739), .I2(n39_adj_4740), 
            .I3(n50627), .O(n50079));
    defparam i35127_4_lut.LUT_INIT = 16'haaab;
    SB_LUT4 i35660_4_lut (.I0(n50240), .I1(n50489), .I2(n45_adj_4741), 
            .I3(n50077), .O(n50613));   // verilog/motorControl.v(38[19:35])
    defparam i35660_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35296_3_lut (.I0(n50640), .I1(n257[20]), .I2(n41_adj_4739), 
            .I3(GND_net), .O(n50248));   // verilog/motorControl.v(38[19:35])
    defparam i35296_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35662_4_lut (.I0(n50248), .I1(n50613), .I2(n45_adj_4741), 
            .I3(n50079), .O(n50615));   // verilog/motorControl.v(38[19:35])
    defparam i35662_4_lut.LUT_INIT = 16'hccca;
    SB_LUT4 i35663_3_lut (.I0(n50615), .I1(duty_23__N_3672[23]), .I2(n257[23]), 
            .I3(GND_net), .O(n256_adj_4552));   // verilog/motorControl.v(38[19:35])
    defparam i35663_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 mux_17_i1_3_lut (.I0(duty_23__N_3672[0]), .I1(n257[0]), .I2(n256_adj_4552), 
            .I3(GND_net), .O(duty_23__N_3647[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam mux_17_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 duty_23__I_0_i1_3_lut (.I0(duty_23__N_3647[0]), .I1(PWMLimit[0]), 
            .I2(duty_23__N_3671), .I3(GND_net), .O(duty_23__N_3548[0]));   // verilog/motorControl.v(38[16] 40[10])
    defparam duty_23__I_0_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mult_10_i506_2_lut (.I0(\Kp[10] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n752_adj_4371));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i506_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i277_2_lut (.I0(\Kp[5] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n411));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i277_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i10_1_lut (.I0(PWMLimit[9]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[9]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i10_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i102_2_lut (.I0(\Kp[2] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n150_adj_4361));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i102_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i555_2_lut (.I0(\Kp[11] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n825_adj_4360));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i555_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i151_2_lut (.I0(\Kp[3] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n223_adj_4358));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i151_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i414_2_lut (.I0(\Kp[8] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n615));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i414_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i11_1_lut (.I0(PWMLimit[10]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[10]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i11_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i12_1_lut (.I0(PWMLimit[11]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[11]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i12_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_10_i326_2_lut (.I0(\Kp[6] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n484));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i326_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i132_2_lut (.I0(\Kp[2] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n195_adj_4646));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i132_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20698_2_lut (.I0(n1[9]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[9]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20698_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i59_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n86_adj_4645));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i59_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i375_2_lut (.I0(\Kp[7] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n557));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i375_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i12_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [5]), 
            .I2(GND_net), .I3(GND_net), .O(n17_adj_4644));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i12_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i424_2_lut (.I0(\Kp[8] ), .I1(n1[15]), .I2(GND_net), 
            .I3(GND_net), .O(n630));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i424_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20697_2_lut (.I0(n1[10]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[10]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20697_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i55_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n80));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i55_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i8_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [3]), 
            .I2(GND_net), .I3(GND_net), .O(n11_adj_4355));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i8_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i13_1_lut (.I0(PWMLimit[12]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[12]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i13_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 unary_minus_16_inv_0_i14_1_lut (.I0(PWMLimit[13]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[13]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i14_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i65_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n95));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i65_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i18_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [8]), 
            .I2(GND_net), .I3(GND_net), .O(n26_adj_4354));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i18_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i604_2_lut (.I0(\Kp[12] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n898_adj_4353));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i604_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i114_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n168));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i114_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 IntegralLimit_23__I_0_i8_3_lut_3_lut (.I0(IntegralLimit[4]), .I1(IntegralLimit[8]), 
            .I2(\PID_CONTROLLER.integral [8]), .I3(GND_net), .O(n8_adj_4432));   // verilog/motorControl.v(31[10:34])
    defparam IntegralLimit_23__I_0_i8_3_lut_3_lut.LUT_INIT = 16'h8e8e;
    SB_LUT4 i25827_3_lut_4_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [18]), 
            .I2(n4_adj_4766), .I3(n19005[1]), .O(n6_adj_4372));   // verilog/motorControl.v(34[25:36])
    defparam i25827_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1534 (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [18]), 
            .I2(n19005[1]), .I3(n4_adj_4766), .O(n18945[2]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1534.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_1535 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [18]), 
            .I2(n19005[0]), .I3(n38833), .O(n18945[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1535.LUT_INIT = 16'h8778;
    SB_LUT4 i25819_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [18]), 
            .I2(n38833), .I3(n19005[0]), .O(n4_adj_4766));   // verilog/motorControl.v(34[25:36])
    defparam i25819_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i25806_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3572 [18]), .I3(\Ki[1] ), 
            .O(n18945[0]));   // verilog/motorControl.v(34[25:36])
    defparam i25806_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i25808_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [19]), 
            .I2(\PID_CONTROLLER.integral_23__N_3572 [18]), .I3(\Ki[1] ), 
            .O(n38833));   // verilog/motorControl.v(34[25:36])
    defparam i25808_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i25775_2_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [20]), 
            .I2(\Ki[1] ), .I3(\PID_CONTROLLER.integral_23__N_3572 [19]), 
            .O(n19005[0]));   // verilog/motorControl.v(34[25:36])
    defparam i25775_2_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i25750_3_lut_4_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [20]), 
            .I2(n38758), .I3(n19069[0]), .O(n4_adj_4385));   // verilog/motorControl.v(34[25:36])
    defparam i25750_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i2_3_lut_4_lut_adj_1536 (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [20]), 
            .I2(n19069[0]), .I3(n38758), .O(n19045[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1536.LUT_INIT = 16'h8778;
    SB_LUT4 i2_3_lut_4_lut_adj_1537 (.I0(n62), .I1(n131), .I2(n19045[0]), 
            .I3(n204), .O(n19005[1]));   // verilog/motorControl.v(34[25:36])
    defparam i2_3_lut_4_lut_adj_1537.LUT_INIT = 16'h8778;
    SB_LUT4 i25788_3_lut_4_lut (.I0(n62), .I1(n131), .I2(n204), .I3(n19045[0]), 
            .O(n4_adj_4376));   // verilog/motorControl.v(34[25:36])
    defparam i25788_3_lut_4_lut.LUT_INIT = 16'hf880;
    SB_LUT4 i25737_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3572 [20]), .I3(\Ki[1] ), 
            .O(n19045[0]));   // verilog/motorControl.v(34[25:36])
    defparam i25737_2_lut_3_lut_4_lut.LUT_INIT = 16'h7888;
    SB_LUT4 i25739_2_lut_3_lut_4_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [21]), 
            .I2(\PID_CONTROLLER.integral_23__N_3572 [20]), .I3(\Ki[1] ), 
            .O(n38758));   // verilog/motorControl.v(34[25:36])
    defparam i25739_2_lut_3_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i20696_2_lut (.I0(n1[11]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[11]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20696_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i181_2_lut (.I0(\Kp[3] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n268_adj_4636));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i181_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i230_2_lut (.I0(\Kp[4] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n341_adj_4635));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i230_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i108_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n159_adj_4634));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i108_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i157_2_lut (.I0(\Ki[3] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n232_adj_4633));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i157_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i279_2_lut (.I0(\Kp[5] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n414_adj_4632));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i279_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i206_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n305_adj_4631));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i206_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20695_2_lut (.I0(n1[12]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[12]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20695_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i467_2_lut (.I0(\Kp[9] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n694_adj_4630));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i467_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i463_2_lut (.I0(\Kp[9] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n688));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i463_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i328_2_lut (.I0(\Kp[6] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n487_adj_4629));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i328_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i377_2_lut (.I0(\Kp[7] ), .I1(n1[16]), .I2(GND_net), 
            .I3(GND_net), .O(n560_adj_4628));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i377_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i516_2_lut (.I0(\Kp[10] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n767_adj_4627));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i516_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i255_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n378_adj_4626));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i255_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i565_2_lut (.I0(\Kp[11] ), .I1(n1[12]), .I2(GND_net), 
            .I3(GND_net), .O(n840_adj_4625));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i565_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i204_2_lut (.I0(\Kp[4] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n302_adj_4624));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i204_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i304_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n451_adj_4623));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i304_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20694_2_lut (.I0(n1[13]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[13]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20694_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i512_2_lut (.I0(\Kp[10] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n761));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i512_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i353_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n524_adj_4621));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i353_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i402_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n597_adj_4620));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i402_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i561_2_lut (.I0(\Kp[11] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n834));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i561_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i253_2_lut (.I0(\Kp[5] ), .I1(n1[3]), .I2(GND_net), 
            .I3(GND_net), .O(n375_adj_4619));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i253_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i451_2_lut (.I0(\Ki[9] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [4]), 
            .I2(GND_net), .I3(GND_net), .O(n670_adj_4618));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i451_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i610_2_lut (.I0(\Kp[12] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n907));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i610_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i20693_2_lut (.I0(n1[14]), .I1(\PID_CONTROLLER.integral_23__N_3620 ), 
            .I2(GND_net), .I3(GND_net), .O(n3616[14]));   // verilog/motorControl.v(31[7] 33[10])
    defparam i20693_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i659_2_lut (.I0(\Kp[13] ), .I1(n1[10]), .I2(GND_net), 
            .I3(GND_net), .O(n980));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i659_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i396_2_lut (.I0(\Kp[8] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n588_adj_4712));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i396_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i445_2_lut (.I0(\Kp[9] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n661_adj_4711));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i445_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i212_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n314_adj_4710));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i212_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i494_2_lut (.I0(\Kp[10] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n734_adj_4709));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i494_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i63_2_lut (.I0(\Kp[1] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n92_adj_4708));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i63_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i16_2_lut (.I0(\Kp[0] ), .I1(n1[7]), .I2(GND_net), 
            .I3(GND_net), .O(n23_adj_4707));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i16_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i543_2_lut (.I0(\Kp[11] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n807_adj_4706));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i543_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i592_2_lut (.I0(\Kp[12] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n880_adj_4705));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i592_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i641_2_lut (.I0(\Kp[13] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n953_adj_4704));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i641_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i690_2_lut (.I0(\Kp[14] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1026_adj_4703));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i690_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i112_2_lut (.I0(\Kp[2] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n165_adj_4702));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i112_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i739_2_lut (.I0(\Kp[15] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n1099_adj_4701));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i739_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i261_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n387_adj_4700));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i261_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i161_2_lut (.I0(\Kp[3] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n238_adj_4699));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i161_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i202_2_lut (.I0(\Ki[4] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n299_adj_4698));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i202_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i210_2_lut (.I0(\Kp[4] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n311_adj_4697));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i210_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i259_2_lut (.I0(\Kp[5] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n384_adj_4696));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i259_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i251_2_lut (.I0(\Ki[5] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n372_adj_4695));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i251_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i308_2_lut (.I0(\Kp[6] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n457_adj_4694));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i308_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i75_2_lut (.I0(\Ki[1] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n110_adj_4693));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i75_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i28_2_lut (.I0(\Ki[0] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [13]), 
            .I2(GND_net), .I3(GND_net), .O(n41_adj_4692));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i28_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i310_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n460_adj_4691));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i310_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i357_2_lut (.I0(\Kp[7] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n530_adj_4690));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i357_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i16_1_lut (.I0(PWMLimit[15]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[15]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i16_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i300_2_lut (.I0(\Ki[6] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n445_adj_4688));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i300_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i359_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n533_adj_4687));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i359_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i406_2_lut (.I0(\Kp[8] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n603_adj_4686));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i406_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i455_2_lut (.I0(\Kp[9] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n676_adj_4685));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i455_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i408_2_lut (.I0(\Ki[8] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [7]), 
            .I2(GND_net), .I3(GND_net), .O(n606_adj_4684));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i408_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 unary_minus_16_inv_0_i17_1_lut (.I0(PWMLimit[16]), .I1(GND_net), 
            .I2(GND_net), .I3(GND_net), .O(n1_adj_4767[16]));   // verilog/motorControl.v(39[18:27])
    defparam unary_minus_16_inv_0_i17_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 mult_11_i124_2_lut (.I0(\Ki[2] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [12]), 
            .I2(GND_net), .I3(GND_net), .O(n183_adj_4682));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i124_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_11_i349_2_lut (.I0(\Ki[7] ), .I1(\PID_CONTROLLER.integral_23__N_3572 [2]), 
            .I2(GND_net), .I3(GND_net), .O(n518_adj_4681));   // verilog/motorControl.v(34[25:36])
    defparam mult_11_i349_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i504_2_lut (.I0(\Kp[10] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n749_adj_4680));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i504_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i553_2_lut (.I0(\Kp[11] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n822_adj_4679));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i553_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i51_2_lut (.I0(\Kp[1] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n74_adj_4678));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i51_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i4_2_lut (.I0(\Kp[0] ), .I1(n1[1]), .I2(GND_net), 
            .I3(GND_net), .O(n5_adj_4677));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i4_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i100_2_lut (.I0(\Kp[2] ), .I1(n1[0]), .I2(GND_net), 
            .I3(GND_net), .O(n147_adj_4676));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i100_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 mult_10_i602_2_lut (.I0(\Kp[12] ), .I1(n1[6]), .I2(GND_net), 
            .I3(GND_net), .O(n895_adj_4675));   // verilog/motorControl.v(34[16:22])
    defparam mult_10_i602_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module coms
//

module coms (rx_data, CLK_c, \data_out_frame[9] , \data_out_frame[4] , 
            GND_net, \data_out_frame[8] , \data_out_frame[13] , \data_out_frame[18] , 
            \data_out_frame[16] , \data_out_frame[20] , \data_out_frame[25] , 
            \data_out_frame[11] , \data_out_frame[15] , \data_out_frame[23] , 
            \data_out_frame[14] , \data_out_frame[7] , \data_out_frame[12] , 
            \data_out_frame[5] , \data_out_frame[10] , \data_out_frame[17] , 
            \data_out_frame[19] , \data_out_frame[6] , \byte_transmit_counter[2] , 
            \FRAME_MATCHER.state , \data_in_frame[2] , \data_in_frame[1] , 
            \data_in_frame[8] , n44058, n33302, n23831, n46759, n40, 
            n33308, n5728, n44035, n61, n76, n2482, n29985, n63, 
            n51904, \FRAME_MATCHER.i_31__N_2524 , n3303, n5, \FRAME_MATCHER.i_31__N_2526 , 
            n4452, n7, \data_in_frame[9] , \displacement[17] , n23935, 
            rx_data_ready, n33298, \FRAME_MATCHER.state[0] , n73, setpoint, 
            \byte_transmit_counter[0] , tx_transmit_N_3413, \data_in_frame[10] , 
            \FRAME_MATCHER.i[31] , \data_in_frame[11] , n28284, control_mode, 
            n28283, n28282, n28281, n28280, n28279, n771, n26687, 
            n1476, n28278, n28277, PWMLimit, n28276, n28275, n28274, 
            n28273, n26489, \data_in[3] , \data_in[1] , \data_in[0] , 
            \data_in[2] , n28272, n28271, \data_in_frame[12] , \data_in_frame[3] , 
            \data_in_frame[13] , n28270, n28269, n28268, n28267, n28266, 
            n28265, n28264, n28263, n28262, n28261, n28260, n28259, 
            n28258, n28257, n28256, n28255, n51636, n51637, \state[2] , 
            \state[3] , n10, n27771, n43485, n49817, \data_out_frame[24] , 
            n51546, \data_out_frame[18][0] , n28214, n27546, DE_c, 
            LED_c, n74, n28213, n44240, n28211, neopxl_color, n28210, 
            \Ki[0] , n28209, \Kp[0] , n28208, n28759, IntegralLimit, 
            n28758, n28757, n28756, n28755, n28754, n28753, n28752, 
            n28751, n28750, n28749, n28748, n28747, n28746, n28745, 
            n28744, n28743, n28742, n28741, n28740, n28739, n28738, 
            n28737, n28736, n28735, n28734, n28733, n28732, n28731, 
            n28730, n28729, n28728, n28727, \data_in_frame[5] , \data_in_frame[6] , 
            \data_in_frame[4] , n28726, n28725, n28724, n28723, n28722, 
            n28721, n28720, n28719, n28718, n28717, n28716, n28715, 
            n28714, n28713, n28712, n28711, n28710, n28709, n28708, 
            n28707, n28706, n28705, \Kp[1] , n28704, \Kp[2] , n28703, 
            \Kp[3] , n28702, \Kp[4] , n28701, \Kp[5] , n28700, \Kp[6] , 
            n28699, \Kp[7] , n28698, \Kp[8] , n28697, \Kp[9] , n28696, 
            \Kp[10] , n28695, \Kp[11] , n28694, \Kp[12] , n28693, 
            \Kp[13] , n28692, \Kp[14] , n28691, \Kp[15] , n28690, 
            \Ki[1] , n28689, \Ki[2] , n28688, \Ki[3] , n28687, \Ki[4] , 
            n28686, \Ki[5] , n28685, \Ki[6] , n28684, \Ki[7] , n28683, 
            \Ki[8] , n28682, \Ki[9] , n28681, \Ki[10] , n28680, 
            \Ki[11] , n28679, \Ki[12] , n28678, \Ki[13] , n28677, 
            \Ki[14] , n28676, \Ki[15] , n28675, n28674, n28673, 
            n28672, n28671, n28670, n28669, n28668, n28667, n28666, 
            n28665, n28664, n28663, n28662, n28661, n28660, n28659, 
            n28658, n28657, n28656, n28655, n28654, n28653, n28652, 
            n28651, n28650, n28649, n28648, n28647, n28646, n28645, 
            n28644, n28643, n28642, n28641, n28640, n28639, n28638, 
            n28637, n28636, n28635, n28634, n28633, n28632, n28631, 
            n28630, n28629, n28628, n28627, n28626, n28625, n28624, 
            n28623, n28622, n28621, n28620, n28619, n28618, n28617, 
            n28616, n28615, n28614, n28613, n28612, n28611, n28610, 
            n28609, n28608, n28607, n28606, n28605, n28604, n28603, 
            n28602, n28601, n28600, n28599, n28598, n28597, n28596, 
            n28595, n28594, n28593, n28592, n28591, n28590, n28589, 
            n28588, n28587, n28586, n28585, n28584, n28583, n28582, 
            n28581, n28580, n28579, n28578, n28577, n28576, n28575, 
            n28574, n28573, n28572, n28571, n28570, n28569, n28568, 
            n28567, n28566, n28565, n28564, n28563, n28561, \data_out_frame[18][2] , 
            n28560, n28559, n28558, n28557, n28556, n28555, n28554, 
            n28553, n28552, n28551, n28550, n28549, n28548, n28547, 
            n28546, n28545, n28544, n28543, n28542, n28541, n28540, 
            n28539, n28538, n28537, n28536, n28535, n28534, n28533, 
            n28532, n28531, n28530, n28529, n28528, n28527, n28526, 
            n28525, n28524, n28523, n28522, n28189, n28521, n28520, 
            n28519, n28518, n28517, n28516, n28515, n28514, n28513, 
            n28512, n28511, n28510, n28509, n28508, n28507, n28506, 
            n28505, n28504, n28503, n28502, n28501, n28500, n28499, 
            n28498, n28497, n28496, n28495, n28494, n28493, n46360, 
            ID, n39, \state[0] , n6014, n44092, n44436, n44685, 
            n26881, n49818, n49819, n15, tx_o, VCC_net, tx_enable, 
            r_SM_Main, \r_SM_Main_2__N_3442[2] , \r_Bit_Index[0] , n26629, 
            n4, r_Rx_Data, RX_N_10, n27846, n28246, n43659, n28250, 
            n28223, n28222, n28221, n28219, n28218, n43968, n28203, 
            n28202, n44048, n4_adj_10, n4_adj_11, n26624, n33765) /* synthesis syn_module_defined=1 */ ;
    output [7:0]rx_data;
    input CLK_c;
    output [7:0]\data_out_frame[9] ;
    output [7:0]\data_out_frame[4] ;
    input GND_net;
    output [7:0]\data_out_frame[8] ;
    output [7:0]\data_out_frame[13] ;
    output [7:0]\data_out_frame[18] ;
    output [7:0]\data_out_frame[16] ;
    output [7:0]\data_out_frame[20] ;
    output [7:0]\data_out_frame[25] ;
    output [7:0]\data_out_frame[11] ;
    output [7:0]\data_out_frame[15] ;
    output [7:0]\data_out_frame[23] ;
    output [7:0]\data_out_frame[14] ;
    output [7:0]\data_out_frame[7] ;
    output [7:0]\data_out_frame[12] ;
    output [7:0]\data_out_frame[5] ;
    output [7:0]\data_out_frame[10] ;
    output [7:0]\data_out_frame[17] ;
    output [7:0]\data_out_frame[19] ;
    output [7:0]\data_out_frame[6] ;
    output \byte_transmit_counter[2] ;
    output [31:0]\FRAME_MATCHER.state ;
    output [7:0]\data_in_frame[2] ;
    output [7:0]\data_in_frame[1] ;
    output [7:0]\data_in_frame[8] ;
    input n44058;
    output n33302;
    output n23831;
    output n46759;
    output n40;
    output n33308;
    output n5728;
    output n44035;
    output n61;
    output n76;
    output n2482;
    output n29985;
    output n63;
    output n51904;
    output \FRAME_MATCHER.i_31__N_2524 ;
    output n3303;
    output n5;
    output \FRAME_MATCHER.i_31__N_2526 ;
    output n4452;
    output n7;
    output [7:0]\data_in_frame[9] ;
    input \displacement[17] ;
    output n23935;
    output rx_data_ready;
    output n33298;
    output \FRAME_MATCHER.state[0] ;
    output n73;
    output [23:0]setpoint;
    output \byte_transmit_counter[0] ;
    output tx_transmit_N_3413;
    output [7:0]\data_in_frame[10] ;
    output \FRAME_MATCHER.i[31] ;
    output [7:0]\data_in_frame[11] ;
    input n28284;
    output [7:0]control_mode;
    input n28283;
    input n28282;
    input n28281;
    input n28280;
    input n28279;
    output n771;
    output n26687;
    output n1476;
    input n28278;
    input n28277;
    output [23:0]PWMLimit;
    input n28276;
    input n28275;
    input n28274;
    input n28273;
    output n26489;
    output [7:0]\data_in[3] ;
    output [7:0]\data_in[1] ;
    output [7:0]\data_in[0] ;
    output [7:0]\data_in[2] ;
    input n28272;
    input n28271;
    output [7:0]\data_in_frame[12] ;
    output [7:0]\data_in_frame[3] ;
    output [7:0]\data_in_frame[13] ;
    input n28270;
    input n28269;
    input n28268;
    input n28267;
    input n28266;
    input n28265;
    input n28264;
    input n28263;
    input n28262;
    input n28261;
    input n28260;
    input n28259;
    input n28258;
    input n28257;
    input n28256;
    input n28255;
    input n51636;
    input n51637;
    input \state[2] ;
    input \state[3] ;
    output n10;
    output n27771;
    input n43485;
    input n49817;
    output [7:0]\data_out_frame[24] ;
    output n51546;
    output \data_out_frame[18][0] ;
    input n28214;
    output n27546;
    output DE_c;
    output LED_c;
    output n74;
    input n28213;
    output n44240;
    input n28211;
    output [23:0]neopxl_color;
    input n28210;
    output \Ki[0] ;
    input n28209;
    output \Kp[0] ;
    input n28208;
    input n28759;
    output [23:0]IntegralLimit;
    input n28758;
    input n28757;
    input n28756;
    input n28755;
    input n28754;
    input n28753;
    input n28752;
    input n28751;
    input n28750;
    input n28749;
    input n28748;
    input n28747;
    input n28746;
    input n28745;
    input n28744;
    input n28743;
    input n28742;
    input n28741;
    input n28740;
    input n28739;
    input n28738;
    input n28737;
    input n28736;
    input n28735;
    input n28734;
    input n28733;
    input n28732;
    input n28731;
    input n28730;
    input n28729;
    input n28728;
    input n28727;
    output [7:0]\data_in_frame[5] ;
    output [7:0]\data_in_frame[6] ;
    output [7:0]\data_in_frame[4] ;
    input n28726;
    input n28725;
    input n28724;
    input n28723;
    input n28722;
    input n28721;
    input n28720;
    input n28719;
    input n28718;
    input n28717;
    input n28716;
    input n28715;
    input n28714;
    input n28713;
    input n28712;
    input n28711;
    input n28710;
    input n28709;
    input n28708;
    input n28707;
    input n28706;
    input n28705;
    output \Kp[1] ;
    input n28704;
    output \Kp[2] ;
    input n28703;
    output \Kp[3] ;
    input n28702;
    output \Kp[4] ;
    input n28701;
    output \Kp[5] ;
    input n28700;
    output \Kp[6] ;
    input n28699;
    output \Kp[7] ;
    input n28698;
    output \Kp[8] ;
    input n28697;
    output \Kp[9] ;
    input n28696;
    output \Kp[10] ;
    input n28695;
    output \Kp[11] ;
    input n28694;
    output \Kp[12] ;
    input n28693;
    output \Kp[13] ;
    input n28692;
    output \Kp[14] ;
    input n28691;
    output \Kp[15] ;
    input n28690;
    output \Ki[1] ;
    input n28689;
    output \Ki[2] ;
    input n28688;
    output \Ki[3] ;
    input n28687;
    output \Ki[4] ;
    input n28686;
    output \Ki[5] ;
    input n28685;
    output \Ki[6] ;
    input n28684;
    output \Ki[7] ;
    input n28683;
    output \Ki[8] ;
    input n28682;
    output \Ki[9] ;
    input n28681;
    output \Ki[10] ;
    input n28680;
    output \Ki[11] ;
    input n28679;
    output \Ki[12] ;
    input n28678;
    output \Ki[13] ;
    input n28677;
    output \Ki[14] ;
    input n28676;
    output \Ki[15] ;
    input n28675;
    input n28674;
    input n28673;
    input n28672;
    input n28671;
    input n28670;
    input n28669;
    input n28668;
    input n28667;
    input n28666;
    input n28665;
    input n28664;
    input n28663;
    input n28662;
    input n28661;
    input n28660;
    input n28659;
    input n28658;
    input n28657;
    input n28656;
    input n28655;
    input n28654;
    input n28653;
    input n28652;
    input n28651;
    input n28650;
    input n28649;
    input n28648;
    input n28647;
    input n28646;
    input n28645;
    input n28644;
    input n28643;
    input n28642;
    input n28641;
    input n28640;
    input n28639;
    input n28638;
    input n28637;
    input n28636;
    input n28635;
    input n28634;
    input n28633;
    input n28632;
    input n28631;
    input n28630;
    input n28629;
    input n28628;
    input n28627;
    input n28626;
    input n28625;
    input n28624;
    input n28623;
    input n28622;
    input n28621;
    input n28620;
    input n28619;
    input n28618;
    input n28617;
    input n28616;
    input n28615;
    input n28614;
    input n28613;
    input n28612;
    input n28611;
    input n28610;
    input n28609;
    input n28608;
    input n28607;
    input n28606;
    input n28605;
    input n28604;
    input n28603;
    input n28602;
    input n28601;
    input n28600;
    input n28599;
    input n28598;
    input n28597;
    input n28596;
    input n28595;
    input n28594;
    input n28593;
    input n28592;
    input n28591;
    input n28590;
    input n28589;
    input n28588;
    input n28587;
    input n28586;
    input n28585;
    input n28584;
    input n28583;
    input n28582;
    input n28581;
    input n28580;
    input n28579;
    input n28578;
    input n28577;
    input n28576;
    input n28575;
    input n28574;
    input n28573;
    input n28572;
    input n28571;
    input n28570;
    input n28569;
    input n28568;
    input n28567;
    input n28566;
    input n28565;
    input n28564;
    input n28563;
    input n28561;
    output \data_out_frame[18][2] ;
    input n28560;
    input n28559;
    input n28558;
    input n28557;
    input n28556;
    input n28555;
    input n28554;
    input n28553;
    input n28552;
    input n28551;
    input n28550;
    input n28549;
    input n28548;
    input n28547;
    input n28546;
    input n28545;
    input n28544;
    input n28543;
    input n28542;
    input n28541;
    input n28540;
    input n28539;
    input n28538;
    input n28537;
    input n28536;
    input n28535;
    input n28534;
    input n28533;
    input n28532;
    input n28531;
    input n28530;
    input n28529;
    input n28528;
    input n28527;
    input n28526;
    input n28525;
    input n28524;
    input n28523;
    input n28522;
    input n28189;
    input n28521;
    input n28520;
    input n28519;
    input n28518;
    input n28517;
    input n28516;
    input n28515;
    input n28514;
    input n28513;
    input n28512;
    input n28511;
    input n28510;
    input n28509;
    input n28508;
    input n28507;
    input n28506;
    input n28505;
    input n28504;
    input n28503;
    input n28502;
    input n28501;
    input n28500;
    input n28499;
    input n28498;
    input n28497;
    input n28496;
    input n28495;
    input n28494;
    input n28493;
    output n46360;
    input [7:0]ID;
    output n39;
    input \state[0] ;
    output n6014;
    output n44092;
    input n44436;
    input n44685;
    output n26881;
    input n49818;
    input n49819;
    input n15;
    output tx_o;
    input VCC_net;
    output tx_enable;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3442[2] ;
    output \r_Bit_Index[0] ;
    output n26629;
    output n4;
    output r_Rx_Data;
    input RX_N_10;
    output n27846;
    input n28246;
    input n43659;
    input n28250;
    input n28223;
    input n28222;
    input n28221;
    input n28219;
    input n28218;
    output n43968;
    input n28203;
    input n28202;
    input n44048;
    output n4_adj_10;
    output n4_adj_11;
    output n26624;
    output n33765;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    
    wire n34417, n44104;
    wire [7:0]\data_in_frame[7] ;   // verilog/coms.v(96[12:25])
    
    wire n28428, n28320;
    wire [7:0]\data_in_frame[21] ;   // verilog/coms.v(96[12:25])
    
    wire n28319, n28318, n28317, n44218, n28316, n44176, n27539, 
        n27558, n27407, n14, n44321, n10_c, n26226, n27110, n50682, 
        n27561, n44351, n6, n44697, n28429, n44333, n6_adj_4111, 
        n50676, n44509, n45876, n44518, n42312, n41225, n45674, 
        n44489, n27212, n14_adj_4112, n10_adj_4113, n44297, n41601, 
        n26380, n45778, n27603, n41540, n41615, n2;
    wire [31:0]\FRAME_MATCHER.i ;   // verilog/coms.v(115[11:12])
    
    wire n3, n11, n9, n44497, n42416, n42300, n44264, n44151, 
        n27484, n27093, n27666, n24830, n44721, n44597, n44258, 
        n1699, n42493, n44318, n41571, n26809, n46253, n44534, 
        n28430, n44621, n44612, n6_adj_4114, n44268, n14_adj_4115, 
        n26755, n26724, n44543, n44703, n15_c, n44700, n28431, 
        n26281, n44366, n44255, n15_adj_4116, n44471, n14_adj_4117, 
        n44201, n42346, n41486, n44491, n6_adj_4118, n2122, n46081, 
        n27152, n41597, n44727, n44576, n44600, n44215, n12, n44724, 
        n41455, n44204, n44285, n14_adj_4119, n10_adj_4120, n44609, 
        n1510, n27321, n44409, n6_adj_4121, n41589, n1794, n10_adj_4122, 
        n41553, n28432, n26846, n6_adj_4123, n44387, n44546, n10_adj_4124, 
        n44304, n28433, n27288, n14_adj_4125, n1519, n10_adj_4126, 
        n44198, n41480, n1516, n27220, n44477, n1168, n44384, 
        n44579, n24, n44559, n34, n44573, n22, n38, n26712, 
        n36, n37, n44330, n35, n42075;
    wire [7:0]n8825;
    
    wire n27787;
    wire [7:0]byte_transmit_counter;   // verilog/coms.v(102[12:33])
    
    wire n33303, n27269, n44342, n27403, n44630, n12_adj_4127, n42387, 
        n44136, n28434, n16, n17, n44224, n44139, n44606, n44582, 
        n10_adj_4128, n44461, n44524, n15_adj_4129, n14_adj_4130, 
        n42285, n42365, n44424, n42378, n44445, n28435, n44688, 
        n8, n42393, n44427, n42339, n34047, n44929, n27912, n44428, 
        n39109, n39110;
    wire [7:0]\data_in_frame[0] ;   // verilog/coms.v(96[12:25])
    
    wire n44373, n44261, n44142, Kp_23__N_869, n44271, n27356, n7_c, 
        n48791, n20, n27, n24_adj_4131, n27337, n30, n24120, n22_adj_4132, 
        n31, n48673;
    wire [31:0]\FRAME_MATCHER.state_31__N_2624 ;
    
    wire n33307, n81;
    wire [31:0]\FRAME_MATCHER.state_c ;   // verilog/coms.v(112[11:16])
    
    wire n10_adj_4133, n8_adj_4134, n44095, n28420, n6_adj_4135, n72, 
        n43481, n9_adj_4136, n43547, n43545, n43543, n43541, n43539, 
        n43537, n43535, n43533, n43531, n43529, n43527, n43525, 
        n43523, n44042, n44113, n43521, n43519, n43975, n43517, 
        n58, n39108, n28421, n28422, n28423, n28424, n28425, n28426, 
        n28427;
    wire [2:0]r_SM_Main_2__N_3516;
    
    wire tx_active, n27687, n4_c, n1, n6_adj_4137;
    wire [0:0]n3912;
    
    wire n44977, n63_c, n63_adj_4138, n8_adj_4141, n28412, n28413;
    wire [7:0]\data_out_frame[18]_c ;   // verilog/coms.v(97[12:26])
    
    wire n28562, \FRAME_MATCHER.rx_data_ready_prev , n5786, n27781, 
        n28414, n39107, n28415, n28416, n28417, n28418, n39106, 
        n28419, n8_adj_4142, n28404, n2_adj_4143, n39105, n2_adj_4144, 
        n39104, n28405, n28406, n2_adj_4145, n39103, n28407, n44947, 
        n28408, n28409, n28410, n2_adj_4146, n39102, n28411, n8_adj_4147, 
        n28396, n2_adj_4148, n39101, n28397, n2_adj_4149, n39100, 
        n28398, n5_adj_4150, n28399, n33752, n26686, n68, n44, 
        n42, n2_adj_4151, n39099, n43, n41, n40_adj_4152, n39_c, 
        n50, n45, n2_adj_4153, n39098, n14_adj_4154, n26689, n15_adj_4155, 
        n26510, n16_adj_4156, n17_adj_4157, n26621, n10_adj_4158, 
        n5809, n10_adj_4159, n14_adj_4160, n5808, n5807, n5806, 
        n5805, n5804, n5803, n5802, n5801, n5800, n26692, n18, 
        n5799, n20_adj_4161, n15_adj_4162, n5798, n5797, n5796, 
        n5795, n16_adj_4163, n5794, n5793, n5792, n17_adj_4164, 
        n2_adj_4165, n39097, n5791, n5790, n5789, n5788, n5787, 
        n20_adj_4166, n19, n48787, n2_adj_4167, n39096, n44079, 
        n2_adj_4168, n39095, n4_adj_4169, n43489, n43587, n2_adj_4170, 
        n39094, n2_adj_4171, n39093, n28400, n28401, n28402, n2_adj_4172, 
        n39092, n2_adj_4173, n39091, n2_adj_4174, n39090, n28403, 
        n8_adj_4175, n28388, n28389, n28390, n28391, n28392, n28393, 
        n28394;
    wire [7:0]\data_in_frame[19] ;   // verilog/coms.v(96[12:25])
    
    wire n5785, n2_adj_4176, n39089, n28395;
    wire [7:0]\data_in_frame[18] ;   // verilog/coms.v(96[12:25])
    
    wire n8_adj_4177, n28380, n2_adj_4178, n39088, n28381, n2_adj_4179, 
        n39087;
    wire [7:0]\data_in_frame[17] ;   // verilog/coms.v(96[12:25])
    
    wire n28382, n2_adj_4180, n39086, n48967, n48968, n49019, n42434, 
        n45731, n49018, n48982, n48983, n48977, n48976, n28383, 
        n28384, n28385, n48985, n48986, n48923, n48922, n48988, 
        n48989, n48887, n48886, n48991, n48992, n2_adj_4181, n39085, 
        n49001, n49000, n49003, n49004, n48857, n48856, n49006, 
        n49007, n7_adj_4183, n43477, n2_adj_4184, n39084, n31_adj_4185, 
        n44979, n69, n46802, n23701, n45946, n2_adj_4186, n39083, 
        n33576, n34368, n43627, n43511, n33574, n34366, n43625, 
        n43513, n33572, n34364, n43623, n43515, n43621, n7_adj_4187, 
        n8_adj_4188, n7_adj_4189, n33570, n43619, n2_adj_4190, n39082, 
        n33568, n34362, n43617, n43615, n43613, n43611, n43609, 
        n43607, n43605, n43603, n43601, n43599, n43597, n43595, 
        n43593, n43591, n43589, n43491, n28386, n14_adj_4191, n2_adj_4192, 
        n39081, n34823, n44989, n12_adj_4193, n67, n28031, n28032, 
        n28387, n48854, n48853, n27172, n2_adj_4194, n39080;
    wire [7:0]\data_out_frame[27] ;   // verilog/coms.v(97[12:26])
    
    wire n45719, n42395, n42381, n41565, n45769;
    wire [7:0]\data_out_frame[26] ;   // verilog/coms.v(97[12:26])
    
    wire n45628, n46698, n46700, n45867, n45555, n45401, n46095, 
        n2_adj_4195, n39079, n2_adj_4196, n39078, n3_adj_4197, n3_adj_4198, 
        n3_adj_4199, n3_adj_4200, n3_adj_4201, n3_adj_4202, n3_adj_4203, 
        n3_adj_4204, n3_adj_4205, n3_adj_4206, n3_adj_4207, n3_adj_4208, 
        n3_adj_4209, n3_adj_4210, n3_adj_4211, n3_adj_4212, n3_adj_4213, 
        n3_adj_4214, n3_adj_4215, n3_adj_4216, n3_adj_4217, n3_adj_4218, 
        n3_adj_4219, n3_adj_4220, n3_adj_4221, n3_adj_4222, n3_adj_4223, 
        n3_adj_4224, n2_adj_4225, n3_adj_4226, n2_adj_4227, n3_adj_4228, 
        n2_adj_4229, n3_adj_4230, n39077, n39076, n50305, n49814, 
        n51627, n51510, n7_adj_4231;
    wire [7:0]tx_data;   // verilog/coms.v(105[13:20])
    
    wire n8_adj_4232;
    wire [7:0]\data_in_frame[14] ;   // verilog/coms.v(96[12:25])
    
    wire n28372, n50303, n49811, n51621, n51504, n7_adj_4233, n50299, 
        n49808, n51615, n48970, n39075, n161, n48971, n49016, 
        n49015, n48914, n48915, n48913, n28373, n51582, n49820, 
        n48884, n51432, n50421, n51498, n7_adj_4234, n28374, n51414, 
        n49805, n51603, n51492, n7_adj_4235, n51420, n49802, n51597, 
        n51486, n7_adj_4236, n51426, n51591, n51480, n7_adj_4237, 
        n50287, n49799, n51585, n51516, n7_adj_4238, n51579, n51573, 
        n51576, n51567, n51570, n51561, n51564, n28375, n51555, 
        n51558, n51549, n51552, n51543, n51537, n51540, n51531, 
        n51474, n7_adj_4239, n51513, n10_adj_4240, n42361, n26249, 
        n42427, n44195, n14_adj_4241, n44694, n34527, n6_adj_4242, 
        n44506, n27497, n41521, n10_adj_4243, n41525, n42363, n26472, 
        n51507, n44_adj_4244, n51501, n42444, n51495, n51489, n44531, 
        n51483, n6_adj_4245, n42333, n33565, n51477, n51471, n26473, 
        n26834, n44055, n42291, n42322, n46232, n44537, n48957, 
        n48955, n44662, n26749, n26890, n44129, n23, n48908, n51456, 
        n44687, n41437, n44381, n48951, n48949;
    wire [7:0]\data_in_frame[15] ;   // verilog/coms.v(96[12:25])
    wire [7:0]\data_in_frame[16] ;   // verilog/coms.v(96[12:25])
    
    wire n44585, n48944, n48945, n48943, n48411, n44754, n48423, 
        n41447, n26854, n27312, n28, n48413, n48938, n44521, Kp_23__N_1402, 
        n48427, n26857, n48433, n44645, n44624, n44324, n48435, 
        n44757, n41445, n44353, n27425, n26, n44766, n22_adj_4246, 
        n44677, n30_adj_4247, n44357, n44668, n48441, n44603, n25, 
        n48379, n44769, n44763, Kp_23__N_1398, n48385, n44680, n44474, 
        n42126, n48391, n44483, n44745, n44656, n48395, n48443, 
        n48939, n48937, n44500, Kp_23__N_1653, n44691, n48399, n45717, 
        n41435, n44715, n48367, n42281, n44230, n42407, n27178, 
        n44390, n42418, Kp_23__N_1644, n44378, Kp_23__N_761, n48523, 
        n28212, n44085, n28322, n42374, n44418, n44712, n28323, 
        n28376, n28321, n41723, n44403, n48653, n28377, n28378, 
        n44549, n46390, n6_adj_4248, n44659, n8_adj_4249, n27347, 
        n27606, n44671, n41580, n44448, n42354, n44652, n44406, 
        n4_adj_4250, n44742, n48559, Kp_23__N_1095, n44527, n46677, 
        n27459, n41956, n41474, n44515, n44458, n27023, n48461, 
        n44503, n42350, Kp_23__N_1221, n27597, n48933, n48931, n44327, 
        n48647, n41494, n42442, n48918, n48916, n44591, n48593, 
        n26978, n44154, n44706, n48599, n44567, n44282, n44639, 
        n48603, n48609, n44512, n42348, n48577, n27587, Kp_23__N_1233, 
        n44718, n48583, n44246, n42367, n6_adj_4251, n44363, n44360, 
        n27650, n44760, n20_adj_4252, n48927, n48925, n44730, n19_adj_4253, 
        n34355, n34549, n34685, n44615, n21, n51453, n41449, n18_adj_4254, 
        n44170, n16_adj_4255, n20_adj_4256, n44553, n44294, n44648, 
        n44739, n27414, n42295, n12_adj_4257, n10_adj_4258, n14_adj_4259, 
        n9_adj_4260, n48477, n26770, n44627, n44736, n27411, n26746, 
        n27010, n48447, n27063, n27584, n44207, n14_adj_4261, n10_adj_4262, 
        n44243, n27360, n48351, n25051, n45701, n44636, n44348, 
        n28379, n25836, Kp_23__N_888, n27198, n44148, n41451, n27297, 
        n44464, n44161, n44642, n10_adj_4263, n44307, n42133, n10_adj_4264, 
        n6_adj_4265, n26866, n44439, n10_adj_4266, n27660, n44674, 
        n10_adj_4267, n44665, n48361, n44251, n41468, n27579, n14_adj_4268, 
        n44454, n44234, n27530, n44556, n26966, n10_adj_4269, n44301, 
        n26996, n44751, n44310, n10_adj_4270, n44339, Kp_23__N_881, 
        n44594, n10_adj_4271, n7_adj_4272, n8_adj_4273, n44345, n44227, 
        n12_adj_4274, Kp_23__N_1647, n44398, n44412, n27465, n41569, 
        n27394, n27058, n44772, Kp_23__N_1114, n28492, n28491, n28490, 
        n28489, n28488, n28485, n28484, n28483, n28482, n28481, 
        n28480, n28479, n28478, n28477, n26938, n28476, n28475, 
        n28474, n28473, n28472, n28471, n28470, n28469, n28468, 
        n28467, n44190, n28466, n28465, n28464, n28463, n28462, 
        n28461, n28460, n28459, n28458, n28457, n28456, n28455, 
        n28454, n28453, Kp_23__N_836, n28452, n28451, n28450, n28449, 
        n28448, n28447, n28446, n28445, n28444, n28443, n28442, 
        n28441, n28440, n28439, n28438, n28437, n28436, n12_adj_4275, 
        n27334, n6_adj_4276, n12_adj_4277, n44709, n8_adj_4278, Kp_23__N_996, 
        n28371, n28370, n28369, n28368, n28367, n28366, n28365, 
        n28364, n28363, Kp_23__N_999, n28362, n28361, n28360, n28359, 
        n28358, n28357, n28356, n28355, n28354, n28353, n28352, 
        n28351, n28350, n28349, n28348, n28347, n28346, n28345, 
        n28344, n28343, n28342, n28341, n28340, n28339, n28338, 
        n28337, n28336, n28335, n28334, n28333, n28332, n28331;
    wire [7:0]\data_in_frame[20] ;   // verilog/coms.v(96[12:25])
    
    wire n28330, n28329, n28328, n28327, n28326, n28325, n28324, 
        n48339, n48341, n48347, n45653, n48355, n45673, n41478, 
        n44395, n31_adj_4279, n48453, n44336, n39112, n44184, n44291, 
        n48617, n39111, n6_adj_4280, n27138, n2206, n11_adj_4281, 
        n6_adj_4282, n6_adj_4283, n24_adj_4284, n12_adj_4285, n45516, 
        n28_adj_4286, n26_adj_4287, n27_adj_4288, n25_adj_4289, n12_adj_4290, 
        n6_adj_4291, n45393, n8_adj_4292, n48487, n48489, n48491, 
        n44159, n45788, n45839, n6_adj_4293, n48497, n48545, n48499, 
        n46067, n46491, n44683, n48505, n44419, n48529, n48535, 
        n46266, n48509, n45684, n45508, n12_adj_4294, n10_adj_4295, 
        n11_adj_4296, n9_adj_4297, n48623, n48629, n51447, n51450, 
        n20_adj_4299, n51441, n34409, n51444, n44570, n19_adj_4300, 
        n46506, n48932, n42170, n21_adj_4301, n48899, n48926, n42438, 
        n48896, n48893, n51438, n51435, n44486, n44494, n41846, 
        n12_adj_4302, n44540, n12_adj_4303, n44237, n13, n42487, 
        n6_adj_4304, n6_adj_4305, n45752, n27163, n44748, n18_adj_4306, 
        n16_adj_4307, n20_adj_4308, n44421, n27244, n46294, n44480, 
        n44433, n30_adj_4309, n34_adj_4310, n32, n33, n31_adj_4311, 
        n45838, n16_adj_4312, n51429, n17_adj_4313, n51423, n17_adj_4314, 
        n49803, n49804, n51417, n17_adj_4316, n16_adj_4317, n49806, 
        n49807, n51411, n17_adj_4318, n16_adj_4319, n13_adj_4320, 
        n44451, n6_adj_4321, n42448, n26_adj_4322, n24_adj_4323, n25_adj_4324, 
        n10_adj_4325, n14_adj_4326, n46282, n44221, n15_adj_4327, 
        n46733, n12_adj_4328, n44564, n42344, n12_adj_4329, n14_adj_4330, 
        n44210, n46, n44_adj_4331, n45_adj_4332, n43_adj_4333, n42_adj_4334, 
        n41_adj_4335, n52, n47, n16_adj_4336, n22_adj_4337, n20_adj_4338, 
        n24_adj_4339, n45357, n7_adj_4340, n16_adj_4341, n17_adj_4342;
    
    SB_LUT4 i15365_3_lut_4_lut (.I0(n34417), .I1(n44104), .I2(rx_data[7]), 
            .I3(\data_in_frame[7] [7]), .O(n28428));
    defparam i15365_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0__i172 (.Q(\data_in_frame[21] [3]), .C(CLK_c), 
           .D(n28320));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i173 (.Q(\data_in_frame[21] [4]), .C(CLK_c), 
           .D(n28319));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i174 (.Q(\data_in_frame[21] [5]), .C(CLK_c), 
           .D(n28318));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i175 (.Q(\data_in_frame[21] [6]), .C(CLK_c), 
           .D(n28317));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[4] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n44218));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i176 (.Q(\data_in_frame[21] [7]), .C(CLK_c), 
           .D(n28316));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut (.I0(n44176), .I1(n27539), .I2(n27558), .I3(n27407), 
            .O(n14));
    defparam i6_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut (.I0(n44321), .I1(n14), .I2(n10_c), .I3(\data_out_frame[8] [6]), 
            .O(n26226));
    defparam i7_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i35729_2_lut (.I0(n27110), .I1(\data_out_frame[13] [4]), .I2(GND_net), 
            .I3(GND_net), .O(n50682));   // verilog/coms.v(97[12:26])
    defparam i35729_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut (.I0(n26226), .I1(n27561), .I2(\data_out_frame[13] [6]), 
            .I3(n50682), .O(n44351));
    defparam i3_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut (.I0(n6), .I1(n44351), .I2(\data_out_frame[18] [3]), 
            .I3(\data_out_frame[16] [2]), .O(n44697));
    defparam i1_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15366_3_lut_4_lut (.I0(n34417), .I1(n44104), .I2(rx_data[6]), 
            .I3(\data_in_frame[7] [6]), .O(n28429));
    defparam i15366_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_852 (.I0(n44333), .I1(n44697), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4111));
    defparam i1_2_lut_adj_852.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut (.I0(\data_out_frame[20] [4]), .I1(n50676), .I2(n44509), 
            .I3(n6_adj_4111), .O(n45876));
    defparam i4_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut (.I0(n45876), .I1(n44518), .I2(n42312), .I3(GND_net), 
            .O(n41225));
    defparam i2_3_lut.LUT_INIT = 16'h6969;
    SB_LUT4 i2_4_lut (.I0(n41225), .I1(\data_out_frame[25] [2]), .I2(n45674), 
            .I3(\data_out_frame[25] [3]), .O(n44489));
    defparam i2_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_853 (.I0(\data_out_frame[11] [4]), .I1(n27212), 
            .I2(n44176), .I3(\data_out_frame[11] [3]), .O(n14_adj_4112));
    defparam i6_4_lut_adj_853.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_854 (.I0(\data_out_frame[13] [5]), .I1(n14_adj_4112), 
            .I2(n10_adj_4113), .I3(n44297), .O(n41601));
    defparam i7_4_lut_adj_854.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_855 (.I0(n41601), .I1(\data_out_frame[11] [5]), 
            .I2(n26380), .I3(GND_net), .O(n45778));
    defparam i2_3_lut_adj_855.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_856 (.I0(\data_out_frame[15] [7]), .I1(n27603), 
            .I2(\data_out_frame[13] [7]), .I3(n45778), .O(n41540));
    defparam i3_4_lut_adj_856.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_857 (.I0(\data_out_frame[16] [1]), .I1(n41540), 
            .I2(GND_net), .I3(GND_net), .O(n41615));
    defparam i1_2_lut_adj_857.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_858 (.I0(\data_out_frame[20] [6]), .I1(n42312), 
            .I2(GND_net), .I3(GND_net), .O(n44509));
    defparam i1_2_lut_adj_858.LUT_INIT = 16'h9999;
    SB_DFFSS \FRAME_MATCHER.i_i0  (.Q(\FRAME_MATCHER.i [0]), .C(CLK_c), 
            .D(n2), .S(n3));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_859 (.I0(n11), .I1(n9), .I2(n44497), .I3(n42416), 
            .O(n42300));
    defparam i6_4_lut_adj_859.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_860 (.I0(\data_out_frame[23] [2]), .I1(\data_out_frame[23] [1]), 
            .I2(n42300), .I3(GND_net), .O(n45674));
    defparam i2_3_lut_adj_860.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_861 (.I0(\data_out_frame[9] [2]), .I1(n44264), 
            .I2(n44151), .I3(\data_out_frame[4] [4]), .O(n27484));   // verilog/coms.v(85[17:70])
    defparam i3_4_lut_adj_861.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_862 (.I0(\data_out_frame[9] [3]), .I1(n27093), 
            .I2(n27666), .I3(n27484), .O(n24830));
    defparam i3_4_lut_adj_862.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_863 (.I0(\data_out_frame[14] [0]), .I1(n44721), 
            .I2(n44597), .I3(n44258), .O(n27603));
    defparam i3_4_lut_adj_863.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_864 (.I0(\data_out_frame[14] [1]), .I1(n27603), 
            .I2(n24830), .I3(\data_out_frame[11] [4]), .O(n6));   // verilog/coms.v(85[17:70])
    defparam i3_4_lut_adj_864.LUT_INIT = 16'h6996;
    SB_LUT4 i911_2_lut (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n1699));   // verilog/coms.v(71[16:27])
    defparam i911_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i35723_2_lut (.I0(n6), .I1(n42493), .I2(GND_net), .I3(GND_net), 
            .O(n50676));
    defparam i35723_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_865 (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[18] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44318));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_865.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_866 (.I0(n41571), .I1(n44497), .I2(\data_out_frame[20] [6]), 
            .I3(n26809), .O(n46253));
    defparam i3_4_lut_adj_866.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_867 (.I0(\data_out_frame[23] [2]), .I1(n46253), 
            .I2(GND_net), .I3(GND_net), .O(n44534));
    defparam i1_2_lut_adj_867.LUT_INIT = 16'h9999;
    SB_LUT4 i15367_3_lut_4_lut (.I0(n34417), .I1(n44104), .I2(rx_data[5]), 
            .I3(\data_in_frame[7] [5]), .O(n28430));
    defparam i15367_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_868 (.I0(\data_out_frame[11] [0]), .I1(\data_out_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44621));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_868.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_869 (.I0(\data_out_frame[11] [3]), .I1(\data_out_frame[11] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44321));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_869.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_870 (.I0(\data_out_frame[7] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(n44612), .I3(n6_adj_4114), .O(n26380));
    defparam i4_4_lut_adj_870.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut (.I0(n26380), .I1(\data_out_frame[11] [4]), .I2(n44268), 
            .I3(GND_net), .O(n14_adj_4115));
    defparam i5_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_871 (.I0(n26755), .I1(n26724), .I2(n44543), .I3(n44703), 
            .O(n15_c));
    defparam i6_4_lut_adj_871.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_872 (.I0(n15_c), .I1(\data_out_frame[12] [3]), 
            .I2(n14_adj_4115), .I3(GND_net), .O(n44700));
    defparam i1_4_lut_adj_872.LUT_INIT = 16'h9696;
    SB_LUT4 i15368_3_lut_4_lut (.I0(n34417), .I1(n44104), .I2(rx_data[4]), 
            .I3(\data_in_frame[7] [4]), .O(n28431));
    defparam i15368_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_873 (.I0(n44321), .I1(n44621), .I2(\data_out_frame[11] [7]), 
            .I3(\data_out_frame[11] [6]), .O(n44703));   // verilog/coms.v(71[16:27])
    defparam i3_4_lut_adj_873.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_874 (.I0(n26281), .I1(\data_out_frame[14] [1]), 
            .I2(\data_out_frame[14] [2]), .I3(GND_net), .O(n44366));
    defparam i2_3_lut_adj_874.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_875 (.I0(n44703), .I1(\data_out_frame[13] [7]), 
            .I2(n44255), .I3(n44700), .O(n15_adj_4116));
    defparam i6_4_lut_adj_875.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut (.I0(n15_adj_4116), .I1(n44471), .I2(n14_adj_4117), 
            .I3(n44201), .O(n42346));
    defparam i8_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_876 (.I0(n42346), .I1(n44366), .I2(\data_out_frame[16] [3]), 
            .I3(GND_net), .O(n42416));
    defparam i2_3_lut_adj_876.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_877 (.I0(n41486), .I1(n41571), .I2(\data_out_frame[16] [5]), 
            .I3(GND_net), .O(n44491));
    defparam i2_3_lut_adj_877.LUT_INIT = 16'h6969;
    SB_LUT4 i4_4_lut_adj_878 (.I0(\data_out_frame[18] [6]), .I1(n42416), 
            .I2(\data_out_frame[18] [5]), .I3(n6_adj_4118), .O(n42312));
    defparam i4_4_lut_adj_878.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_879 (.I0(n42312), .I1(n2122), .I2(\data_out_frame[23] [3]), 
            .I3(GND_net), .O(n46081));
    defparam i2_3_lut_adj_879.LUT_INIT = 16'h6969;
    SB_LUT4 i2_3_lut_adj_880 (.I0(n2122), .I1(n27152), .I2(\data_out_frame[23] [4]), 
            .I3(GND_net), .O(n41597));
    defparam i2_3_lut_adj_880.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_881 (.I0(\data_out_frame[5] [1]), .I1(n44727), 
            .I2(GND_net), .I3(GND_net), .O(n27093));
    defparam i1_2_lut_adj_881.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut (.I0(n44576), .I1(n44600), .I2(\data_out_frame[12] [0]), 
            .I3(n44215), .O(n12));   // verilog/coms.v(71[16:27])
    defparam i5_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_882 (.I0(\data_out_frame[10] [0]), .I1(n12), .I2(n44724), 
            .I3(\data_out_frame[7] [6]), .O(n26281));   // verilog/coms.v(71[16:27])
    defparam i6_4_lut_adj_882.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_883 (.I0(n26281), .I1(\data_out_frame[14] [2]), 
            .I2(n41455), .I3(GND_net), .O(n42493));
    defparam i2_3_lut_adj_883.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_884 (.I0(\data_out_frame[18] [6]), .I1(\data_out_frame[16] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44204));
    defparam i1_2_lut_adj_884.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_885 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[12] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26755));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_885.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_886 (.I0(\data_out_frame[11] [7]), .I1(\data_out_frame[5] [5]), 
            .I2(n44285), .I3(\data_out_frame[9] [5]), .O(n14_adj_4119));
    defparam i6_4_lut_adj_886.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_887 (.I0(n26755), .I1(n14_adj_4119), .I2(n10_adj_4120), 
            .I3(n44609), .O(n44471));
    defparam i7_4_lut_adj_887.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_888 (.I0(n1510), .I1(n44471), .I2(\data_out_frame[14] [3]), 
            .I3(GND_net), .O(n41455));
    defparam i2_3_lut_adj_888.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_889 (.I0(n27321), .I1(\data_out_frame[18] [7]), 
            .I2(\data_out_frame[16] [5]), .I3(GND_net), .O(n44409));
    defparam i2_3_lut_adj_889.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_890 (.I0(\data_out_frame[17] [0]), .I1(\data_out_frame[16] [7]), 
            .I2(n41455), .I3(n6_adj_4121), .O(n41589));
    defparam i4_4_lut_adj_890.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_891 (.I0(\data_out_frame[19] [0]), .I1(n44204), 
            .I2(n42493), .I3(n1794), .O(n10_adj_4122));
    defparam i4_4_lut_adj_891.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_adj_892 (.I0(\data_out_frame[18] [7]), .I1(n10_adj_4122), 
            .I2(\data_out_frame[16] [6]), .I3(GND_net), .O(n41571));
    defparam i5_3_lut_adj_892.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut (.I0(\data_out_frame[25] [5]), .I1(n41597), .I2(n46081), 
            .I3(GND_net), .O(n41553));
    defparam i1_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i15369_3_lut_4_lut (.I0(n34417), .I1(n44104), .I2(rx_data[3]), 
            .I3(\data_in_frame[7] [3]), .O(n28432));
    defparam i15369_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_893 (.I0(\data_out_frame[23] [5]), .I1(\data_out_frame[23] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26846));
    defparam i1_2_lut_adj_893.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_894 (.I0(\data_out_frame[7] [4]), .I1(\data_out_frame[5] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44721));
    defparam i1_2_lut_adj_894.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_895 (.I0(\data_out_frame[9] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(n44285), .I3(n6_adj_4123), .O(n1510));   // verilog/coms.v(74[16:27])
    defparam i4_4_lut_adj_895.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_896 (.I0(n1510), .I1(n44387), .I2(GND_net), .I3(GND_net), 
            .O(n44255));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_896.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_897 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[5] [7]), 
            .I2(\data_out_frame[7] [5]), .I3(n44546), .O(n10_adj_4124));   // verilog/coms.v(75[16:27])
    defparam i4_4_lut_adj_897.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_898 (.I0(n44304), .I1(\data_out_frame[12] [3]), 
            .I2(\data_out_frame[9] [7]), .I3(GND_net), .O(n44387));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_898.LUT_INIT = 16'h9696;
    SB_LUT4 i15370_3_lut_4_lut (.I0(n34417), .I1(n44104), .I2(rx_data[2]), 
            .I3(\data_in_frame[7] [2]), .O(n28433));
    defparam i15370_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_899 (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[4] [2]), 
            .I2(\data_out_frame[10] [4]), .I3(n27288), .O(n14_adj_4125));   // verilog/coms.v(73[16:42])
    defparam i6_4_lut_adj_899.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_900 (.I0(n1519), .I1(n14_adj_4125), .I2(n10_adj_4126), 
            .I3(n44198), .O(n44268));   // verilog/coms.v(73[16:42])
    defparam i7_4_lut_adj_900.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_901 (.I0(\data_out_frame[12] [6]), .I1(n44268), 
            .I2(\data_out_frame[12] [5]), .I3(\data_out_frame[14] [7]), 
            .O(n41480));
    defparam i3_4_lut_adj_901.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_902 (.I0(\data_out_frame[14] [5]), .I1(n44387), 
            .I2(n1516), .I3(\data_out_frame[12] [4]), .O(n27220));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_902.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_903 (.I0(n27220), .I1(n41480), .I2(\data_out_frame[15] [0]), 
            .I3(GND_net), .O(n44477));
    defparam i2_3_lut_adj_903.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_904 (.I0(\data_out_frame[9] [4]), .I1(\data_out_frame[9] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n44724));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_904.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_905 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[5] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44215));   // verilog/coms.v(71[16:62])
    defparam i1_2_lut_adj_905.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_906 (.I0(\data_out_frame[5] [0]), .I1(n1168), .I2(GND_net), 
            .I3(GND_net), .O(n44264));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_906.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_907 (.I0(\data_out_frame[6] [7]), .I1(\data_out_frame[6] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44151));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_907.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_908 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44198));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_908.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_909 (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[4] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44384));
    defparam i1_2_lut_adj_909.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_910 (.I0(\data_out_frame[7] [6]), .I1(\data_out_frame[7] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44609));
    defparam i1_2_lut_adj_910.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_911 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[8] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44579));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_911.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_912 (.I0(\data_out_frame[5] [0]), .I1(\data_out_frame[7] [2]), 
            .I2(\data_out_frame[4] [6]), .I3(GND_net), .O(n44727));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_912.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_913 (.I0(n27666), .I1(\data_out_frame[7] [1]), 
            .I2(\data_out_frame[8] [7]), .I3(GND_net), .O(n44176));   // verilog/coms.v(75[16:27])
    defparam i2_3_lut_adj_913.LUT_INIT = 16'h9696;
    SB_LUT4 i3_2_lut (.I0(n44176), .I1(\data_out_frame[8] [2]), .I2(GND_net), 
            .I3(GND_net), .O(n24));
    defparam i3_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i13_4_lut (.I0(n44727), .I1(n44559), .I2(n44579), .I3(\data_out_frame[4] [6]), 
            .O(n34));
    defparam i13_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_914 (.I0(n44573), .I1(\data_out_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n22));
    defparam i1_2_lut_adj_914.LUT_INIT = 16'h6666;
    SB_LUT4 i17_4_lut (.I0(\data_out_frame[8] [5]), .I1(n34), .I2(n24), 
            .I3(n44609), .O(n38));
    defparam i17_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut (.I0(\data_out_frame[5] [5]), .I1(n44384), .I2(n26712), 
            .I3(n44198), .O(n36));
    defparam i15_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[6] [0]), 
            .I2(\data_out_frame[4] [7]), .I3(n22), .O(n37));
    defparam i16_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut (.I0(\data_out_frame[7] [4]), .I1(n44330), .I2(\data_out_frame[8] [0]), 
            .I3(n27558), .O(n35));
    defparam i14_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut (.I0(n35), .I1(n37), .I2(n36), .I3(n38), .O(n42075));
    defparam i20_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_915 (.I0(\data_out_frame[9] [7]), .I1(\data_out_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44600));
    defparam i1_2_lut_adj_915.LUT_INIT = 16'h6666;
    SB_DFFESR byte_transmit_counter_i0_i1 (.Q(byte_transmit_counter[1]), .C(CLK_c), 
            .E(n27787), .D(n8825[1]), .R(n33303));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_916 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[4] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44330));
    defparam i1_2_lut_adj_916.LUT_INIT = 16'h6666;
    SB_DFFESR byte_transmit_counter_i0_i2 (.Q(\byte_transmit_counter[2] ), 
            .C(CLK_c), .E(n27787), .D(n8825[2]), .R(n33303));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_917 (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[10] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27269));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_917.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_918 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n44342));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_918.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_919 (.I0(n27403), .I1(n44342), .I2(n27269), .I3(n44630), 
            .O(n12_adj_4127));   // verilog/coms.v(85[17:63])
    defparam i5_4_lut_adj_919.LUT_INIT = 16'h6996;
    SB_DFFESR byte_transmit_counter_i0_i3 (.Q(byte_transmit_counter[3]), .C(CLK_c), 
            .E(n27787), .D(n8825[3]), .R(n33303));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i4 (.Q(byte_transmit_counter[4]), .C(CLK_c), 
            .E(n27787), .D(n8825[4]), .R(n33303));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i5 (.Q(byte_transmit_counter[5]), .C(CLK_c), 
            .E(n27787), .D(n8825[5]), .R(n33303));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i6 (.Q(byte_transmit_counter[6]), .C(CLK_c), 
            .E(n27787), .D(n8825[6]), .R(n33303));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i7 (.Q(byte_transmit_counter[7]), .C(CLK_c), 
            .E(n27787), .D(n8825[7]), .R(n33303));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_920 (.I0(\data_out_frame[10] [6]), .I1(n12_adj_4127), 
            .I2(\data_out_frame[10] [0]), .I3(n42387), .O(n44136));   // verilog/coms.v(85[17:63])
    defparam i6_4_lut_adj_920.LUT_INIT = 16'h9669;
    SB_LUT4 i15371_3_lut_4_lut (.I0(n34417), .I1(n44104), .I2(rx_data[1]), 
            .I3(\data_in_frame[7] [1]), .O(n28434));
    defparam i15371_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i6_4_lut_adj_921 (.I0(\data_out_frame[9] [0]), .I1(\data_out_frame[9] [2]), 
            .I2(n44258), .I3(\data_out_frame[9] [1]), .O(n16));
    defparam i6_4_lut_adj_921.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_922 (.I0(\data_out_frame[9] [3]), .I1(\data_out_frame[5] [4]), 
            .I2(n44600), .I3(n42075), .O(n17));
    defparam i7_4_lut_adj_922.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut (.I0(n17), .I1(\data_out_frame[7] [5]), .I2(n16), 
            .I3(n27403), .O(n42387));
    defparam i9_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_923 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[8] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44546));   // verilog/coms.v(72[16:27])
    defparam i1_2_lut_adj_923.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_924 (.I0(\data_out_frame[6] [1]), .I1(\data_out_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n44224));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_924.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_925 (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44630));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_925.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_926 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44139));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_926.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_927 (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n44559));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_adj_927.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_928 (.I0(\data_out_frame[5] [4]), .I1(n44606), 
            .I2(n44582), .I3(n44224), .O(n1516));   // verilog/coms.v(85[17:70])
    defparam i3_4_lut_adj_928.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_929 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n26724));   // verilog/coms.v(85[17:63])
    defparam i1_2_lut_adj_929.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_930 (.I0(n44559), .I1(n44139), .I2(\data_out_frame[6] [1]), 
            .I3(n44630), .O(n10_adj_4128));   // verilog/coms.v(72[16:27])
    defparam i4_4_lut_adj_930.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_931 (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[10] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n27288));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_931.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_932 (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44461));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_932.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_933 (.I0(n44524), .I1(n44582), .I2(\data_out_frame[10] [1]), 
            .I3(n26712), .O(n15_adj_4129));
    defparam i6_4_lut_adj_933.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_934 (.I0(n15_adj_4129), .I1(n42387), .I2(n14_adj_4130), 
            .I3(n44136), .O(n42285));
    defparam i8_4_lut_adj_934.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_935 (.I0(n42285), .I1(\data_out_frame[13] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n42365));
    defparam i1_2_lut_adj_935.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_936 (.I0(n1519), .I1(n44201), .I2(\data_out_frame[14] [6]), 
            .I3(GND_net), .O(n27321));
    defparam i2_3_lut_adj_936.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_937 (.I0(\data_out_frame[15] [0]), .I1(\data_out_frame[15] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44424));
    defparam i1_2_lut_adj_937.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_938 (.I0(\data_out_frame[17] [2]), .I1(n44424), 
            .I2(n27321), .I3(n42365), .O(n42378));
    defparam i3_4_lut_adj_938.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_939 (.I0(n44477), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [7]), .I3(GND_net), .O(n44445));
    defparam i2_3_lut_adj_939.LUT_INIT = 16'h9696;
    SB_LUT4 i15372_3_lut_4_lut (.I0(n34417), .I1(n44104), .I2(rx_data[0]), 
            .I3(\data_in_frame[7] [0]), .O(n28435));
    defparam i15372_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_3_lut (.I0(n27321), .I1(\data_out_frame[17] [0]), .I2(n44688), 
            .I3(GND_net), .O(n8));
    defparam i3_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_940 (.I0(\data_out_frame[19] [2]), .I1(\data_out_frame[16] [6]), 
            .I2(n8), .I3(n44477), .O(n42393));
    defparam i1_4_lut_adj_940.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_941 (.I0(n26846), .I1(n41553), .I2(n2122), .I3(\data_out_frame[25] [6]), 
            .O(n44427));
    defparam i3_4_lut_adj_941.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_942 (.I0(n42393), .I1(n44445), .I2(n42378), .I3(\data_out_frame[19] [3]), 
            .O(n42339));
    defparam i3_4_lut_adj_942.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_943 (.I0(n34047), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n44929), .I3(GND_net), .O(n27912));
    defparam i3_3_lut_adj_943.LUT_INIT = 16'h0404;
    SB_LUT4 i1_2_lut_adj_944 (.I0(n42339), .I1(n44427), .I2(GND_net), 
            .I3(GND_net), .O(n44428));
    defparam i1_2_lut_adj_944.LUT_INIT = 16'h9999;
    SB_CARRY add_3971_6 (.CI(n39109), .I0(byte_transmit_counter[4]), .I1(GND_net), 
            .CO(n39110));
    SB_LUT4 i1_2_lut_adj_945 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[0] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n44373));   // verilog/coms.v(77[16:27])
    defparam i1_2_lut_adj_945.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_946 (.I0(\data_in_frame[0] [7]), .I1(n44373), .I2(n44261), 
            .I3(n44142), .O(Kp_23__N_869));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_946.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_947 (.I0(\data_in_frame[0] [0]), .I1(Kp_23__N_869), 
            .I2(GND_net), .I3(GND_net), .O(n44271));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_adj_947.LUT_INIT = 16'h6666;
    SB_LUT4 i33897_4_lut (.I0(\data_in_frame[2] [0]), .I1(n27356), .I2(n44271), 
            .I3(n7_c), .O(n48791));
    defparam i33897_4_lut.LUT_INIT = 16'hffde;
    SB_LUT4 i3_2_lut_adj_948 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[1] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n20));
    defparam i3_2_lut_adj_948.LUT_INIT = 16'h8888;
    SB_LUT4 i10_4_lut (.I0(\data_in_frame[1] [7]), .I1(n20), .I2(\data_in_frame[1] [3]), 
            .I3(n44271), .O(n27));
    defparam i10_4_lut.LUT_INIT = 16'h4080;
    SB_LUT4 i7_4_lut_adj_949 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[1] [1]), 
            .I2(n44373), .I3(\data_in_frame[0] [7]), .O(n24_adj_4131));
    defparam i7_4_lut_adj_949.LUT_INIT = 16'h8421;
    SB_LUT4 i13_4_lut_adj_950 (.I0(Kp_23__N_869), .I1(n48791), .I2(n27337), 
            .I3(\data_in_frame[2] [1]), .O(n30));
    defparam i13_4_lut_adj_950.LUT_INIT = 16'h0102;
    SB_LUT4 i14_4_lut_adj_951 (.I0(n27), .I1(n24120), .I2(n22_adj_4132), 
            .I3(\data_in_frame[1] [4]), .O(n31));
    defparam i14_4_lut_adj_951.LUT_INIT = 16'h2000;
    SB_LUT4 i16_4_lut_adj_952 (.I0(n31), .I1(n48673), .I2(n30), .I3(n24_adj_4131), 
            .O(\FRAME_MATCHER.state_31__N_2624 [3]));
    defparam i16_4_lut_adj_952.LUT_INIT = 16'h2000;
    SB_LUT4 i84_4_lut (.I0(n33307), .I1(n81), .I2(\FRAME_MATCHER.state_31__N_2624 [3]), 
            .I3(\FRAME_MATCHER.state_c [2]), .O(n10_adj_4133));
    defparam i84_4_lut.LUT_INIT = 16'hccdc;
    SB_LUT4 i15357_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44095), .I2(rx_data[7]), 
            .I3(\data_in_frame[8] [7]), .O(n28420));
    defparam i15357_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_adj_953 (.I0(\FRAME_MATCHER.state [3]), .I1(n6_adj_4135), 
            .I2(n72), .I3(GND_net), .O(n43481));
    defparam i1_3_lut_adj_953.LUT_INIT = 16'ha8a8;
    SB_LUT4 i1_2_lut_adj_954 (.I0(\FRAME_MATCHER.state_c [5]), .I1(n9_adj_4136), 
            .I2(GND_net), .I3(GND_net), .O(n43547));
    defparam i1_2_lut_adj_954.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_955 (.I0(\FRAME_MATCHER.state_c [6]), .I1(n9_adj_4136), 
            .I2(GND_net), .I3(GND_net), .O(n43545));
    defparam i1_2_lut_adj_955.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_956 (.I0(\FRAME_MATCHER.state_c [7]), .I1(n9_adj_4136), 
            .I2(GND_net), .I3(GND_net), .O(n43543));
    defparam i1_2_lut_adj_956.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_957 (.I0(\FRAME_MATCHER.state_c [8]), .I1(n9_adj_4136), 
            .I2(GND_net), .I3(GND_net), .O(n43541));
    defparam i1_2_lut_adj_957.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_958 (.I0(\FRAME_MATCHER.state_c [9]), .I1(n9_adj_4136), 
            .I2(GND_net), .I3(GND_net), .O(n43539));
    defparam i1_2_lut_adj_958.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_959 (.I0(\FRAME_MATCHER.state_c [10]), .I1(n9_adj_4136), 
            .I2(GND_net), .I3(GND_net), .O(n43537));
    defparam i1_2_lut_adj_959.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_960 (.I0(\FRAME_MATCHER.state_c [11]), .I1(n9_adj_4136), 
            .I2(GND_net), .I3(GND_net), .O(n43535));
    defparam i1_2_lut_adj_960.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_961 (.I0(\FRAME_MATCHER.state_c [12]), .I1(n9_adj_4136), 
            .I2(GND_net), .I3(GND_net), .O(n43533));
    defparam i1_2_lut_adj_961.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_962 (.I0(\FRAME_MATCHER.state_c [13]), .I1(n9_adj_4136), 
            .I2(GND_net), .I3(GND_net), .O(n43531));
    defparam i1_2_lut_adj_962.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_963 (.I0(\FRAME_MATCHER.state_c [14]), .I1(n9_adj_4136), 
            .I2(GND_net), .I3(GND_net), .O(n43529));
    defparam i1_2_lut_adj_963.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_964 (.I0(\FRAME_MATCHER.state_c [15]), .I1(n9_adj_4136), 
            .I2(GND_net), .I3(GND_net), .O(n43527));
    defparam i1_2_lut_adj_964.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_965 (.I0(\FRAME_MATCHER.state_c [16]), .I1(n9_adj_4136), 
            .I2(GND_net), .I3(GND_net), .O(n43525));
    defparam i1_2_lut_adj_965.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_966 (.I0(\FRAME_MATCHER.state_c [17]), .I1(n9_adj_4136), 
            .I2(GND_net), .I3(GND_net), .O(n43523));
    defparam i1_2_lut_adj_966.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_967 (.I0(\FRAME_MATCHER.state_c [18]), .I1(n44042), 
            .I2(n44113), .I3(n44058), .O(n43521));
    defparam i1_4_lut_adj_967.LUT_INIT = 16'ha8a0;
    SB_LUT4 i1_2_lut_adj_968 (.I0(\FRAME_MATCHER.state_c [20]), .I1(n9_adj_4136), 
            .I2(GND_net), .I3(GND_net), .O(n43519));
    defparam i1_2_lut_adj_968.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_969 (.I0(n33307), .I1(n44113), .I2(n33302), .I3(n43975), 
            .O(n9_adj_4136));
    defparam i1_4_lut_adj_969.LUT_INIT = 16'heccc;
    SB_LUT4 i1_2_lut_adj_970 (.I0(\FRAME_MATCHER.state_c [23]), .I1(n9_adj_4136), 
            .I2(GND_net), .I3(GND_net), .O(n43517));
    defparam i1_2_lut_adj_970.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_adj_971 (.I0(n23831), .I1(n46759), .I2(GND_net), 
            .I3(GND_net), .O(n58));
    defparam i1_2_lut_adj_971.LUT_INIT = 16'h2222;
    SB_LUT4 add_3971_5_lut (.I0(GND_net), .I1(byte_transmit_counter[3]), 
            .I2(GND_net), .I3(n39108), .O(n8825[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15358_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44095), .I2(rx_data[6]), 
            .I3(\data_in_frame[8] [6]), .O(n28421));
    defparam i15358_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15359_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44095), .I2(rx_data[5]), 
            .I3(\data_in_frame[8] [5]), .O(n28422));
    defparam i15359_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15360_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44095), .I2(rx_data[4]), 
            .I3(\data_in_frame[8] [4]), .O(n28423));
    defparam i15360_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15361_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44095), .I2(rx_data[3]), 
            .I3(\data_in_frame[8] [3]), .O(n28424));
    defparam i15361_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15362_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44095), .I2(rx_data[2]), 
            .I3(\data_in_frame[8] [2]), .O(n28425));
    defparam i15362_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15363_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44095), .I2(rx_data[1]), 
            .I3(\data_in_frame[8] [1]), .O(n28426));
    defparam i15363_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15364_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44095), .I2(rx_data[0]), 
            .I3(\data_in_frame[8] [0]), .O(n28427));
    defparam i15364_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_972 (.I0(r_SM_Main_2__N_3516[0]), .I1(tx_active), 
            .I2(GND_net), .I3(GND_net), .O(n40));
    defparam i1_2_lut_adj_972.LUT_INIT = 16'heeee;
    SB_LUT4 i2_3_lut_4_lut (.I0(n26712), .I1(\data_out_frame[6] [1]), .I2(\data_out_frame[4] [0]), 
            .I3(\data_out_frame[5] [7]), .O(n27687));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_973 (.I0(n4_c), .I1(n1), .I2(GND_net), .I3(GND_net), 
            .O(n44113));
    defparam i1_2_lut_adj_973.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_974 (.I0(n43975), .I1(n33308), .I2(n5728), .I3(n44035), 
            .O(n6_adj_4135));
    defparam i2_4_lut_adj_974.LUT_INIT = 16'h88a8;
    SB_LUT4 i1_2_lut_adj_975 (.I0(n61), .I1(n76), .I2(GND_net), .I3(GND_net), 
            .O(n6_adj_4137));
    defparam i1_2_lut_adj_975.LUT_INIT = 16'hbbbb;
    SB_DFFSR tx_transmit_3871 (.Q(r_SM_Main_2__N_3516[0]), .C(CLK_c), .D(n3912[0]), 
            .R(n44977));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_976 (.I0(n2482), .I1(n33307), .I2(n33302), .I3(n6_adj_4137), 
            .O(n46759));
    defparam i4_4_lut_adj_976.LUT_INIT = 16'hffbf;
    SB_LUT4 i1_3_lut_adj_977 (.I0(\FRAME_MATCHER.state_c [2]), .I1(n63_c), 
            .I2(n63_adj_4138), .I3(GND_net), .O(n29985));   // verilog/coms.v(112[11:16])
    defparam i1_3_lut_adj_977.LUT_INIT = 16'hb3b3;
    SB_LUT4 i1_rep_231_2_lut (.I0(n63), .I1(n29985), .I2(GND_net), .I3(GND_net), 
            .O(n51904));   // verilog/coms.v(112[11:16])
    defparam i1_rep_231_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 select_455_Select_2_i5_4_lut (.I0(n63), .I1(\FRAME_MATCHER.i_31__N_2524 ), 
            .I2(n3303), .I3(n29985), .O(n5));
    defparam select_455_Select_2_i5_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 select_455_Select_2_i7_4_lut (.I0(n63), .I1(\FRAME_MATCHER.i_31__N_2526 ), 
            .I2(n4452), .I3(n29985), .O(n7));
    defparam select_455_Select_2_i7_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 i15349_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44095), .I2(rx_data[7]), 
            .I3(\data_in_frame[9] [7]), .O(n28412));
    defparam i15349_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15350_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44095), .I2(rx_data[6]), 
            .I3(\data_in_frame[9] [6]), .O(n28413));
    defparam i15350_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut (.I0(n1168), .I1(\data_out_frame[4] [7]), .I2(\data_out_frame[9] [3]), 
            .I3(GND_net), .O(n44297));   // verilog/coms.v(71[16:69])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i17138_3_lut (.I0(\data_out_frame[18]_c [1]), .I1(\displacement[17] ), 
            .I2(n23935), .I3(GND_net), .O(n28562));
    defparam i17138_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_3971_5 (.CI(n39108), .I0(byte_transmit_counter[3]), .I1(GND_net), 
            .CO(n39109));
    SB_DFF \FRAME_MATCHER.rx_data_ready_prev_3872  (.Q(\FRAME_MATCHER.rx_data_ready_prev ), 
           .C(CLK_c), .D(rx_data_ready));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_978 (.I0(\FRAME_MATCHER.state [3]), .I1(n33298), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(n73), .O(n76));
    defparam i3_4_lut_adj_978.LUT_INIT = 16'hfdff;
    SB_DFFE setpoint__i0 (.Q(setpoint[0]), .C(CLK_c), .E(n27781), .D(n5786));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15351_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44095), .I2(rx_data[5]), 
            .I3(\data_in_frame[9] [5]), .O(n28414));
    defparam i15351_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_3971_4_lut (.I0(GND_net), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(n39107), .O(n8825[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_4_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15352_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44095), .I2(rx_data[4]), 
            .I3(\data_in_frame[9] [4]), .O(n28415));
    defparam i15352_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15353_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44095), .I2(rx_data[3]), 
            .I3(\data_in_frame[9] [3]), .O(n28416));
    defparam i15353_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15354_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44095), .I2(rx_data[2]), 
            .I3(\data_in_frame[9] [2]), .O(n28417));
    defparam i15354_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15355_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44095), .I2(rx_data[1]), 
            .I3(\data_in_frame[9] [1]), .O(n28418));
    defparam i15355_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_979 (.I0(n33302), .I1(n76), .I2(GND_net), .I3(GND_net), 
            .O(n33303));
    defparam i1_2_lut_adj_979.LUT_INIT = 16'h2222;
    SB_LUT4 i2_2_lut_3_lut (.I0(n1168), .I1(\data_out_frame[4] [7]), .I2(n27484), 
            .I3(GND_net), .O(n10_c));   // verilog/coms.v(71[16:69])
    defparam i2_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_CARRY add_3971_4 (.CI(n39107), .I0(\byte_transmit_counter[2] ), .I1(GND_net), 
            .CO(n39108));
    SB_LUT4 add_3971_3_lut (.I0(GND_net), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(n39106), .O(n8825[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_3 (.CI(n39106), .I0(byte_transmit_counter[1]), .I1(GND_net), 
            .CO(n39107));
    SB_LUT4 add_3971_2_lut (.I0(GND_net), .I1(\byte_transmit_counter[0] ), 
            .I2(tx_transmit_N_3413), .I3(GND_net), .O(n8825[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15356_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44095), .I2(rx_data[0]), 
            .I3(\data_in_frame[9] [0]), .O(n28419));
    defparam i15356_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15341_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44095), .I2(rx_data[7]), 
            .I3(\data_in_frame[10] [7]), .O(n28404));
    defparam i15341_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_3971_2 (.CI(GND_net), .I0(\byte_transmit_counter[0] ), 
            .I1(tx_transmit_N_3413), .CO(n39106));
    SB_LUT4 add_43_33_lut (.I0(n2482), .I1(\FRAME_MATCHER.i[31] ), .I2(GND_net), 
            .I3(n39105), .O(n2_adj_4143)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_33_lut.LUT_INIT = 16'h8228;
    SB_LUT4 add_43_32_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [30]), .I2(GND_net), 
            .I3(n39104), .O(n2_adj_4144)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_32_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15342_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44095), .I2(rx_data[6]), 
            .I3(\data_in_frame[10] [6]), .O(n28405));
    defparam i15342_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15343_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44095), .I2(rx_data[5]), 
            .I3(\data_in_frame[10] [5]), .O(n28406));
    defparam i15343_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_32 (.CI(n39104), .I0(\FRAME_MATCHER.i [30]), .I1(GND_net), 
            .CO(n39105));
    SB_LUT4 add_43_31_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [29]), .I2(GND_net), 
            .I3(n39103), .O(n2_adj_4145)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_31_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15344_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44095), .I2(rx_data[4]), 
            .I3(\data_in_frame[10] [4]), .O(n28407));
    defparam i15344_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_980 (.I0(n44947), .I1(\FRAME_MATCHER.state [3]), 
            .I2(\FRAME_MATCHER.state_c [1]), .I3(\FRAME_MATCHER.state_31__N_2624 [3]), 
            .O(n23935));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_980.LUT_INIT = 16'h1000;
    SB_LUT4 i15345_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44095), .I2(rx_data[3]), 
            .I3(\data_in_frame[10] [3]), .O(n28408));
    defparam i15345_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15346_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44095), .I2(rx_data[2]), 
            .I3(\data_in_frame[10] [2]), .O(n28409));
    defparam i15346_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15347_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44095), .I2(rx_data[1]), 
            .I3(\data_in_frame[10] [1]), .O(n28410));
    defparam i15347_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_31 (.CI(n39103), .I0(\FRAME_MATCHER.i [29]), .I1(GND_net), 
            .CO(n39104));
    SB_LUT4 add_43_30_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [28]), .I2(GND_net), 
            .I3(n39102), .O(n2_adj_4146)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_30_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15348_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44095), .I2(rx_data[0]), 
            .I3(\data_in_frame[10] [0]), .O(n28411));
    defparam i15348_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15333_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44095), .I2(rx_data[7]), 
            .I3(\data_in_frame[11] [7]), .O(n28396));
    defparam i15333_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF control_mode_i0_i1 (.Q(control_mode[1]), .C(CLK_c), .D(n28284));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i2 (.Q(control_mode[2]), .C(CLK_c), .D(n28283));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i3 (.Q(control_mode[3]), .C(CLK_c), .D(n28282));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i4 (.Q(control_mode[4]), .C(CLK_c), .D(n28281));   // verilog/coms.v(127[12] 300[6])
    SB_DFF control_mode_i0_i5 (.Q(control_mode[5]), .C(CLK_c), .D(n28280));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_30 (.CI(n39102), .I0(\FRAME_MATCHER.i [28]), .I1(GND_net), 
            .CO(n39103));
    SB_LUT4 add_43_29_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [27]), .I2(GND_net), 
            .I3(n39101), .O(n2_adj_4148)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_29_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_29 (.CI(n39101), .I0(\FRAME_MATCHER.i [27]), .I1(GND_net), 
            .CO(n39102));
    SB_LUT4 i15334_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44095), .I2(rx_data[6]), 
            .I3(\data_in_frame[11] [6]), .O(n28397));
    defparam i15334_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF control_mode_i0_i6 (.Q(control_mode[6]), .C(CLK_c), .D(n28279));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_28_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [26]), .I2(GND_net), 
            .I3(n39100), .O(n2_adj_4149)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_28_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i15335_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44095), .I2(rx_data[5]), 
            .I3(\data_in_frame[11] [5]), .O(n28398));
    defparam i15335_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i20819_4_lut (.I0(n5_adj_4150), .I1(\FRAME_MATCHER.i[31] ), 
            .I2(\FRAME_MATCHER.i [3]), .I3(\FRAME_MATCHER.i [2]), .O(n771));   // verilog/coms.v(157[9:60])
    defparam i20819_4_lut.LUT_INIT = 16'h3332;
    SB_LUT4 i15336_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44095), .I2(rx_data[4]), 
            .I3(\data_in_frame[11] [4]), .O(n28399));
    defparam i15336_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i20702_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(GND_net), .I3(GND_net), .O(n33752));
    defparam i20702_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut_adj_981 (.I0(n33752), .I1(n26686), .I2(\FRAME_MATCHER.i [4]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n26687));
    defparam i1_4_lut_adj_981.LUT_INIT = 16'hfcec;
    SB_LUT4 i20822_2_lut (.I0(n26687), .I1(\FRAME_MATCHER.i[31] ), .I2(GND_net), 
            .I3(GND_net), .O(n4452));   // verilog/coms.v(259[9:58])
    defparam i20822_2_lut.LUT_INIT = 16'h2222;
    SB_CARRY add_43_28 (.CI(n39100), .I0(\FRAME_MATCHER.i [26]), .I1(GND_net), 
            .CO(n39101));
    SB_LUT4 i104_3_lut (.I0(n33302), .I1(n1476), .I2(n23831), .I3(GND_net), 
            .O(n68));   // verilog/coms.v(115[11:12])
    defparam i104_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i18_4_lut (.I0(\FRAME_MATCHER.i [30]), .I1(\FRAME_MATCHER.i [21]), 
            .I2(\FRAME_MATCHER.i [24]), .I3(\FRAME_MATCHER.i [17]), .O(n44));
    defparam i18_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i16_4_lut_adj_982 (.I0(\FRAME_MATCHER.i [29]), .I1(\FRAME_MATCHER.i [6]), 
            .I2(\FRAME_MATCHER.i [18]), .I3(\FRAME_MATCHER.i [23]), .O(n42));
    defparam i16_4_lut_adj_982.LUT_INIT = 16'hfffe;
    SB_LUT4 add_43_27_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [25]), .I2(GND_net), 
            .I3(n39099), .O(n2_adj_4151)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_27_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i17_4_lut_adj_983 (.I0(\FRAME_MATCHER.i [7]), .I1(\FRAME_MATCHER.i [20]), 
            .I2(\FRAME_MATCHER.i [12]), .I3(\FRAME_MATCHER.i [14]), .O(n43));
    defparam i17_4_lut_adj_983.LUT_INIT = 16'hfffe;
    SB_DFF control_mode_i0_i7 (.Q(control_mode[7]), .C(CLK_c), .D(n28278));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i1 (.Q(PWMLimit[1]), .C(CLK_c), .D(n28277));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i2 (.Q(PWMLimit[2]), .C(CLK_c), .D(n28276));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i3 (.Q(PWMLimit[3]), .C(CLK_c), .D(n28275));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i4 (.Q(PWMLimit[4]), .C(CLK_c), .D(n28274));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i5 (.Q(PWMLimit[5]), .C(CLK_c), .D(n28273));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15_4_lut_adj_984 (.I0(\FRAME_MATCHER.i [22]), .I1(\FRAME_MATCHER.i [11]), 
            .I2(\FRAME_MATCHER.i [26]), .I3(\FRAME_MATCHER.i [16]), .O(n41));
    defparam i15_4_lut_adj_984.LUT_INIT = 16'hfffe;
    SB_LUT4 i14_4_lut_adj_985 (.I0(\FRAME_MATCHER.i [13]), .I1(\FRAME_MATCHER.i [15]), 
            .I2(\FRAME_MATCHER.i [10]), .I3(\FRAME_MATCHER.i [28]), .O(n40_adj_4152));
    defparam i14_4_lut_adj_985.LUT_INIT = 16'hfffe;
    SB_LUT4 i13_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(\FRAME_MATCHER.i [27]), 
            .I2(GND_net), .I3(GND_net), .O(n39_c));
    defparam i13_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i24_4_lut (.I0(n41), .I1(n43), .I2(n42), .I3(n44), .O(n50));
    defparam i24_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i19_4_lut (.I0(\FRAME_MATCHER.i [8]), .I1(\FRAME_MATCHER.i [25]), 
            .I2(\FRAME_MATCHER.i [5]), .I3(\FRAME_MATCHER.i [19]), .O(n45));
    defparam i19_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY add_43_27 (.CI(n39099), .I0(\FRAME_MATCHER.i [25]), .I1(GND_net), 
            .CO(n39100));
    SB_LUT4 i25_4_lut (.I0(n45), .I1(n50), .I2(n39_c), .I3(n40_adj_4152), 
            .O(n26686));
    defparam i25_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 add_43_26_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [24]), .I2(GND_net), 
            .I3(n39098), .O(n2_adj_4153)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_26_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_26 (.CI(n39098), .I0(\FRAME_MATCHER.i [24]), .I1(GND_net), 
            .CO(n39099));
    SB_LUT4 i20821_2_lut (.I0(n26489), .I1(\FRAME_MATCHER.i[31] ), .I2(GND_net), 
            .I3(GND_net), .O(n3303));   // verilog/coms.v(227[9:54])
    defparam i20821_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i5_3_lut_adj_986 (.I0(\data_in[3] [0]), .I1(\data_in[1] [4]), 
            .I2(\data_in[1] [5]), .I3(GND_net), .O(n14_adj_4154));
    defparam i5_3_lut_adj_986.LUT_INIT = 16'hdfdf;
    SB_LUT4 i6_4_lut_adj_987 (.I0(\data_in[0] [6]), .I1(n26689), .I2(\data_in[2] [4]), 
            .I3(\data_in[1] [0]), .O(n15_adj_4155));
    defparam i6_4_lut_adj_987.LUT_INIT = 16'hfeff;
    SB_LUT4 i8_4_lut_adj_988 (.I0(n15_adj_4155), .I1(\data_in[2] [2]), .I2(n14_adj_4154), 
            .I3(\data_in[0] [3]), .O(n26510));
    defparam i8_4_lut_adj_988.LUT_INIT = 16'hfbff;
    SB_LUT4 i6_4_lut_adj_989 (.I0(\data_in[1] [3]), .I1(\data_in[0] [1]), 
            .I2(\data_in[3] [2]), .I3(\data_in[0] [5]), .O(n16_adj_4156));
    defparam i6_4_lut_adj_989.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_4_lut_adj_990 (.I0(\data_in[2] [6]), .I1(\data_in[2] [5]), 
            .I2(\data_in[2] [0]), .I3(\data_in[1] [2]), .O(n17_adj_4157));
    defparam i7_4_lut_adj_990.LUT_INIT = 16'hfffd;
    SB_LUT4 i9_4_lut_adj_991 (.I0(n17_adj_4157), .I1(\data_in[1] [6]), .I2(n16_adj_4156), 
            .I3(\data_in[3] [7]), .O(n26621));
    defparam i9_4_lut_adj_991.LUT_INIT = 16'hfbff;
    SB_LUT4 i4_4_lut_adj_992 (.I0(\data_in[1] [7]), .I1(\data_in[0] [0]), 
            .I2(\data_in[1] [1]), .I3(\data_in[0] [4]), .O(n10_adj_4158));
    defparam i4_4_lut_adj_992.LUT_INIT = 16'hfdff;
    SB_DFFE setpoint__i23 (.Q(setpoint[23]), .C(CLK_c), .E(n27781), .D(n5809));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_3_lut_adj_993 (.I0(\data_in[3] [4]), .I1(n10_adj_4158), .I2(\data_in[2] [7]), 
            .I3(GND_net), .O(n26689));
    defparam i5_3_lut_adj_993.LUT_INIT = 16'hdfdf;
    SB_LUT4 i2_2_lut (.I0(\data_in[2] [3]), .I1(\data_in[3] [5]), .I2(GND_net), 
            .I3(GND_net), .O(n10_adj_4159));
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i6_4_lut_adj_994 (.I0(\data_in[0] [2]), .I1(\data_in[3] [3]), 
            .I2(\data_in[3] [1]), .I3(\data_in[0] [7]), .O(n14_adj_4160));
    defparam i6_4_lut_adj_994.LUT_INIT = 16'hfeff;
    SB_DFFE setpoint__i22 (.Q(setpoint[22]), .C(CLK_c), .E(n27781), .D(n5808));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i21 (.Q(setpoint[21]), .C(CLK_c), .E(n27781), .D(n5807));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i20 (.Q(setpoint[20]), .C(CLK_c), .E(n27781), .D(n5806));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i19 (.Q(setpoint[19]), .C(CLK_c), .E(n27781), .D(n5805));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i18 (.Q(setpoint[18]), .C(CLK_c), .E(n27781), .D(n5804));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i17 (.Q(setpoint[17]), .C(CLK_c), .E(n27781), .D(n5803));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i16 (.Q(setpoint[16]), .C(CLK_c), .E(n27781), .D(n5802));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i15 (.Q(setpoint[15]), .C(CLK_c), .E(n27781), .D(n5801));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i14 (.Q(setpoint[14]), .C(CLK_c), .E(n27781), .D(n5800));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i7_4_lut_adj_995 (.I0(\data_in[3] [6]), .I1(n14_adj_4160), .I2(n10_adj_4159), 
            .I3(\data_in[2] [1]), .O(n26692));
    defparam i7_4_lut_adj_995.LUT_INIT = 16'hfffd;
    SB_LUT4 i7_4_lut_adj_996 (.I0(\data_in[2] [4]), .I1(n26692), .I2(\data_in[1] [5]), 
            .I3(n26689), .O(n18));
    defparam i7_4_lut_adj_996.LUT_INIT = 16'hfffd;
    SB_DFFE setpoint__i13 (.Q(setpoint[13]), .C(CLK_c), .E(n27781), .D(n5799));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i9_4_lut_adj_997 (.I0(\data_in[0] [6]), .I1(n18), .I2(\data_in[3] [0]), 
            .I3(n26621), .O(n20_adj_4161));
    defparam i9_4_lut_adj_997.LUT_INIT = 16'hfffd;
    SB_LUT4 i4_2_lut (.I0(\data_in[1] [0]), .I1(\data_in[0] [3]), .I2(GND_net), 
            .I3(GND_net), .O(n15_adj_4162));
    defparam i4_2_lut.LUT_INIT = 16'heeee;
    SB_DFFE setpoint__i12 (.Q(setpoint[12]), .C(CLK_c), .E(n27781), .D(n5798));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i11 (.Q(setpoint[11]), .C(CLK_c), .E(n27781), .D(n5797));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i10_4_lut_adj_998 (.I0(n15_adj_4162), .I1(n20_adj_4161), .I2(\data_in[2] [2]), 
            .I3(\data_in[1] [4]), .O(n63_c));
    defparam i10_4_lut_adj_998.LUT_INIT = 16'hfeff;
    SB_DFFE setpoint__i10 (.Q(setpoint[10]), .C(CLK_c), .E(n27781), .D(n5796));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i9 (.Q(setpoint[9]), .C(CLK_c), .E(n27781), .D(n5795));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i6_4_lut_adj_999 (.I0(\data_in[3] [6]), .I1(\data_in[0] [7]), 
            .I2(\data_in[2] [1]), .I3(n26510), .O(n16_adj_4163));
    defparam i6_4_lut_adj_999.LUT_INIT = 16'hffef;
    SB_DFFE setpoint__i8 (.Q(setpoint[8]), .C(CLK_c), .E(n27781), .D(n5794));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i7 (.Q(setpoint[7]), .C(CLK_c), .E(n27781), .D(n5793));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i6 (.Q(setpoint[6]), .C(CLK_c), .E(n27781), .D(n5792));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i7_4_lut_adj_1000 (.I0(n26621), .I1(\data_in[2] [3]), .I2(\data_in[0] [2]), 
            .I3(\data_in[3] [5]), .O(n17_adj_4164));
    defparam i7_4_lut_adj_1000.LUT_INIT = 16'hbfff;
    SB_LUT4 add_43_25_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [23]), .I2(GND_net), 
            .I3(n39097), .O(n2_adj_4165)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_25_lut.LUT_INIT = 16'h8228;
    SB_DFFE setpoint__i5 (.Q(setpoint[5]), .C(CLK_c), .E(n27781), .D(n5791));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i4 (.Q(setpoint[4]), .C(CLK_c), .E(n27781), .D(n5790));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i3 (.Q(setpoint[3]), .C(CLK_c), .E(n27781), .D(n5789));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i9_4_lut_adj_1001 (.I0(n17_adj_4164), .I1(\data_in[3] [3]), 
            .I2(n16_adj_4163), .I3(\data_in[3] [1]), .O(n63_adj_4138));
    defparam i9_4_lut_adj_1001.LUT_INIT = 16'hfbff;
    SB_DFFE setpoint__i2 (.Q(setpoint[2]), .C(CLK_c), .E(n27781), .D(n5788));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE setpoint__i1 (.Q(setpoint[1]), .C(CLK_c), .E(n27781), .D(n5787));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i8_4_lut_adj_1002 (.I0(n26692), .I1(\data_in[1] [3]), .I2(n26510), 
            .I3(\data_in[1] [2]), .O(n20_adj_4166));
    defparam i8_4_lut_adj_1002.LUT_INIT = 16'hfbff;
    SB_LUT4 i7_4_lut_adj_1003 (.I0(\data_in[2] [6]), .I1(\data_in[1] [6]), 
            .I2(\data_in[3] [7]), .I3(\data_in[0] [1]), .O(n19));
    defparam i7_4_lut_adj_1003.LUT_INIT = 16'hfeff;
    SB_LUT4 i33893_4_lut (.I0(\data_in[2] [0]), .I1(\data_in[2] [5]), .I2(\data_in[0] [5]), 
            .I3(\data_in[3] [2]), .O(n48787));
    defparam i33893_4_lut.LUT_INIT = 16'h8000;
    SB_CARRY add_43_25 (.CI(n39097), .I0(\FRAME_MATCHER.i [23]), .I1(GND_net), 
            .CO(n39098));
    SB_LUT4 i11_3_lut (.I0(n48787), .I1(n19), .I2(n20_adj_4166), .I3(GND_net), 
            .O(n63));
    defparam i11_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i1_2_lut_adj_1004 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(GND_net), .I3(GND_net), .O(n5728));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1004.LUT_INIT = 16'hbbbb;
    SB_LUT4 add_43_24_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [22]), .I2(GND_net), 
            .I3(n39096), .O(n2_adj_4167)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_24_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_4_lut_adj_1005 (.I0(n4_c), .I1(n61), .I2(n44042), .I3(n33307), 
            .O(n44079));
    defparam i1_4_lut_adj_1005.LUT_INIT = 16'hbaaa;
    SB_CARRY add_43_24 (.CI(n39096), .I0(\FRAME_MATCHER.i [22]), .I1(GND_net), 
            .CO(n39097));
    SB_LUT4 add_43_23_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [21]), .I2(GND_net), 
            .I3(n39095), .O(n2_adj_4168)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_23_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_23 (.CI(n39095), .I0(\FRAME_MATCHER.i [21]), .I1(GND_net), 
            .CO(n39096));
    SB_LUT4 i1_4_lut_adj_1006 (.I0(\FRAME_MATCHER.state_c [31]), .I1(\FRAME_MATCHER.state[0] ), 
            .I2(n44079), .I3(n4_adj_4169), .O(n43489));
    defparam i1_4_lut_adj_1006.LUT_INIT = 16'ha8a0;
    SB_DFFSS \FRAME_MATCHER.state_i31  (.Q(\FRAME_MATCHER.state_c [31]), .C(CLK_c), 
            .D(n43587), .S(n43489));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_22_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [20]), .I2(GND_net), 
            .I3(n39094), .O(n2_adj_4170)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_22_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_22 (.CI(n39094), .I0(\FRAME_MATCHER.i [20]), .I1(GND_net), 
            .CO(n39095));
    SB_LUT4 add_43_21_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [19]), .I2(GND_net), 
            .I3(n39093), .O(n2_adj_4171)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_21_lut.LUT_INIT = 16'h8228;
    SB_DFF PWMLimit_i0_i6 (.Q(PWMLimit[6]), .C(CLK_c), .D(n28272));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15337_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44095), .I2(rx_data[3]), 
            .I3(\data_in_frame[11] [3]), .O(n28400));
    defparam i15337_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15338_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44095), .I2(rx_data[2]), 
            .I3(\data_in_frame[11] [2]), .O(n28401));
    defparam i15338_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i7 (.Q(PWMLimit[7]), .C(CLK_c), .D(n28271));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15339_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44095), .I2(rx_data[1]), 
            .I3(\data_in_frame[11] [1]), .O(n28402));
    defparam i15339_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_21 (.CI(n39093), .I0(\FRAME_MATCHER.i [19]), .I1(GND_net), 
            .CO(n39094));
    SB_LUT4 add_43_20_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [18]), .I2(GND_net), 
            .I3(n39092), .O(n2_adj_4172)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_20_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_20 (.CI(n39092), .I0(\FRAME_MATCHER.i [18]), .I1(GND_net), 
            .CO(n39093));
    SB_LUT4 add_43_19_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [17]), .I2(GND_net), 
            .I3(n39091), .O(n2_adj_4173)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_19_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_19 (.CI(n39091), .I0(\FRAME_MATCHER.i [17]), .I1(GND_net), 
            .CO(n39092));
    SB_LUT4 add_43_18_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [16]), .I2(GND_net), 
            .I3(n39090), .O(n2_adj_4174)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_18_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_18 (.CI(n39090), .I0(\FRAME_MATCHER.i [16]), .I1(GND_net), 
            .CO(n39091));
    SB_LUT4 i15340_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44095), .I2(rx_data[0]), 
            .I3(\data_in_frame[11] [0]), .O(n28403));
    defparam i15340_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15325_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44095), .I2(rx_data[7]), 
            .I3(\data_in_frame[12] [7]), .O(n28388));
    defparam i15325_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15326_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44095), .I2(rx_data[6]), 
            .I3(\data_in_frame[12] [6]), .O(n28389));
    defparam i15326_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15327_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44095), .I2(rx_data[5]), 
            .I3(\data_in_frame[12] [5]), .O(n28390));
    defparam i15327_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15328_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44095), .I2(rx_data[4]), 
            .I3(\data_in_frame[12] [4]), .O(n28391));
    defparam i15328_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15329_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44095), .I2(rx_data[3]), 
            .I3(\data_in_frame[12] [3]), .O(n28392));
    defparam i15329_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15330_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44095), .I2(rx_data[2]), 
            .I3(\data_in_frame[12] [2]), .O(n28393));
    defparam i15330_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15331_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44095), .I2(rx_data[1]), 
            .I3(\data_in_frame[12] [1]), .O(n28394));
    defparam i15331_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1361_i2_3_lut (.I0(\data_in_frame[19] [1]), .I1(\data_in_frame[3] [1]), 
            .I2(n5785), .I3(GND_net), .O(n5787));
    defparam mux_1361_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_43_17_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [15]), .I2(GND_net), 
            .I3(n39089), .O(n2_adj_4176)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_17_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mux_1361_i3_3_lut (.I0(\data_in_frame[19] [2]), .I1(\data_in_frame[3] [2]), 
            .I2(n5785), .I3(GND_net), .O(n5788));
    defparam mux_1361_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1361_i4_3_lut (.I0(\data_in_frame[19] [3]), .I1(\data_in_frame[3] [3]), 
            .I2(n5785), .I3(GND_net), .O(n5789));
    defparam mux_1361_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1361_i5_3_lut (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[3] [4]), 
            .I2(n5785), .I3(GND_net), .O(n5790));
    defparam mux_1361_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1361_i6_3_lut (.I0(\data_in_frame[19] [5]), .I1(\data_in_frame[3] [5]), 
            .I2(n5785), .I3(GND_net), .O(n5791));
    defparam mux_1361_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1361_i7_3_lut (.I0(\data_in_frame[19] [6]), .I1(\data_in_frame[3] [6]), 
            .I2(n5785), .I3(GND_net), .O(n5792));
    defparam mux_1361_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15332_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44095), .I2(rx_data[0]), 
            .I3(\data_in_frame[12] [0]), .O(n28395));
    defparam i15332_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1361_i8_3_lut (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[3] [7]), 
            .I2(n5785), .I3(GND_net), .O(n5793));
    defparam mux_1361_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1361_i9_3_lut (.I0(\data_in_frame[18] [0]), .I1(\data_in_frame[2] [0]), 
            .I2(n5785), .I3(GND_net), .O(n5794));
    defparam mux_1361_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_17 (.CI(n39089), .I0(\FRAME_MATCHER.i [15]), .I1(GND_net), 
            .CO(n39090));
    SB_LUT4 i15317_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44095), .I2(rx_data[7]), 
            .I3(\data_in_frame[13] [7]), .O(n28380));
    defparam i15317_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1361_i10_3_lut (.I0(\data_in_frame[18] [1]), .I1(\data_in_frame[2] [1]), 
            .I2(n5785), .I3(GND_net), .O(n5795));
    defparam mux_1361_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1361_i11_3_lut (.I0(\data_in_frame[18] [2]), .I1(\data_in_frame[2] [2]), 
            .I2(n5785), .I3(GND_net), .O(n5796));
    defparam mux_1361_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1361_i12_3_lut (.I0(\data_in_frame[18] [3]), .I1(\data_in_frame[2] [3]), 
            .I2(n5785), .I3(GND_net), .O(n5797));
    defparam mux_1361_i12_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1361_i13_3_lut (.I0(\data_in_frame[18] [4]), .I1(\data_in_frame[2] [4]), 
            .I2(n5785), .I3(GND_net), .O(n5798));
    defparam mux_1361_i13_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_43_16_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [14]), .I2(GND_net), 
            .I3(n39088), .O(n2_adj_4178)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_16_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mux_1361_i14_3_lut (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[2] [5]), 
            .I2(n5785), .I3(GND_net), .O(n5799));
    defparam mux_1361_i14_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_16 (.CI(n39088), .I0(\FRAME_MATCHER.i [14]), .I1(GND_net), 
            .CO(n39089));
    SB_LUT4 i15318_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44095), .I2(rx_data[6]), 
            .I3(\data_in_frame[13] [6]), .O(n28381));
    defparam i15318_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 add_43_15_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [13]), .I2(GND_net), 
            .I3(n39087), .O(n2_adj_4179)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_15_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_15 (.CI(n39087), .I0(\FRAME_MATCHER.i [13]), .I1(GND_net), 
            .CO(n39088));
    SB_LUT4 mux_1361_i15_3_lut (.I0(\data_in_frame[18] [6]), .I1(\data_in_frame[2] [6]), 
            .I2(n5785), .I3(GND_net), .O(n5800));
    defparam mux_1361_i15_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1361_i16_3_lut (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[2] [7]), 
            .I2(n5785), .I3(GND_net), .O(n5801));
    defparam mux_1361_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1361_i17_3_lut (.I0(\data_in_frame[17] [0]), .I1(\data_in_frame[1] [0]), 
            .I2(n5785), .I3(GND_net), .O(n5802));
    defparam mux_1361_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1361_i18_3_lut (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[1] [1]), 
            .I2(n5785), .I3(GND_net), .O(n5803));
    defparam mux_1361_i18_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15319_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44095), .I2(rx_data[5]), 
            .I3(\data_in_frame[13] [5]), .O(n28382));
    defparam i15319_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1361_i19_3_lut (.I0(\data_in_frame[17] [2]), .I1(\data_in_frame[1] [2]), 
            .I2(n5785), .I3(GND_net), .O(n5804));
    defparam mux_1361_i19_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_43_14_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [12]), .I2(GND_net), 
            .I3(n39086), .O(n2_adj_4180)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_14_lut.LUT_INIT = 16'h8228;
    SB_LUT4 mux_1361_i20_3_lut (.I0(\data_in_frame[17] [3]), .I1(\data_in_frame[1] [3]), 
            .I2(n5785), .I3(GND_net), .O(n5805));
    defparam mux_1361_i20_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1361_i21_3_lut (.I0(\data_in_frame[17] [4]), .I1(\data_in_frame[1] [4]), 
            .I2(n5785), .I3(GND_net), .O(n5806));
    defparam mux_1361_i21_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34015_3_lut (.I0(\data_out_frame[8] [0]), .I1(\data_out_frame[9] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48967));
    defparam i34015_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34016_3_lut (.I0(\data_out_frame[10] [0]), .I1(\data_out_frame[11] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48968));
    defparam i34016_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34067_3_lut (.I0(\data_out_frame[14] [0]), .I1(\data_out_frame[15] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n49019));
    defparam i34067_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1007 (.I0(n42434), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[25] [3]), .I3(n45674), .O(n45731));
    defparam i2_3_lut_4_lut_adj_1007.LUT_INIT = 16'h9669;
    SB_LUT4 i34066_3_lut (.I0(\data_out_frame[12] [0]), .I1(\data_out_frame[13] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n49018));
    defparam i34066_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34030_3_lut (.I0(\data_out_frame[8] [6]), .I1(\data_out_frame[9] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48982));
    defparam i34030_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34031_3_lut (.I0(\data_out_frame[10] [6]), .I1(\data_out_frame[11] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48983));
    defparam i34031_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34025_3_lut (.I0(\data_out_frame[14] [6]), .I1(\data_out_frame[15] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48977));
    defparam i34025_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34024_3_lut (.I0(\data_out_frame[12] [6]), .I1(\data_out_frame[13] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48976));
    defparam i34024_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1361_i22_3_lut (.I0(\data_in_frame[17] [5]), .I1(\data_in_frame[1] [5]), 
            .I2(n5785), .I3(GND_net), .O(n5807));
    defparam mux_1361_i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 mux_1361_i23_3_lut (.I0(\data_in_frame[17] [6]), .I1(\data_in_frame[1] [6]), 
            .I2(n5785), .I3(GND_net), .O(n5808));
    defparam mux_1361_i23_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15320_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44095), .I2(rx_data[4]), 
            .I3(\data_in_frame[13] [4]), .O(n28383));
    defparam i15320_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 mux_1361_i24_3_lut (.I0(\data_in_frame[17] [7]), .I1(\data_in_frame[1] [7]), 
            .I2(n5785), .I3(GND_net), .O(n5809));
    defparam mux_1361_i24_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15321_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44095), .I2(rx_data[3]), 
            .I3(\data_in_frame[13] [3]), .O(n28384));
    defparam i15321_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF PWMLimit_i0_i8 (.Q(PWMLimit[8]), .C(CLK_c), .D(n28270));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i9 (.Q(PWMLimit[9]), .C(CLK_c), .D(n28269));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i10 (.Q(PWMLimit[10]), .C(CLK_c), .D(n28268));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i11 (.Q(PWMLimit[11]), .C(CLK_c), .D(n28267));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i12 (.Q(PWMLimit[12]), .C(CLK_c), .D(n28266));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i13 (.Q(PWMLimit[13]), .C(CLK_c), .D(n28265));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i14 (.Q(PWMLimit[14]), .C(CLK_c), .D(n28264));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i15 (.Q(PWMLimit[15]), .C(CLK_c), .D(n28263));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i16 (.Q(PWMLimit[16]), .C(CLK_c), .D(n28262));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i17 (.Q(PWMLimit[17]), .C(CLK_c), .D(n28261));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i18 (.Q(PWMLimit[18]), .C(CLK_c), .D(n28260));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i19 (.Q(PWMLimit[19]), .C(CLK_c), .D(n28259));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i20 (.Q(PWMLimit[20]), .C(CLK_c), .D(n28258));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i21 (.Q(PWMLimit[21]), .C(CLK_c), .D(n28257));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i22 (.Q(PWMLimit[22]), .C(CLK_c), .D(n28256));   // verilog/coms.v(127[12] 300[6])
    SB_DFF PWMLimit_i0_i23 (.Q(PWMLimit[23]), .C(CLK_c), .D(n28255));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i1  (.Q(\FRAME_MATCHER.state_c [1]), .C(CLK_c), 
           .D(n51636));   // verilog/coms.v(127[12] 300[6])
    SB_DFF \FRAME_MATCHER.state_i2  (.Q(\FRAME_MATCHER.state_c [2]), .C(CLK_c), 
           .D(n51637));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR byte_transmit_counter_i0_i0 (.Q(\byte_transmit_counter[0] ), 
            .C(CLK_c), .E(n27787), .D(n8825[0]), .R(n33303));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15322_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44095), .I2(rx_data[2]), 
            .I3(\data_in_frame[13] [2]), .O(n28385));
    defparam i15322_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i34033_3_lut (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[9] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48985));
    defparam i34033_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34034_3_lut (.I0(\data_out_frame[10] [5]), .I1(\data_out_frame[11] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48986));
    defparam i34034_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33971_3_lut (.I0(\data_out_frame[14] [5]), .I1(\data_out_frame[15] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48923));
    defparam i33971_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33970_3_lut (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[13] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48922));
    defparam i33970_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34036_3_lut (.I0(\data_out_frame[8] [4]), .I1(\data_out_frame[9] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48988));
    defparam i34036_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34037_3_lut (.I0(\data_out_frame[10] [4]), .I1(\data_out_frame[11] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48989));
    defparam i34037_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33935_3_lut (.I0(\data_out_frame[14] [4]), .I1(\data_out_frame[15] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48887));
    defparam i33935_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_14 (.CI(n39086), .I0(\FRAME_MATCHER.i [12]), .I1(GND_net), 
            .CO(n39087));
    SB_LUT4 i33934_3_lut (.I0(\data_out_frame[12] [4]), .I1(\data_out_frame[13] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48886));
    defparam i33934_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34039_3_lut (.I0(\data_out_frame[8] [3]), .I1(\data_out_frame[9] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48991));
    defparam i34039_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34040_3_lut (.I0(\data_out_frame[10] [3]), .I1(\data_out_frame[11] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48992));
    defparam i34040_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 add_43_13_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [11]), .I2(GND_net), 
            .I3(n39085), .O(n2_adj_4181)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_13_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i34049_3_lut (.I0(\data_out_frame[14] [3]), .I1(\data_out_frame[15] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n49001));
    defparam i34049_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34048_3_lut (.I0(\data_out_frame[12] [3]), .I1(\data_out_frame[13] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n49000));
    defparam i34048_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34051_3_lut (.I0(\data_out_frame[8] [2]), .I1(\data_out_frame[9] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n49003));
    defparam i34051_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34052_3_lut (.I0(\data_out_frame[10] [2]), .I1(\data_out_frame[11] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n49004));
    defparam i34052_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33905_3_lut (.I0(\data_out_frame[14] [2]), .I1(\data_out_frame[15] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48857));
    defparam i33905_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33904_3_lut (.I0(\data_out_frame[12] [2]), .I1(\data_out_frame[13] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48856));
    defparam i33904_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34054_3_lut (.I0(\data_out_frame[8] [1]), .I1(\data_out_frame[9] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n49006));
    defparam i34054_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20647_2_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n10));
    defparam i20647_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i34055_3_lut (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[11] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n49007));
    defparam i34055_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_13 (.CI(n39085), .I0(\FRAME_MATCHER.i [11]), .I1(GND_net), 
            .CO(n39086));
    SB_DFFSS \FRAME_MATCHER.state_i30  (.Q(\FRAME_MATCHER.state_c [30]), .C(CLK_c), 
            .D(n7_adj_4183), .S(n43477));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_12_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [10]), .I2(GND_net), 
            .I3(n39084), .O(n2_adj_4184)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_12_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i1_3_lut_adj_1008 (.I0(n61), .I1(n31_adj_4185), .I2(n24120), 
            .I3(GND_net), .O(n27771));
    defparam i1_3_lut_adj_1008.LUT_INIT = 16'h0202;
    SB_LUT4 i2_4_lut_adj_1009 (.I0(n44947), .I1(n44979), .I2(\FRAME_MATCHER.state_c [1]), 
            .I3(n69), .O(n46802));
    defparam i2_4_lut_adj_1009.LUT_INIT = 16'h0501;
    SB_CARRY add_43_12 (.CI(n39084), .I0(\FRAME_MATCHER.i [10]), .I1(GND_net), 
            .CO(n39085));
    SB_LUT4 i1_4_lut_adj_1010 (.I0(\FRAME_MATCHER.state[0] ), .I1(n24120), 
            .I2(\FRAME_MATCHER.state_c [2]), .I3(n23701), .O(n45946));
    defparam i1_4_lut_adj_1010.LUT_INIT = 16'h5040;
    SB_LUT4 add_43_11_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [9]), .I2(GND_net), 
            .I3(n39083), .O(n2_adj_4186)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_11_lut.LUT_INIT = 16'h8228;
    SB_DFFSS \FRAME_MATCHER.state_i29  (.Q(\FRAME_MATCHER.state_c [29]), .C(CLK_c), 
            .D(n33576), .S(n34368));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i28  (.Q(\FRAME_MATCHER.state_c [28]), .C(CLK_c), 
            .D(n43627), .S(n43511));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i27  (.Q(\FRAME_MATCHER.state_c [27]), .C(CLK_c), 
            .D(n33574), .S(n34366));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i26  (.Q(\FRAME_MATCHER.state_c [26]), .C(CLK_c), 
            .D(n43625), .S(n43513));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i25  (.Q(\FRAME_MATCHER.state_c [25]), .C(CLK_c), 
            .D(n33572), .S(n34364));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i24  (.Q(\FRAME_MATCHER.state_c [24]), .C(CLK_c), 
            .D(n43623), .S(n43515));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i23  (.Q(\FRAME_MATCHER.state_c [23]), .C(CLK_c), 
            .D(n43621), .S(n43517));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i22  (.Q(\FRAME_MATCHER.state_c [22]), .C(CLK_c), 
            .D(n7_adj_4187), .S(n8_adj_4188));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i21  (.Q(\FRAME_MATCHER.state_c [21]), .C(CLK_c), 
            .D(n7_adj_4189), .S(n33570));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i20  (.Q(\FRAME_MATCHER.state_c [20]), .C(CLK_c), 
            .D(n43619), .S(n43519));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_11 (.CI(n39083), .I0(\FRAME_MATCHER.i [9]), .I1(GND_net), 
            .CO(n39084));
    SB_LUT4 add_43_10_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [8]), .I2(GND_net), 
            .I3(n39082), .O(n2_adj_4190)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_10_lut.LUT_INIT = 16'h8228;
    SB_DFFSS \FRAME_MATCHER.state_i19  (.Q(\FRAME_MATCHER.state_c [19]), .C(CLK_c), 
            .D(n33568), .S(n34362));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i18  (.Q(\FRAME_MATCHER.state_c [18]), .C(CLK_c), 
            .D(n43617), .S(n43521));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i17  (.Q(\FRAME_MATCHER.state_c [17]), .C(CLK_c), 
            .D(n43615), .S(n43523));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i16  (.Q(\FRAME_MATCHER.state_c [16]), .C(CLK_c), 
            .D(n43613), .S(n43525));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i15  (.Q(\FRAME_MATCHER.state_c [15]), .C(CLK_c), 
            .D(n43611), .S(n43527));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i14  (.Q(\FRAME_MATCHER.state_c [14]), .C(CLK_c), 
            .D(n43609), .S(n43529));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i13  (.Q(\FRAME_MATCHER.state_c [13]), .C(CLK_c), 
            .D(n43607), .S(n43531));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i12  (.Q(\FRAME_MATCHER.state_c [12]), .C(CLK_c), 
            .D(n43605), .S(n43533));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i11  (.Q(\FRAME_MATCHER.state_c [11]), .C(CLK_c), 
            .D(n43603), .S(n43535));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i10  (.Q(\FRAME_MATCHER.state_c [10]), .C(CLK_c), 
            .D(n43601), .S(n43537));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i9  (.Q(\FRAME_MATCHER.state_c [9]), .C(CLK_c), 
            .D(n43599), .S(n43539));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i8  (.Q(\FRAME_MATCHER.state_c [8]), .C(CLK_c), 
            .D(n43597), .S(n43541));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i7  (.Q(\FRAME_MATCHER.state_c [7]), .C(CLK_c), 
            .D(n43595), .S(n43543));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i6  (.Q(\FRAME_MATCHER.state_c [6]), .C(CLK_c), 
            .D(n43593), .S(n43545));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i5  (.Q(\FRAME_MATCHER.state_c [5]), .C(CLK_c), 
            .D(n43591), .S(n43547));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i4  (.Q(\FRAME_MATCHER.state_c [4]), .C(CLK_c), 
            .D(n43589), .S(n43491));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.state_i3  (.Q(\FRAME_MATCHER.state [3]), .C(CLK_c), 
            .D(n43481), .S(n10_adj_4133));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15323_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44095), .I2(rx_data[1]), 
            .I3(\data_in_frame[13] [1]), .O(n28386));
    defparam i15323_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_CARRY add_43_10 (.CI(n39082), .I0(\FRAME_MATCHER.i [8]), .I1(GND_net), 
            .CO(n39083));
    SB_LUT4 i1_4_lut_adj_1011 (.I0(n45946), .I1(n5728), .I2(\FRAME_MATCHER.state_c [2]), 
            .I3(\FRAME_MATCHER.state_31__N_2624 [3]), .O(n14_adj_4191));
    defparam i1_4_lut_adj_1011.LUT_INIT = 16'haaab;
    SB_LUT4 add_43_9_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [7]), .I2(GND_net), 
            .I3(n39081), .O(n2_adj_4192)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_9_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i36073_4_lut (.I0(n69), .I1(n34823), .I2(n44989), .I3(n14_adj_4191), 
            .O(n12_adj_4193));
    defparam i36073_4_lut.LUT_INIT = 16'h23af;
    SB_CARRY add_43_9 (.CI(n39081), .I0(\FRAME_MATCHER.i [7]), .I1(GND_net), 
            .CO(n39082));
    SB_LUT4 i30089_2_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n44977), .I2(GND_net), 
            .I3(GND_net), .O(n44979));
    defparam i30089_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1_2_lut_adj_1012 (.I0(n44977), .I1(n34823), .I2(GND_net), 
            .I3(GND_net), .O(n67));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1012.LUT_INIT = 16'h4444;
    SB_LUT4 i14969_2_lut (.I0(n28031), .I1(n34823), .I2(GND_net), .I3(GND_net), 
            .O(n28032));   // verilog/coms.v(127[12] 300[6])
    defparam i14969_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_4_lut_adj_1013 (.I0(\FRAME_MATCHER.state_c [1]), .I1(n44989), 
            .I2(\FRAME_MATCHER.state_c [2]), .I3(n67), .O(n28031));
    defparam i1_4_lut_adj_1013.LUT_INIT = 16'h3733;
    SB_LUT4 i15324_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44095), .I2(rx_data[0]), 
            .I3(\data_in_frame[13] [0]), .O(n28387));
    defparam i15324_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i33902_3_lut (.I0(\data_out_frame[14] [1]), .I1(\data_out_frame[15] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48854));
    defparam i33902_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33901_3_lut (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[13] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48853));
    defparam i33901_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1014 (.I0(n42434), .I1(\data_out_frame[25] [4]), 
            .I2(n41553), .I3(GND_net), .O(n27172));
    defparam i1_2_lut_3_lut_adj_1014.LUT_INIT = 16'h9696;
    SB_LUT4 add_43_8_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [6]), .I2(GND_net), 
            .I3(n39080), .O(n2_adj_4194)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_8_lut.LUT_INIT = 16'h8228;
    SB_DFFE data_out_frame_0___i224 (.Q(\data_out_frame[27] [7]), .C(CLK_c), 
            .E(n27912), .D(n44428));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_8 (.CI(n39080), .I0(\FRAME_MATCHER.i [6]), .I1(GND_net), 
            .CO(n39081));
    SB_DFFE data_out_frame_0___i223 (.Q(\data_out_frame[27] [6]), .C(CLK_c), 
            .E(n27912), .D(n27172));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i222 (.Q(\data_out_frame[27] [5]), .C(CLK_c), 
            .E(n27912), .D(n45731));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i221 (.Q(\data_out_frame[27] [4]), .C(CLK_c), 
            .E(n27912), .D(n44489));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i220 (.Q(\data_out_frame[27] [3]), .C(CLK_c), 
            .E(n27912), .D(n45719));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i219 (.Q(\data_out_frame[27] [2]), .C(CLK_c), 
            .E(n27912), .D(n42395));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i218 (.Q(\data_out_frame[27] [1]), .C(CLK_c), 
            .E(n27912), .D(n42381));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i217 (.Q(\data_out_frame[27] [0]), .C(CLK_c), 
            .E(n27912), .D(n41565));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i216 (.Q(\data_out_frame[26] [7]), .C(CLK_c), 
            .E(n27912), .D(n45769));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i215 (.Q(\data_out_frame[26] [6]), .C(CLK_c), 
            .E(n27912), .D(n45628));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i214 (.Q(\data_out_frame[26] [5]), .C(CLK_c), 
            .E(n27912), .D(n46698));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i213 (.Q(\data_out_frame[26] [4]), .C(CLK_c), 
            .E(n27912), .D(n46700));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i212 (.Q(\data_out_frame[26] [3]), .C(CLK_c), 
            .E(n27912), .D(n45867));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i211 (.Q(\data_out_frame[26] [2]), .C(CLK_c), 
            .E(n27912), .D(n45555));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i210 (.Q(\data_out_frame[26] [1]), .C(CLK_c), 
            .E(n27912), .D(n45401));   // verilog/coms.v(127[12] 300[6])
    SB_DFFE data_out_frame_0___i209 (.Q(\data_out_frame[26] [0]), .C(CLK_c), 
            .E(n27912), .D(n46095));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 add_43_7_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [5]), .I2(GND_net), 
            .I3(n39079), .O(n2_adj_4195)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_7_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_7 (.CI(n39079), .I0(\FRAME_MATCHER.i [5]), .I1(GND_net), 
            .CO(n39080));
    SB_LUT4 add_43_6_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [4]), .I2(GND_net), 
            .I3(n39078), .O(n2_adj_4196)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_6_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i4_3_lut_4_lut (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[18] [5]), 
            .I2(\data_out_frame[18] [3]), .I3(n41615), .O(n11));   // verilog/coms.v(85[17:28])
    defparam i4_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFFSS \FRAME_MATCHER.i_i31  (.Q(\FRAME_MATCHER.i[31] ), .C(CLK_c), 
            .D(n2_adj_4143), .S(n3_adj_4197));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i30  (.Q(\FRAME_MATCHER.i [30]), .C(CLK_c), 
            .D(n2_adj_4144), .S(n3_adj_4198));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i29  (.Q(\FRAME_MATCHER.i [29]), .C(CLK_c), 
            .D(n2_adj_4145), .S(n3_adj_4199));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i28  (.Q(\FRAME_MATCHER.i [28]), .C(CLK_c), 
            .D(n2_adj_4146), .S(n3_adj_4200));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i27  (.Q(\FRAME_MATCHER.i [27]), .C(CLK_c), 
            .D(n2_adj_4148), .S(n3_adj_4201));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i26  (.Q(\FRAME_MATCHER.i [26]), .C(CLK_c), 
            .D(n2_adj_4149), .S(n3_adj_4202));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i25  (.Q(\FRAME_MATCHER.i [25]), .C(CLK_c), 
            .D(n2_adj_4151), .S(n3_adj_4203));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i24  (.Q(\FRAME_MATCHER.i [24]), .C(CLK_c), 
            .D(n2_adj_4153), .S(n3_adj_4204));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i23  (.Q(\FRAME_MATCHER.i [23]), .C(CLK_c), 
            .D(n2_adj_4165), .S(n3_adj_4205));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i22  (.Q(\FRAME_MATCHER.i [22]), .C(CLK_c), 
            .D(n2_adj_4167), .S(n3_adj_4206));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i21  (.Q(\FRAME_MATCHER.i [21]), .C(CLK_c), 
            .D(n2_adj_4168), .S(n3_adj_4207));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i20  (.Q(\FRAME_MATCHER.i [20]), .C(CLK_c), 
            .D(n2_adj_4170), .S(n3_adj_4208));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i19  (.Q(\FRAME_MATCHER.i [19]), .C(CLK_c), 
            .D(n2_adj_4171), .S(n3_adj_4209));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i18  (.Q(\FRAME_MATCHER.i [18]), .C(CLK_c), 
            .D(n2_adj_4172), .S(n3_adj_4210));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i17  (.Q(\FRAME_MATCHER.i [17]), .C(CLK_c), 
            .D(n2_adj_4173), .S(n3_adj_4211));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i16  (.Q(\FRAME_MATCHER.i [16]), .C(CLK_c), 
            .D(n2_adj_4174), .S(n3_adj_4212));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i15  (.Q(\FRAME_MATCHER.i [15]), .C(CLK_c), 
            .D(n2_adj_4176), .S(n3_adj_4213));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i14  (.Q(\FRAME_MATCHER.i [14]), .C(CLK_c), 
            .D(n2_adj_4178), .S(n3_adj_4214));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i13  (.Q(\FRAME_MATCHER.i [13]), .C(CLK_c), 
            .D(n2_adj_4179), .S(n3_adj_4215));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i12  (.Q(\FRAME_MATCHER.i [12]), .C(CLK_c), 
            .D(n2_adj_4180), .S(n3_adj_4216));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i11  (.Q(\FRAME_MATCHER.i [11]), .C(CLK_c), 
            .D(n2_adj_4181), .S(n3_adj_4217));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i10  (.Q(\FRAME_MATCHER.i [10]), .C(CLK_c), 
            .D(n2_adj_4184), .S(n3_adj_4218));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i9  (.Q(\FRAME_MATCHER.i [9]), .C(CLK_c), 
            .D(n2_adj_4186), .S(n3_adj_4219));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i8  (.Q(\FRAME_MATCHER.i [8]), .C(CLK_c), 
            .D(n2_adj_4190), .S(n3_adj_4220));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i7  (.Q(\FRAME_MATCHER.i [7]), .C(CLK_c), 
            .D(n2_adj_4192), .S(n3_adj_4221));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i6  (.Q(\FRAME_MATCHER.i [6]), .C(CLK_c), 
            .D(n2_adj_4194), .S(n3_adj_4222));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i5  (.Q(\FRAME_MATCHER.i [5]), .C(CLK_c), 
            .D(n2_adj_4195), .S(n3_adj_4223));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i4  (.Q(\FRAME_MATCHER.i [4]), .C(CLK_c), 
            .D(n2_adj_4196), .S(n3_adj_4224));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i3  (.Q(\FRAME_MATCHER.i [3]), .C(CLK_c), 
            .D(n2_adj_4225), .S(n3_adj_4226));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i2  (.Q(\FRAME_MATCHER.i [2]), .C(CLK_c), 
            .D(n2_adj_4227), .S(n3_adj_4228));   // verilog/coms.v(127[12] 300[6])
    SB_DFFSS \FRAME_MATCHER.i_i1  (.Q(\FRAME_MATCHER.i [1]), .C(CLK_c), 
            .D(n2_adj_4229), .S(n3_adj_4230));   // verilog/coms.v(127[12] 300[6])
    SB_CARRY add_43_6 (.CI(n39078), .I0(\FRAME_MATCHER.i [4]), .I1(GND_net), 
            .CO(n39079));
    SB_LUT4 add_43_5_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [3]), .I2(GND_net), 
            .I3(n39077), .O(n2_adj_4225)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_5_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_5 (.CI(n39077), .I0(\FRAME_MATCHER.i [3]), .I1(GND_net), 
            .CO(n39078));
    SB_LUT4 add_43_4_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [2]), .I2(GND_net), 
            .I3(n39076), .O(n2_adj_4227)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_4_lut.LUT_INIT = 16'h8228;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut (.I0(byte_transmit_counter[3]), 
            .I1(n50305), .I2(n49814), .I3(byte_transmit_counter[4]), .O(n51627));
    defparam byte_transmit_counter_3__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n51627_bdd_4_lut (.I0(n51627), .I1(n51510), .I2(n7_adj_4231), 
            .I3(byte_transmit_counter[4]), .O(tx_data[1]));
    defparam n51627_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15309_3_lut_4_lut (.I0(n8_adj_4232), .I1(n44095), .I2(rx_data[7]), 
            .I3(\data_in_frame[14] [7]), .O(n28372));
    defparam i15309_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_36635 (.I0(byte_transmit_counter[3]), 
            .I1(n50303), .I2(n49811), .I3(byte_transmit_counter[4]), .O(n51621));
    defparam byte_transmit_counter_3__bdd_4_lut_36635.LUT_INIT = 16'he4aa;
    SB_LUT4 n51621_bdd_4_lut (.I0(n51621), .I1(n51504), .I2(n7_adj_4233), 
            .I3(byte_transmit_counter[4]), .O(tx_data[2]));
    defparam n51621_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_36630 (.I0(byte_transmit_counter[3]), 
            .I1(n50299), .I2(n49808), .I3(byte_transmit_counter[4]), .O(n51615));
    defparam byte_transmit_counter_3__bdd_4_lut_36630.LUT_INIT = 16'he4aa;
    SB_LUT4 i34018_3_lut (.I0(\data_out_frame[8] [7]), .I1(\data_out_frame[9] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48970));
    defparam i34018_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_4 (.CI(n39076), .I0(\FRAME_MATCHER.i [2]), .I1(GND_net), 
            .CO(n39077));
    SB_LUT4 add_43_3_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [1]), .I2(GND_net), 
            .I3(n39075), .O(n2_adj_4229)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_3_lut.LUT_INIT = 16'h8228;
    SB_CARRY add_43_3 (.CI(n39075), .I0(\FRAME_MATCHER.i [1]), .I1(GND_net), 
            .CO(n39076));
    SB_LUT4 add_43_2_lut (.I0(n2482), .I1(\FRAME_MATCHER.i [0]), .I2(n161), 
            .I3(GND_net), .O(n2)) /* synthesis syn_instantiated=1 */ ;
    defparam add_43_2_lut.LUT_INIT = 16'h8228;
    SB_LUT4 i34019_3_lut (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[11] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48971));
    defparam i34019_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34064_3_lut (.I0(\data_out_frame[14] [7]), .I1(\data_out_frame[15] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n49016));
    defparam i34064_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34063_3_lut (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[13] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n49015));
    defparam i34063_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33962_3_lut (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[7] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48914));
    defparam i33962_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33963_4_lut (.I0(n48914), .I1(byte_transmit_counter[1]), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n48915));
    defparam i33963_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i33961_3_lut (.I0(\data_out_frame[4] [0]), .I1(\data_out_frame[5] [0]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48913));
    defparam i33961_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15310_3_lut_4_lut (.I0(n8_adj_4232), .I1(n44095), .I2(rx_data[6]), 
            .I3(\data_in_frame[14] [6]), .O(n28373));
    defparam i15310_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i35051_2_lut (.I0(n51582), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n49820));
    defparam i35051_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i33932_4_lut (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[23] [0]), 
            .I2(byte_transmit_counter[1]), .I3(\byte_transmit_counter[0] ), 
            .O(n48884));
    defparam i33932_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i35468_3_lut (.I0(n51432), .I1(n48884), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n50421));
    defparam i35468_3_lut.LUT_INIT = 16'hcaca;
    SB_CARRY add_43_2 (.CI(GND_net), .I0(\FRAME_MATCHER.i [0]), .I1(n161), 
            .CO(n39075));
    SB_LUT4 n51615_bdd_4_lut (.I0(n51615), .I1(n51498), .I2(n7_adj_4234), 
            .I3(byte_transmit_counter[4]), .O(tx_data[3]));
    defparam n51615_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF \FRAME_MATCHER.state_i0  (.Q(\FRAME_MATCHER.state[0] ), .C(CLK_c), 
           .D(n43485));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15311_3_lut_4_lut (.I0(n8_adj_4232), .I1(n44095), .I2(rx_data[5]), 
            .I3(\data_in_frame[14] [5]), .O(n28374));
    defparam i15311_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_36625 (.I0(byte_transmit_counter[3]), 
            .I1(n51414), .I2(n49805), .I3(byte_transmit_counter[4]), .O(n51603));
    defparam byte_transmit_counter_3__bdd_4_lut_36625.LUT_INIT = 16'he4aa;
    SB_LUT4 n51603_bdd_4_lut (.I0(n51603), .I1(n51492), .I2(n7_adj_4235), 
            .I3(byte_transmit_counter[4]), .O(tx_data[4]));
    defparam n51603_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_36615 (.I0(byte_transmit_counter[3]), 
            .I1(n51420), .I2(n49802), .I3(byte_transmit_counter[4]), .O(n51597));
    defparam byte_transmit_counter_3__bdd_4_lut_36615.LUT_INIT = 16'he4aa;
    SB_LUT4 n51597_bdd_4_lut (.I0(n51597), .I1(n51486), .I2(n7_adj_4236), 
            .I3(byte_transmit_counter[4]), .O(tx_data[5]));
    defparam n51597_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_36610 (.I0(byte_transmit_counter[3]), 
            .I1(n51426), .I2(n49817), .I3(byte_transmit_counter[4]), .O(n51591));
    defparam byte_transmit_counter_3__bdd_4_lut_36610.LUT_INIT = 16'he4aa;
    SB_LUT4 n51591_bdd_4_lut (.I0(n51591), .I1(n51480), .I2(n7_adj_4237), 
            .I3(byte_transmit_counter[4]), .O(tx_data[6]));
    defparam n51591_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_36605 (.I0(byte_transmit_counter[3]), 
            .I1(n50287), .I2(n49799), .I3(byte_transmit_counter[4]), .O(n51585));
    defparam byte_transmit_counter_3__bdd_4_lut_36605.LUT_INIT = 16'he4aa;
    SB_LUT4 n51585_bdd_4_lut (.I0(n51585), .I1(n51516), .I2(n7_adj_4238), 
            .I3(byte_transmit_counter[4]), .O(tx_data[7]));
    defparam n51585_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [0]), .I2(\data_out_frame[27] [0]), 
            .I3(byte_transmit_counter[1]), .O(n51579));
    defparam byte_transmit_counter_0__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n51579_bdd_4_lut (.I0(n51579), .I1(\data_out_frame[25] [0]), 
            .I2(\data_out_frame[24] [0]), .I3(byte_transmit_counter[1]), 
            .O(n51582));
    defparam n51579_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36595 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [1]), .I2(\data_out_frame[27] [1]), 
            .I3(byte_transmit_counter[1]), .O(n51573));
    defparam byte_transmit_counter_0__bdd_4_lut_36595.LUT_INIT = 16'he4aa;
    SB_LUT4 n51573_bdd_4_lut (.I0(n51573), .I1(\data_out_frame[25] [1]), 
            .I2(\data_out_frame[24] [1]), .I3(byte_transmit_counter[1]), 
            .O(n51576));
    defparam n51573_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36590 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [2]), .I2(\data_out_frame[27] [2]), 
            .I3(byte_transmit_counter[1]), .O(n51567));
    defparam byte_transmit_counter_0__bdd_4_lut_36590.LUT_INIT = 16'he4aa;
    SB_LUT4 n51567_bdd_4_lut (.I0(n51567), .I1(\data_out_frame[25] [2]), 
            .I2(\data_out_frame[24] [2]), .I3(byte_transmit_counter[1]), 
            .O(n51570));
    defparam n51567_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36585 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [3]), .I2(\data_out_frame[27] [3]), 
            .I3(byte_transmit_counter[1]), .O(n51561));
    defparam byte_transmit_counter_0__bdd_4_lut_36585.LUT_INIT = 16'he4aa;
    SB_LUT4 n51561_bdd_4_lut (.I0(n51561), .I1(\data_out_frame[25] [3]), 
            .I2(\data_out_frame[24] [3]), .I3(byte_transmit_counter[1]), 
            .O(n51564));
    defparam n51561_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15312_3_lut_4_lut (.I0(n8_adj_4232), .I1(n44095), .I2(rx_data[4]), 
            .I3(\data_in_frame[14] [4]), .O(n28375));
    defparam i15312_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36580 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [4]), .I2(\data_out_frame[27] [4]), 
            .I3(byte_transmit_counter[1]), .O(n51555));
    defparam byte_transmit_counter_0__bdd_4_lut_36580.LUT_INIT = 16'he4aa;
    SB_LUT4 n51555_bdd_4_lut (.I0(n51555), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[24] [4]), .I3(byte_transmit_counter[1]), 
            .O(n51558));
    defparam n51555_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36575 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [5]), .I2(\data_out_frame[27] [5]), 
            .I3(byte_transmit_counter[1]), .O(n51549));
    defparam byte_transmit_counter_0__bdd_4_lut_36575.LUT_INIT = 16'he4aa;
    SB_LUT4 n51549_bdd_4_lut (.I0(n51549), .I1(\data_out_frame[25] [5]), 
            .I2(\data_out_frame[24] [5]), .I3(byte_transmit_counter[1]), 
            .O(n51552));
    defparam n51549_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36570 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [6]), .I2(\data_out_frame[27] [6]), 
            .I3(byte_transmit_counter[1]), .O(n51543));
    defparam byte_transmit_counter_0__bdd_4_lut_36570.LUT_INIT = 16'he4aa;
    SB_LUT4 n51543_bdd_4_lut (.I0(n51543), .I1(\data_out_frame[25] [6]), 
            .I2(\data_out_frame[24] [6]), .I3(byte_transmit_counter[1]), 
            .O(n51546));
    defparam n51543_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36565 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[26] [7]), .I2(\data_out_frame[27] [7]), 
            .I3(byte_transmit_counter[1]), .O(n51537));
    defparam byte_transmit_counter_0__bdd_4_lut_36565.LUT_INIT = 16'he4aa;
    SB_LUT4 n51537_bdd_4_lut (.I0(n51537), .I1(\data_out_frame[25] [7]), 
            .I2(\data_out_frame[24] [7]), .I3(byte_transmit_counter[1]), 
            .O(n51540));
    defparam n51537_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_3__bdd_4_lut_36600 (.I0(byte_transmit_counter[3]), 
            .I1(n50421), .I2(n49820), .I3(byte_transmit_counter[4]), .O(n51531));
    defparam byte_transmit_counter_3__bdd_4_lut_36600.LUT_INIT = 16'he4aa;
    SB_LUT4 n51531_bdd_4_lut (.I0(n51531), .I1(n51474), .I2(n7_adj_4239), 
            .I3(byte_transmit_counter[4]), .O(tx_data[0]));
    defparam n51531_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut (.I0(byte_transmit_counter[1]), 
            .I1(n49015), .I2(n49016), .I3(\byte_transmit_counter[2] ), 
            .O(n51513));
    defparam byte_transmit_counter_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n51513_bdd_4_lut (.I0(n51513), .I1(n48971), .I2(n48970), .I3(\byte_transmit_counter[2] ), 
            .O(n51516));
    defparam n51513_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2_2_lut_4_lut (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[10] [7]), 
            .I2(\data_out_frame[13] [3]), .I3(\data_out_frame[8] [7]), .O(n10_adj_4240));   // verilog/coms.v(85[17:28])
    defparam i2_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1015 (.I0(n42361), .I1(\data_out_frame[20] [2]), 
            .I2(n26249), .I3(\data_out_frame[20] [3]), .O(n42427));
    defparam i2_3_lut_4_lut_adj_1015.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1016 (.I0(\data_out_frame[18]_c [1]), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[18][0] ), .I3(\data_out_frame[17] [6]), 
            .O(n44195));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1016.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[6] [2]), 
            .I2(n27539), .I3(\data_out_frame[8] [7]), .O(n14_adj_4241));   // verilog/coms.v(74[16:43])
    defparam i5_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [4]), 
            .I2(\data_out_frame[20] [7]), .I3(\data_out_frame[20] [6]), 
            .O(n44694));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h6996;
    SB_DFF PWMLimit_i0_i0 (.Q(PWMLimit[0]), .C(CLK_c), .D(n28214));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i36410_2_lut (.I0(n34527), .I1(n6_adj_4242), .I2(GND_net), 
            .I3(GND_net), .O(tx_transmit_N_3413));
    defparam i36410_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i1_2_lut_4_lut_adj_1017 (.I0(n27546), .I1(n44506), .I2(n27497), 
            .I3(\data_out_frame[19] [5]), .O(n41521));
    defparam i1_2_lut_4_lut_adj_1017.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_4_lut_adj_1018 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[17] [5]), 
            .I2(n10_adj_4243), .I3(n41525), .O(n42363));
    defparam i5_3_lut_4_lut_adj_1018.LUT_INIT = 16'h6996;
    SB_LUT4 select_427_Select_0_i3_2_lut (.I0(\FRAME_MATCHER.i [0]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3));
    defparam select_427_Select_0_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_36543 (.I0(byte_transmit_counter[1]), 
            .I1(n48853), .I2(n48854), .I3(\byte_transmit_counter[2] ), 
            .O(n51507));
    defparam byte_transmit_counter_1__bdd_4_lut_36543.LUT_INIT = 16'he4aa;
    SB_DFFESR driver_enable_3875 (.Q(DE_c), .C(CLK_c), .E(n28031), .D(n73), 
            .R(n28032));   // verilog/coms.v(127[12] 300[6])
    SB_DFFESR LED_3874 (.Q(LED_c), .C(CLK_c), .E(n12_adj_4193), .D(n44_adj_4244), 
            .R(n46802));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n51507_bdd_4_lut (.I0(n51507), .I1(n49007), .I2(n49006), .I3(\byte_transmit_counter[2] ), 
            .O(n51510));
    defparam n51507_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_36538 (.I0(byte_transmit_counter[1]), 
            .I1(n48856), .I2(n48857), .I3(\byte_transmit_counter[2] ), 
            .O(n51501));
    defparam byte_transmit_counter_1__bdd_4_lut_36538.LUT_INIT = 16'he4aa;
    SB_LUT4 n51501_bdd_4_lut (.I0(n51501), .I1(n49004), .I2(n49003), .I3(\byte_transmit_counter[2] ), 
            .O(n51504));
    defparam n51501_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_4_lut_adj_1019 (.I0(n42363), .I1(\data_out_frame[20] [1]), 
            .I2(\data_out_frame[20] [3]), .I3(n42361), .O(n42444));
    defparam i1_2_lut_4_lut_adj_1019.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_36533 (.I0(byte_transmit_counter[1]), 
            .I1(n49000), .I2(n49001), .I3(\byte_transmit_counter[2] ), 
            .O(n51495));
    defparam byte_transmit_counter_1__bdd_4_lut_36533.LUT_INIT = 16'he4aa;
    SB_LUT4 n51495_bdd_4_lut (.I0(n51495), .I1(n48992), .I2(n48991), .I3(\byte_transmit_counter[2] ), 
            .O(n51498));
    defparam n51495_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_36528 (.I0(byte_transmit_counter[1]), 
            .I1(n48886), .I2(n48887), .I3(\byte_transmit_counter[2] ), 
            .O(n51489));
    defparam byte_transmit_counter_1__bdd_4_lut_36528.LUT_INIT = 16'he4aa;
    SB_LUT4 n51489_bdd_4_lut (.I0(n51489), .I1(n48989), .I2(n48988), .I3(\byte_transmit_counter[2] ), 
            .O(n51492));
    defparam n51489_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1020 (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[20] [3]), 
            .I2(n42361), .I3(GND_net), .O(n44531));
    defparam i1_2_lut_3_lut_adj_1020.LUT_INIT = 16'h9696;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_36523 (.I0(byte_transmit_counter[1]), 
            .I1(n48922), .I2(n48923), .I3(\byte_transmit_counter[2] ), 
            .O(n51483));
    defparam byte_transmit_counter_1__bdd_4_lut_36523.LUT_INIT = 16'he4aa;
    SB_LUT4 n51483_bdd_4_lut (.I0(n51483), .I1(n48986), .I2(n48985), .I3(\byte_transmit_counter[2] ), 
            .O(n51486));
    defparam n51483_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1021 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[19] [6]), 
            .I2(n44506), .I3(GND_net), .O(n6_adj_4245));
    defparam i1_2_lut_3_lut_adj_1021.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut (.I0(n27497), .I1(\data_out_frame[19] [3]), .I2(\data_out_frame[19] [4]), 
            .I3(n44445), .O(n42333));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h9669;
    SB_LUT4 i20520_2_lut_3_lut (.I0(n2482), .I1(rx_data_ready), .I2(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I3(GND_net), .O(n33565));
    defparam i20520_2_lut_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_36518 (.I0(byte_transmit_counter[1]), 
            .I1(n48976), .I2(n48977), .I3(\byte_transmit_counter[2] ), 
            .O(n51477));
    defparam byte_transmit_counter_1__bdd_4_lut_36518.LUT_INIT = 16'he4aa;
    SB_LUT4 n51477_bdd_4_lut (.I0(n51477), .I1(n48983), .I2(n48982), .I3(\byte_transmit_counter[2] ), 
            .O(n51480));
    defparam n51477_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1022 (.I0(\FRAME_MATCHER.i_31__N_2526 ), .I1(\FRAME_MATCHER.i_31__N_2524 ), 
            .I2(n74), .I3(GND_net), .O(n2482));
    defparam i1_2_lut_3_lut_adj_1022.LUT_INIT = 16'hefef;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_36513 (.I0(byte_transmit_counter[1]), 
            .I1(n49018), .I2(n49019), .I3(\byte_transmit_counter[2] ), 
            .O(n51471));
    defparam byte_transmit_counter_1__bdd_4_lut_36513.LUT_INIT = 16'he4aa;
    SB_LUT4 n51471_bdd_4_lut (.I0(n51471), .I1(n48968), .I2(n48967), .I3(\byte_transmit_counter[2] ), 
            .O(n51474));
    defparam n51471_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1023 (.I0(n26473), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(\FRAME_MATCHER.state_c [2]), .I3(GND_net), .O(n74));
    defparam i1_2_lut_3_lut_adj_1023.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_3_lut_adj_1024 (.I0(\FRAME_MATCHER.state[0] ), .I1(n33298), 
            .I2(\FRAME_MATCHER.state [3]), .I3(GND_net), .O(n26473));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1024.LUT_INIT = 16'hfdfd;
    SB_DFF control_mode_i0_i0 (.Q(control_mode[0]), .C(CLK_c), .D(n28213));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i33781_2_lut_3_lut_4_lut (.I0(n26834), .I1(\data_in_frame[2] [5]), 
            .I2(\data_in_frame[0] [4]), .I3(\data_in_frame[0] [3]), .O(n48673));
    defparam i33781_2_lut_3_lut_4_lut.LUT_INIT = 16'hebbe;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(n23831), .I1(n771), .I2(\FRAME_MATCHER.state_c [1]), 
            .I3(\FRAME_MATCHER.state_c [2]), .O(n44055));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_4_lut_adj_1025 (.I0(n42291), .I1(n42322), .I2(n46232), 
            .I3(\data_in_frame[19] [7]), .O(n44537));
    defparam i1_4_lut_adj_1025.LUT_INIT = 16'h6996;
    SB_LUT4 i34005_4_lut (.I0(\data_out_frame[6] [7]), .I1(\byte_transmit_counter[0] ), 
            .I2(\byte_transmit_counter[2] ), .I3(\data_out_frame[7] [7]), 
            .O(n48957));
    defparam i34005_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i34003_3_lut (.I0(\data_out_frame[4] [7]), .I1(\data_out_frame[5] [7]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48955));
    defparam i34003_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1026 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [5]), 
            .I2(n41601), .I3(GND_net), .O(n44662));
    defparam i1_2_lut_3_lut_adj_1026.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1027 (.I0(n23831), .I1(n771), .I2(n26473), 
            .I3(n73), .O(n1));
    defparam i1_2_lut_3_lut_4_lut_adj_1027.LUT_INIT = 16'h0200;
    SB_LUT4 i1_2_lut_adj_1028 (.I0(\data_in_frame[14] [5]), .I1(\data_in_frame[14] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26749));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1028.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1029 (.I0(\data_in_frame[18] [7]), .I1(\data_in_frame[18] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n26890));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1029.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1030 (.I0(\data_out_frame[15] [4]), .I1(\data_out_frame[15] [5]), 
            .I2(\data_out_frame[13] [4]), .I3(n26226), .O(n44240));
    defparam i2_3_lut_4_lut_adj_1030.LUT_INIT = 16'h6996;
    SB_LUT4 i8_3_lut_4_lut (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[24] [2]), 
            .I2(\data_out_frame[24] [0]), .I3(n44129), .O(n23));   // verilog/coms.v(78[16:27])
    defparam i8_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i35041_2_lut (.I0(n51540), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n49799));
    defparam i35041_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i33956_4_lut (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[23] [7]), 
            .I2(byte_transmit_counter[1]), .I3(\byte_transmit_counter[0] ), 
            .O(n48908));
    defparam i33956_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i35334_3_lut (.I0(n51456), .I1(n48908), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n50287));
    defparam i35334_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2_3_lut_4_lut_adj_1031 (.I0(\data_out_frame[24] [1]), .I1(\data_out_frame[24] [2]), 
            .I2(n44687), .I3(n41437), .O(n44381));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_4_lut_adj_1031.LUT_INIT = 16'h9669;
    SB_LUT4 i33999_4_lut (.I0(\data_out_frame[6] [6]), .I1(\byte_transmit_counter[0] ), 
            .I2(\byte_transmit_counter[2] ), .I3(\data_out_frame[7] [6]), 
            .O(n48951));
    defparam i33999_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i33997_3_lut (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [6]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48949));
    defparam i33997_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1032 (.I0(\data_in_frame[15] [7]), .I1(\data_in_frame[16] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n44585));
    defparam i1_2_lut_adj_1032.LUT_INIT = 16'h6666;
    SB_LUT4 i33992_3_lut (.I0(\data_out_frame[6] [5]), .I1(\data_out_frame[7] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48944));
    defparam i33992_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33993_4_lut (.I0(n48944), .I1(byte_transmit_counter[1]), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n48945));
    defparam i33993_4_lut.LUT_INIT = 16'ha3a0;
    SB_LUT4 i33991_3_lut (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [5]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48943));
    defparam i33991_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1033 (.I0(\data_in_frame[15] [4]), .I1(\data_in_frame[15] [2]), 
            .I2(\data_in_frame[14] [1]), .I3(\data_in_frame[14] [3]), .O(n48411));
    defparam i1_4_lut_adj_1033.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1034 (.I0(n48411), .I1(n44754), .I2(\data_in_frame[12] [1]), 
            .I3(\data_in_frame[18] [1]), .O(n48423));
    defparam i1_4_lut_adj_1034.LUT_INIT = 16'h6996;
    SB_LUT4 i35056_2_lut (.I0(n51552), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n49802));
    defparam i35056_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12_4_lut (.I0(\data_in_frame[10] [6]), .I1(n41447), .I2(n26854), 
            .I3(n27312), .O(n28));
    defparam i12_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1035 (.I0(\data_in_frame[12] [0]), .I1(\data_in_frame[16] [4]), 
            .I2(\data_in_frame[13] [5]), .I3(\data_in_frame[16] [5]), .O(n48413));
    defparam i1_4_lut_adj_1035.LUT_INIT = 16'h6996;
    SB_LUT4 i33986_3_lut (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[7] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48938));
    defparam i33986_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1036 (.I0(n44521), .I1(Kp_23__N_1402), .I2(n44585), 
            .I3(n48413), .O(n48427));
    defparam i1_4_lut_adj_1036.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1037 (.I0(n26857), .I1(n48423), .I2(n26890), 
            .I3(n26749), .O(n48433));
    defparam i1_4_lut_adj_1037.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1038 (.I0(n44645), .I1(n48427), .I2(n44624), 
            .I3(n44324), .O(n48435));
    defparam i1_4_lut_adj_1038.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1039 (.I0(n44757), .I1(n41445), .I2(n44353), 
            .I3(n27425), .O(n26));
    defparam i10_4_lut_adj_1039.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1040 (.I0(n44766), .I1(n28), .I2(n22_adj_4246), 
            .I3(n44677), .O(n30_adj_4247));
    defparam i14_4_lut_adj_1040.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1041 (.I0(n44357), .I1(n44668), .I2(n48435), 
            .I3(n48433), .O(n48441));
    defparam i1_4_lut_adj_1041.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1042 (.I0(\data_in_frame[11] [7]), .I1(n44603), 
            .I2(\data_in_frame[11] [0]), .I3(\data_in_frame[9] [6]), .O(n25));
    defparam i9_4_lut_adj_1042.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1043 (.I0(\data_in_frame[17] [1]), .I1(\data_in_frame[10] [3]), 
            .I2(\data_in_frame[14] [7]), .I3(GND_net), .O(n48379));
    defparam i1_3_lut_adj_1043.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1044 (.I0(n44769), .I1(n44763), .I2(Kp_23__N_1398), 
            .I3(n48379), .O(n48385));
    defparam i1_4_lut_adj_1044.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1045 (.I0(n44680), .I1(n44474), .I2(n48385), 
            .I3(n42126), .O(n48391));
    defparam i1_4_lut_adj_1045.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1046 (.I0(n44483), .I1(n44745), .I2(n48391), 
            .I3(n44656), .O(n48395));
    defparam i1_4_lut_adj_1046.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1047 (.I0(n25), .I1(n48441), .I2(n30_adj_4247), 
            .I3(n26), .O(n48443));
    defparam i1_4_lut_adj_1047.LUT_INIT = 16'h9669;
    SB_LUT4 i33987_4_lut (.I0(n48938), .I1(byte_transmit_counter[1]), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n48939));
    defparam i33987_4_lut.LUT_INIT = 16'haca3;
    SB_LUT4 i33985_3_lut (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[5] [4]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48937));
    defparam i33985_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_4_lut_adj_1048 (.I0(n48395), .I1(n44500), .I2(Kp_23__N_1653), 
            .I3(n44691), .O(n48399));
    defparam i1_4_lut_adj_1048.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1049 (.I0(n48399), .I1(n45717), .I2(n41435), 
            .I3(n48443), .O(n42291));
    defparam i1_4_lut_adj_1049.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_adj_1050 (.I0(n44715), .I1(n44585), .I2(\data_in_frame[11] [4]), 
            .I3(GND_net), .O(n48367));
    defparam i1_3_lut_adj_1050.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1051 (.I0(n42281), .I1(n42291), .I2(n44230), 
            .I3(n48367), .O(n42322));
    defparam i1_4_lut_adj_1051.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1052 (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [0]), 
            .I2(n1168), .I3(n44151), .O(n27558));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_4_lut_adj_1052.LUT_INIT = 16'h6996;
    SB_LUT4 i35048_2_lut (.I0(n51558), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n49805));
    defparam i35048_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_4_lut_adj_1053 (.I0(n42407), .I1(n44129), .I2(n27178), 
            .I3(n42444), .O(n45628));
    defparam i2_3_lut_4_lut_adj_1053.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1054 (.I0(n42407), .I1(n44129), .I2(\data_out_frame[24] [4]), 
            .I3(n44390), .O(n46698));
    defparam i2_3_lut_4_lut_adj_1054.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1055 (.I0(n42418), .I1(Kp_23__N_1644), .I2(n44378), 
            .I3(Kp_23__N_761), .O(n48523));
    defparam i1_4_lut_adj_1055.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i1 (.Q(\data_in_frame[0] [0]), .C(CLK_c), .D(n28212));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15259_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44085), .I2(rx_data[1]), 
            .I3(\data_in_frame[21] [1]), .O(n28322));
    defparam i15259_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_4_lut_adj_1056 (.I0(n42374), .I1(n42322), .I2(Kp_23__N_1653), 
            .I3(n48523), .O(n44418));
    defparam i1_4_lut_adj_1056.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1057 (.I0(\data_out_frame[4] [5]), .I1(\data_out_frame[5] [0]), 
            .I2(n1168), .I3(\data_out_frame[6] [7]), .O(n44712));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_4_lut_adj_1057.LUT_INIT = 16'h6996;
    SB_DFF neopxl_color_i0_i0 (.Q(neopxl_color[0]), .C(CLK_c), .D(n28211));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 data_in_frame_17__7__I_0_3899_2_lut (.I0(\data_in_frame[17] [7]), 
            .I1(\data_in_frame[17] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1398));   // verilog/coms.v(70[16:27])
    defparam data_in_frame_17__7__I_0_3899_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i15260_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44085), .I2(rx_data[0]), 
            .I3(\data_in_frame[21] [0]), .O(n28323));
    defparam i15260_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15313_3_lut_4_lut (.I0(n8_adj_4232), .I1(n44095), .I2(rx_data[3]), 
            .I3(\data_in_frame[14] [3]), .O(n28376));
    defparam i15313_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15258_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44085), .I2(rx_data[2]), 
            .I3(\data_in_frame[21] [2]), .O(n28321));
    defparam i15258_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_adj_1058 (.I0(n41723), .I1(n27312), .I2(\data_in_frame[13] [6]), 
            .I3(GND_net), .O(n44715));
    defparam i2_3_lut_adj_1058.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1059 (.I0(n44715), .I1(n41435), .I2(n44403), 
            .I3(n48653), .O(n46232));
    defparam i1_4_lut_adj_1059.LUT_INIT = 16'h6996;
    SB_LUT4 i15314_3_lut_4_lut (.I0(n8_adj_4232), .I1(n44095), .I2(rx_data[2]), 
            .I3(\data_in_frame[14] [2]), .O(n28377));
    defparam i15314_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15253_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44085), .I2(rx_data[7]), 
            .I3(\data_in_frame[21] [7]), .O(n28316));
    defparam i15253_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF Ki_i0 (.Q(\Ki[0] ), .C(CLK_c), .D(n28210));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i0 (.Q(\Kp[0] ), .C(CLK_c), .D(n28209));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i15315_3_lut_4_lut (.I0(n8_adj_4232), .I1(n44095), .I2(rx_data[1]), 
            .I3(\data_in_frame[14] [1]), .O(n28378));
    defparam i15315_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_DFF data_in_0___i1 (.Q(\data_in[0] [0]), .C(CLK_c), .D(n28208));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1060 (.I0(n44230), .I1(n44549), .I2(n46390), 
            .I3(n6_adj_4248), .O(n44659));   // verilog/coms.v(74[16:43])
    defparam i4_4_lut_adj_1060.LUT_INIT = 16'h9669;
    SB_LUT4 i15254_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44085), .I2(rx_data[6]), 
            .I3(\data_in_frame[21] [6]), .O(n28317));
    defparam i15254_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15255_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44085), .I2(rx_data[5]), 
            .I3(\data_in_frame[21] [5]), .O(n28318));
    defparam i15255_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1061 (.I0(\data_in_frame[19] [7]), .I1(\data_in_frame[19] [1]), 
            .I2(\data_in_frame[19] [2]), .I3(\data_in_frame[19] [3]), .O(n8_adj_4249));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_1061.LUT_INIT = 16'h6996;
    SB_LUT4 i15256_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44085), .I2(rx_data[4]), 
            .I3(\data_in_frame[21] [4]), .O(n28319));
    defparam i15256_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15257_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44085), .I2(rx_data[3]), 
            .I3(\data_in_frame[21] [3]), .O(n28320));
    defparam i15257_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_136_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4177));   // verilog/coms.v(154[7:23])
    defparam equal_136_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 equal_137_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4175));   // verilog/coms.v(154[7:23])
    defparam equal_137_i8_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(byte_transmit_counter[1]), .I2(n48915), .I3(n48913), .O(n7_adj_4239));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_0_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(byte_transmit_counter[1]), .I2(n48957), .I3(n48955), .O(n7_adj_4238));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_7_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i4_4_lut_adj_1062 (.I0(\data_in_frame[19] [6]), .I1(n8_adj_4249), 
            .I2(\data_in_frame[19] [4]), .I3(\data_in_frame[19] [5]), .O(Kp_23__N_761));   // verilog/coms.v(85[17:28])
    defparam i4_4_lut_adj_1062.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(byte_transmit_counter[1]), .I2(n48951), .I3(n48949), .O(n7_adj_4237));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_adj_1063 (.I0(n27347), .I1(n27606), .I2(GND_net), 
            .I3(GND_net), .O(n44671));
    defparam i1_2_lut_adj_1063.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1064 (.I0(n41580), .I1(n44448), .I2(n44671), 
            .I3(\data_in_frame[9] [3]), .O(n45717));
    defparam i1_4_lut_adj_1064.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1065 (.I0(\data_in_frame[10] [6]), .I1(n42354), 
            .I2(GND_net), .I3(GND_net), .O(n44652));
    defparam i1_2_lut_adj_1065.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1066 (.I0(n45717), .I1(\data_in_frame[13] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44406));
    defparam i1_2_lut_adj_1066.LUT_INIT = 16'h9999;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(byte_transmit_counter[1]), .I2(n48945), .I3(n48943), .O(n7_adj_4236));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_4_lut_adj_1067 (.I0(n4_adj_4250), .I1(n44742), .I2(\data_in_frame[13] [2]), 
            .I3(\data_in_frame[15] [4]), .O(n48559));
    defparam i1_4_lut_adj_1067.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1068 (.I0(n44406), .I1(n44652), .I2(Kp_23__N_1095), 
            .I3(n48559), .O(n46390));
    defparam i1_4_lut_adj_1068.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1069 (.I0(\data_in_frame[13] [1]), .I1(n44652), 
            .I2(n44527), .I3(\data_in_frame[17] [5]), .O(n44745));
    defparam i3_4_lut_adj_1069.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_adj_1070 (.I0(n44745), .I1(n46390), .I2(\data_in_frame[10] [5]), 
            .I3(GND_net), .O(n42281));
    defparam i1_3_lut_adj_1070.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1071 (.I0(n42281), .I1(n46677), .I2(GND_net), 
            .I3(GND_net), .O(n42374));
    defparam i1_2_lut_adj_1071.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1072 (.I0(n46677), .I1(n27459), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1653));
    defparam i1_2_lut_adj_1072.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_adj_1073 (.I0(n41956), .I1(n41474), .I2(GND_net), 
            .I3(GND_net), .O(n44515));
    defparam i1_2_lut_adj_1073.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(byte_transmit_counter[1]), .I2(n48939), .I3(n48937), .O(n7_adj_4235));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_2_lut_adj_1074 (.I0(\data_in_frame[10] [7]), .I1(\data_in_frame[11] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44677));
    defparam i1_2_lut_adj_1074.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1075 (.I0(\data_out_frame[13] [7]), .I1(\data_out_frame[13] [6]), 
            .I2(n42346), .I3(n50676), .O(n44497));
    defparam i1_2_lut_3_lut_4_lut_adj_1075.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1076 (.I0(n44458), .I1(n27023), .I2(n48461), 
            .I3(n44515), .O(n44448));
    defparam i1_4_lut_adj_1076.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1077 (.I0(n1699), .I1(n42346), .I2(n42427), 
            .I3(n44503), .O(n42350));
    defparam i2_3_lut_4_lut_adj_1077.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1078 (.I0(\data_in_frame[13] [2]), .I1(\data_in_frame[15] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44754));
    defparam i1_2_lut_adj_1078.LUT_INIT = 16'h6666;
    SB_DFF IntegralLimit_i0_i1 (.Q(IntegralLimit[1]), .C(CLK_c), .D(n28759));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i2 (.Q(IntegralLimit[2]), .C(CLK_c), .D(n28758));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_4_lut_adj_1079 (.I0(n41723), .I1(n44448), .I2(Kp_23__N_1221), 
            .I3(n27597), .O(n42354));
    defparam i1_4_lut_adj_1079.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(byte_transmit_counter[1]), .I2(n48933), .I3(n48931), .O(n7_adj_4234));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_3_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_4_lut_adj_1080 (.I0(Kp_23__N_1095), .I1(n44327), .I2(\data_in_frame[13] [0]), 
            .I3(\data_in_frame[17] [4]), .O(n48647));
    defparam i1_4_lut_adj_1080.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1081 (.I0(n44527), .I1(n42354), .I2(n44353), 
            .I3(n48647), .O(n46677));
    defparam i1_4_lut_adj_1081.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1082 (.I0(\data_in_frame[16] [4]), .I1(n41494), 
            .I2(GND_net), .I3(GND_net), .O(n42442));
    defparam i1_2_lut_adj_1082.LUT_INIT = 16'h6666;
    SB_DFF IntegralLimit_i0_i3 (.Q(IntegralLimit[3]), .C(CLK_c), .D(n28757));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i4 (.Q(IntegralLimit[4]), .C(CLK_c), .D(n28756));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i5 (.Q(IntegralLimit[5]), .C(CLK_c), .D(n28755));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i6 (.Q(IntegralLimit[6]), .C(CLK_c), .D(n28754));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i7 (.Q(IntegralLimit[7]), .C(CLK_c), .D(n28753));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i8 (.Q(IntegralLimit[8]), .C(CLK_c), .D(n28752));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i9 (.Q(IntegralLimit[9]), .C(CLK_c), .D(n28751));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i10 (.Q(IntegralLimit[10]), .C(CLK_c), .D(n28750));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i11 (.Q(IntegralLimit[11]), .C(CLK_c), .D(n28749));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i12 (.Q(IntegralLimit[12]), .C(CLK_c), .D(n28748));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i13 (.Q(IntegralLimit[13]), .C(CLK_c), .D(n28747));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i14 (.Q(IntegralLimit[14]), .C(CLK_c), .D(n28746));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i15 (.Q(IntegralLimit[15]), .C(CLK_c), .D(n28745));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i16 (.Q(IntegralLimit[16]), .C(CLK_c), .D(n28744));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i17 (.Q(IntegralLimit[17]), .C(CLK_c), .D(n28743));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i18 (.Q(IntegralLimit[18]), .C(CLK_c), .D(n28742));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i19 (.Q(IntegralLimit[19]), .C(CLK_c), .D(n28741));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i20 (.Q(IntegralLimit[20]), .C(CLK_c), .D(n28740));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i21 (.Q(IntegralLimit[21]), .C(CLK_c), .D(n28739));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i22 (.Q(IntegralLimit[22]), .C(CLK_c), .D(n28738));   // verilog/coms.v(127[12] 300[6])
    SB_DFF IntegralLimit_i0_i23 (.Q(IntegralLimit[23]), .C(CLK_c), .D(n28737));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i2 (.Q(\data_in[0] [1]), .C(CLK_c), .D(n28736));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i3 (.Q(\data_in[0] [2]), .C(CLK_c), .D(n28735));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i4 (.Q(\data_in[0] [3]), .C(CLK_c), .D(n28734));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i5 (.Q(\data_in[0] [4]), .C(CLK_c), .D(n28733));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i6 (.Q(\data_in[0] [5]), .C(CLK_c), .D(n28732));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i7 (.Q(\data_in[0] [6]), .C(CLK_c), .D(n28731));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i8 (.Q(\data_in[0] [7]), .C(CLK_c), .D(n28730));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i9 (.Q(\data_in[1] [0]), .C(CLK_c), .D(n28729));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i10 (.Q(\data_in[1] [1]), .C(CLK_c), .D(n28728));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i11 (.Q(\data_in[1] [2]), .C(CLK_c), .D(n28727));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_4_lut_adj_1083 (.I0(\data_in_frame[11] [6]), .I1(\data_in_frame[9] [6]), 
            .I2(n41956), .I3(\data_in_frame[9] [5]), .O(n44757));
    defparam i1_4_lut_adj_1083.LUT_INIT = 16'h9669;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(byte_transmit_counter[1]), .I2(n48918), .I3(n48916), .O(n7_adj_4231));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_1_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i1_4_lut_adj_1084 (.I0(n44591), .I1(\data_in_frame[5] [0]), 
            .I2(\data_in_frame[6] [0]), .I3(\data_in_frame[10] [0]), .O(n48593));
    defparam i1_4_lut_adj_1084.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1085 (.I0(n48593), .I1(n26978), .I2(n44154), 
            .I3(n44706), .O(n48599));
    defparam i1_4_lut_adj_1085.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1086 (.I0(n44567), .I1(n44282), .I2(n44639), 
            .I3(n48603), .O(n48609));
    defparam i1_4_lut_adj_1086.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1087 (.I0(n44512), .I1(n44757), .I2(n42348), 
            .I3(n48609), .O(n41494));
    defparam i1_4_lut_adj_1087.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1088 (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[16] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44521));
    defparam i1_2_lut_adj_1088.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1089 (.I0(n44521), .I1(\data_in_frame[11] [4]), 
            .I2(\data_in_frame[9] [3]), .I3(\data_in_frame[14] [2]), .O(n48577));   // verilog/coms.v(75[16:43])
    defparam i1_4_lut_adj_1089.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1090 (.I0(n27587), .I1(Kp_23__N_1233), .I2(n48577), 
            .I3(n44718), .O(n48583));   // verilog/coms.v(75[16:43])
    defparam i1_4_lut_adj_1090.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1091 (.I0(\data_in_frame[18] [4]), .I1(n27347), 
            .I2(n41494), .I3(n48583), .O(n44691));
    defparam i1_4_lut_adj_1091.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_adj_1092 (.I0(n44246), .I1(n42367), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4251));
    defparam i2_2_lut_adj_1092.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1093 (.I0(\data_in_frame[18] [5]), .I1(\data_in_frame[16] [4]), 
            .I2(n6_adj_4251), .I3(\data_in_frame[16] [3]), .O(n44500));
    defparam i1_4_lut_adj_1093.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1094 (.I0(\data_in_frame[9] [0]), .I1(\data_in_frame[11] [2]), 
            .I2(Kp_23__N_1095), .I3(GND_net), .O(n44603));   // verilog/coms.v(72[16:41])
    defparam i2_3_lut_adj_1094.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1095 (.I0(\data_in_frame[4] [5]), .I1(n27337), 
            .I2(n44363), .I3(\data_in_frame[1] [7]), .O(n44360));
    defparam i1_2_lut_4_lut_adj_1095.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1096 (.I0(n27650), .I1(\data_in_frame[8] [2]), 
            .I2(Kp_23__N_1095), .I3(n44760), .O(n20_adj_4252));   // verilog/coms.v(78[16:27])
    defparam i8_4_lut_adj_1096.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut (.I0(\byte_transmit_counter[2] ), 
            .I1(byte_transmit_counter[1]), .I2(n48927), .I3(n48925), .O(n7_adj_4233));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_2_i7_3_lut_4_lut.LUT_INIT = 16'hf2d0;
    SB_LUT4 i7_4_lut_adj_1097 (.I0(n41956), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[12] [0]), .I3(n44730), .O(n19_adj_4253));   // verilog/coms.v(78[16:27])
    defparam i7_4_lut_adj_1097.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1098 (.I0(n34355), .I1(n34549), .I2(n34685), 
            .I3(n34047), .O(n34823));   // verilog/coms.v(231[5:23])
    defparam i2_3_lut_4_lut_adj_1098.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut_adj_1099 (.I0(n44615), .I1(\data_in_frame[8] [4]), 
            .I2(\data_in_frame[6] [3]), .I3(\data_in_frame[8] [3]), .O(n21));   // verilog/coms.v(78[16:27])
    defparam i9_4_lut_adj_1099.LUT_INIT = 16'h6996;
    SB_LUT4 i11_3_lut_adj_1100 (.I0(n21), .I1(n19_adj_4253), .I2(n20_adj_4252), 
            .I3(GND_net), .O(n44512));   // verilog/coms.v(78[16:27])
    defparam i11_3_lut_adj_1100.LUT_INIT = 16'h9696;
    SB_LUT4 i2_2_lut_3_lut_adj_1101 (.I0(n34355), .I1(n34549), .I2(n34685), 
            .I3(GND_net), .O(n33298));   // verilog/coms.v(231[5:23])
    defparam i2_2_lut_3_lut_adj_1101.LUT_INIT = 16'hfefe;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36560 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [7]), .I2(\data_out_frame[19] [7]), 
            .I3(byte_transmit_counter[1]), .O(n51453));
    defparam byte_transmit_counter_0__bdd_4_lut_36560.LUT_INIT = 16'he4aa;
    SB_LUT4 i30057_2_lut_3_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state_c [2]), 
            .I2(n44929), .I3(GND_net), .O(n44947));
    defparam i30057_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i7_4_lut_adj_1102 (.I0(n44512), .I1(\data_in_frame[11] [7]), 
            .I2(\data_in_frame[9] [1]), .I3(n41449), .O(n18_adj_4254));
    defparam i7_4_lut_adj_1102.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut (.I0(n44170), .I1(\data_in_frame[9] [7]), .I2(GND_net), 
            .I3(GND_net), .O(n16_adj_4255));
    defparam i5_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1103 (.I0(\data_in_frame[11] [5]), .I1(n18_adj_4254), 
            .I2(\data_in_frame[14] [1]), .I3(\data_in_frame[9] [0]), .O(n20_adj_4256));
    defparam i9_4_lut_adj_1103.LUT_INIT = 16'h6996;
    SB_LUT4 i10_4_lut_adj_1104 (.I0(n44553), .I1(n20_adj_4256), .I2(n16_adj_4255), 
            .I3(\data_in_frame[13] [7]), .O(n44246));
    defparam i10_4_lut_adj_1104.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1105 (.I0(\data_in_frame[6] [7]), .I1(n26834), 
            .I2(n27356), .I3(\data_in_frame[4] [4]), .O(n44294));   // verilog/coms.v(236[9:81])
    defparam i1_2_lut_4_lut_adj_1105.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1106 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state_c [2]), 
            .I2(\FRAME_MATCHER.state_c [1]), .I3(GND_net), .O(n34047));
    defparam i2_2_lut_3_lut_adj_1106.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut_adj_1107 (.I0(\data_in_frame[15] [7]), .I1(n44648), 
            .I2(GND_net), .I3(GND_net), .O(n44739));
    defparam i1_2_lut_adj_1107.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1108 (.I0(\data_in_frame[13] [6]), .I1(\data_in_frame[14] [0]), 
            .I2(\data_in_frame[13] [7]), .I3(GND_net), .O(n44718));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1108.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1109 (.I0(n41445), .I1(n27414), .I2(GND_net), 
            .I3(GND_net), .O(n41449));
    defparam i1_2_lut_adj_1109.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1110 (.I0(\data_in_frame[16] [0]), .I1(n44549), 
            .I2(GND_net), .I3(GND_net), .O(n44403));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1110.LUT_INIT = 16'h6666;
    SB_LUT4 i3_4_lut_adj_1111 (.I0(\data_in_frame[11] [6]), .I1(n42295), 
            .I2(n41580), .I3(\data_in_frame[9] [5]), .O(n27587));
    defparam i3_4_lut_adj_1111.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1112 (.I0(\data_in_frame[15] [6]), .I1(n44718), 
            .I2(\data_in_frame[16] [1]), .I3(GND_net), .O(n44645));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_adj_1112.LUT_INIT = 16'h9696;
    SB_LUT4 i5_4_lut_adj_1113 (.I0(n27606), .I1(n44645), .I2(\data_in_frame[9] [1]), 
            .I3(\data_in_frame[13] [4]), .O(n12_adj_4257));   // verilog/coms.v(70[16:27])
    defparam i5_4_lut_adj_1113.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1114 (.I0(n27587), .I1(n12_adj_4257), .I2(\data_in_frame[18] [2]), 
            .I3(n44403), .O(n44656));   // verilog/coms.v(70[16:27])
    defparam i6_4_lut_adj_1114.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1115 (.I0(n27347), .I1(\data_in_frame[16] [1]), 
            .I2(n44246), .I3(GND_net), .O(n10_adj_4258));
    defparam i2_3_lut_adj_1115.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1116 (.I0(n44739), .I1(n41580), .I2(n44549), 
            .I3(\data_in_frame[11] [5]), .O(n14_adj_4259));
    defparam i6_4_lut_adj_1116.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1117 (.I0(\data_in_frame[16] [2]), .I1(\data_in_frame[13] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n9_adj_4260));
    defparam i1_2_lut_adj_1117.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1118 (.I0(\data_in_frame[18] [3]), .I1(n9_adj_4260), 
            .I2(n14_adj_4259), .I3(n10_adj_4258), .O(n44483));
    defparam i1_4_lut_adj_1118.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1119 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[12] [1]), 
            .I2(n41445), .I3(GND_net), .O(n44567));
    defparam i2_3_lut_adj_1119.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1120 (.I0(\data_in_frame[9] [2]), .I1(\data_in_frame[9] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44154));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1120.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1121 (.I0(\data_in_frame[2] [3]), .I1(\data_in_frame[0] [2]), 
            .I2(\data_in_frame[0] [1]), .I3(GND_net), .O(n27337));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1121.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_4_lut_adj_1122 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[5] [6]), .O(n48477));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_4_lut_adj_1122.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1123 (.I0(\data_in_frame[2] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[0] [3]), .I3(GND_net), .O(n26770));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1123.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1124 (.I0(n27650), .I1(n44627), .I2(n44736), 
            .I3(GND_net), .O(n44766));
    defparam i1_3_lut_adj_1124.LUT_INIT = 16'h6969;
    SB_LUT4 i1_2_lut_adj_1125 (.I0(n27411), .I1(n27414), .I2(GND_net), 
            .I3(GND_net), .O(Kp_23__N_1233));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1125.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1126 (.I0(n26746), .I1(n44766), .I2(n27010), 
            .I3(n48447), .O(n44458));
    defparam i1_4_lut_adj_1126.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1127 (.I0(n41445), .I1(n27023), .I2(GND_net), 
            .I3(GND_net), .O(n42295));
    defparam i1_2_lut_adj_1127.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1128 (.I0(\data_in_frame[3] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[1] [2]), .I3(GND_net), .O(n27063));
    defparam i1_2_lut_3_lut_adj_1128.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1129 (.I0(n26834), .I1(\data_in_frame[2] [3]), 
            .I2(n44142), .I3(\data_in_frame[4] [5]), .O(n27584));   // verilog/coms.v(75[16:43])
    defparam i1_3_lut_4_lut_adj_1129.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1130 (.I0(n27425), .I1(n42348), .I2(n27597), 
            .I3(\data_in_frame[9] [0]), .O(n44207));
    defparam i1_4_lut_adj_1130.LUT_INIT = 16'h9669;
    SB_LUT4 i6_2_lut_3_lut_4_lut (.I0(\data_in_frame[11] [4]), .I1(n44648), 
            .I2(n41956), .I3(n41474), .O(n22_adj_4246));   // verilog/coms.v(74[16:43])
    defparam i6_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1131 (.I0(\data_in_frame[12] [2]), .I1(\data_in_frame[11] [7]), 
            .I2(n44567), .I3(n44207), .O(n14_adj_4261));
    defparam i6_4_lut_adj_1131.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1132 (.I0(\data_in_frame[14] [3]), .I1(n14_adj_4261), 
            .I2(n10_adj_4262), .I3(n41956), .O(n42367));
    defparam i7_4_lut_adj_1132.LUT_INIT = 16'h6996;
    SB_DFF data_in_0___i12 (.Q(\data_in[1] [3]), .C(CLK_c), .D(n28726));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i13 (.Q(\data_in[1] [4]), .C(CLK_c), .D(n28725));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i14 (.Q(\data_in[1] [5]), .C(CLK_c), .D(n28724));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i15 (.Q(\data_in[1] [6]), .C(CLK_c), .D(n28723));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i16 (.Q(\data_in[1] [7]), .C(CLK_c), .D(n28722));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i17 (.Q(\data_in[2] [0]), .C(CLK_c), .D(n28721));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i18 (.Q(\data_in[2] [1]), .C(CLK_c), .D(n28720));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i19 (.Q(\data_in[2] [2]), .C(CLK_c), .D(n28719));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i20 (.Q(\data_in[2] [3]), .C(CLK_c), .D(n28718));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i21 (.Q(\data_in[2] [4]), .C(CLK_c), .D(n28717));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1133 (.I0(\data_in_frame[10] [1]), .I1(\data_in_frame[10] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n26854));
    defparam i1_2_lut_adj_1133.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1134 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [3]), 
            .I2(n44243), .I3(n27360), .O(n48351));   // verilog/coms.v(166[9:87])
    defparam i1_3_lut_4_lut_adj_1134.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1135 (.I0(n25051), .I1(n42367), .I2(GND_net), 
            .I3(GND_net), .O(n44474));
    defparam i1_2_lut_adj_1135.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_3_lut_adj_1136 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [3]), 
            .I2(\data_in_frame[2] [4]), .I3(GND_net), .O(n26834));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_3_lut_adj_1136.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1137 (.I0(\data_in_frame[16] [6]), .I1(n45701), 
            .I2(n44474), .I3(n26854), .O(n44636));
    defparam i3_4_lut_adj_1137.LUT_INIT = 16'h9669;
    SB_LUT4 i3_4_lut_adj_1138 (.I0(\data_in_frame[18] [7]), .I1(n44636), 
            .I2(n44348), .I3(\data_in_frame[16] [5]), .O(n42418));
    defparam i3_4_lut_adj_1138.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1139 (.I0(n27010), .I1(n27023), .I2(GND_net), 
            .I3(GND_net), .O(n44553));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1139.LUT_INIT = 16'h6666;
    SB_LUT4 i15316_3_lut_4_lut (.I0(n8_adj_4232), .I1(n44095), .I2(rx_data[0]), 
            .I3(\data_in_frame[14] [0]), .O(n28379));
    defparam i15316_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1140 (.I0(n25836), .I1(\data_in_frame[2] [7]), 
            .I2(Kp_23__N_888), .I3(\data_in_frame[0] [7]), .O(n27198));
    defparam i2_3_lut_4_lut_adj_1140.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1141 (.I0(\data_in_frame[9] [7]), .I1(\data_in_frame[9] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44148));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1141.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1142 (.I0(\data_in_frame[14] [4]), .I1(\data_in_frame[12] [2]), 
            .I2(\data_in_frame[12] [3]), .I3(GND_net), .O(n44324));
    defparam i2_3_lut_adj_1142.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1143 (.I0(\data_in_frame[10] [0]), .I1(n44148), 
            .I2(\data_in_frame[10] [2]), .I3(n44553), .O(n41447));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_1143.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1144 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[5] [1]), .I3(\data_out_frame[5] [2]), .O(n44573));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_4_lut_adj_1144.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1145 (.I0(n41447), .I1(n44324), .I2(n41451), 
            .I3(GND_net), .O(n27297));
    defparam i2_3_lut_adj_1145.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1146 (.I0(n44464), .I1(\data_in_frame[14] [5]), 
            .I2(n27297), .I3(GND_net), .O(n44348));
    defparam i2_3_lut_adj_1146.LUT_INIT = 16'h9696;
    SB_DFF data_in_0___i22 (.Q(\data_in[2] [5]), .C(CLK_c), .D(n28716));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i23 (.Q(\data_in[2] [6]), .C(CLK_c), .D(n28715));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i24 (.Q(\data_in[2] [7]), .C(CLK_c), .D(n28714));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i25 (.Q(\data_in[3] [0]), .C(CLK_c), .D(n28713));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i26 (.Q(\data_in[3] [1]), .C(CLK_c), .D(n28712));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i27 (.Q(\data_in[3] [2]), .C(CLK_c), .D(n28711));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i28 (.Q(\data_in[3] [3]), .C(CLK_c), .D(n28710));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i29 (.Q(\data_in[3] [4]), .C(CLK_c), .D(n28709));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i30 (.Q(\data_in[3] [5]), .C(CLK_c), .D(n28708));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i31 (.Q(\data_in[3] [6]), .C(CLK_c), .D(n28707));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_0___i32 (.Q(\data_in[3] [7]), .C(CLK_c), .D(n28706));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i1 (.Q(\Kp[1] ), .C(CLK_c), .D(n28705));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i2 (.Q(\Kp[2] ), .C(CLK_c), .D(n28704));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i3 (.Q(\Kp[3] ), .C(CLK_c), .D(n28703));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i4 (.Q(\Kp[4] ), .C(CLK_c), .D(n28702));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i5 (.Q(\Kp[5] ), .C(CLK_c), .D(n28701));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i6 (.Q(\Kp[6] ), .C(CLK_c), .D(n28700));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i7 (.Q(\Kp[7] ), .C(CLK_c), .D(n28699));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i8 (.Q(\Kp[8] ), .C(CLK_c), .D(n28698));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i9 (.Q(\Kp[9] ), .C(CLK_c), .D(n28697));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i10 (.Q(\Kp[10] ), .C(CLK_c), .D(n28696));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i11 (.Q(\Kp[11] ), .C(CLK_c), .D(n28695));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i12 (.Q(\Kp[12] ), .C(CLK_c), .D(n28694));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i13 (.Q(\Kp[13] ), .C(CLK_c), .D(n28693));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i14 (.Q(\Kp[14] ), .C(CLK_c), .D(n28692));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Kp_i15 (.Q(\Kp[15] ), .C(CLK_c), .D(n28691));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i1 (.Q(\Ki[1] ), .C(CLK_c), .D(n28690));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i2 (.Q(\Ki[2] ), .C(CLK_c), .D(n28689));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i3 (.Q(\Ki[3] ), .C(CLK_c), .D(n28688));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i4 (.Q(\Ki[4] ), .C(CLK_c), .D(n28687));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i5 (.Q(\Ki[5] ), .C(CLK_c), .D(n28686));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i6 (.Q(\Ki[6] ), .C(CLK_c), .D(n28685));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i7 (.Q(\Ki[7] ), .C(CLK_c), .D(n28684));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i8 (.Q(\Ki[8] ), .C(CLK_c), .D(n28683));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i9 (.Q(\Ki[9] ), .C(CLK_c), .D(n28682));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i10 (.Q(\Ki[10] ), .C(CLK_c), .D(n28681));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i11 (.Q(\Ki[11] ), .C(CLK_c), .D(n28680));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i12 (.Q(\Ki[12] ), .C(CLK_c), .D(n28679));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i13 (.Q(\Ki[13] ), .C(CLK_c), .D(n28678));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i14 (.Q(\Ki[14] ), .C(CLK_c), .D(n28677));   // verilog/coms.v(127[12] 300[6])
    SB_DFF Ki_i15 (.Q(\Ki[15] ), .C(CLK_c), .D(n28676));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i33 (.Q(\data_out_frame[4] [0]), .C(CLK_c), 
           .D(n28675));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i34 (.Q(\data_out_frame[4] [1]), .C(CLK_c), 
           .D(n28674));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i35 (.Q(\data_out_frame[4] [2]), .C(CLK_c), 
           .D(n28673));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i36 (.Q(\data_out_frame[4] [3]), .C(CLK_c), 
           .D(n28672));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i37 (.Q(\data_out_frame[4] [4]), .C(CLK_c), 
           .D(n28671));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i38 (.Q(\data_out_frame[4] [5]), .C(CLK_c), 
           .D(n28670));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i39 (.Q(\data_out_frame[4] [6]), .C(CLK_c), 
           .D(n28669));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i40 (.Q(\data_out_frame[4] [7]), .C(CLK_c), 
           .D(n28668));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i41 (.Q(\data_out_frame[5] [0]), .C(CLK_c), 
           .D(n28667));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i42 (.Q(\data_out_frame[5] [1]), .C(CLK_c), 
           .D(n28666));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i43 (.Q(\data_out_frame[5] [2]), .C(CLK_c), 
           .D(n28665));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i44 (.Q(\data_out_frame[5] [3]), .C(CLK_c), 
           .D(n28664));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i45 (.Q(\data_out_frame[5] [4]), .C(CLK_c), 
           .D(n28663));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i46 (.Q(\data_out_frame[5] [5]), .C(CLK_c), 
           .D(n28662));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i47 (.Q(\data_out_frame[5] [6]), .C(CLK_c), 
           .D(n28661));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i48 (.Q(\data_out_frame[5] [7]), .C(CLK_c), 
           .D(n28660));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i49 (.Q(\data_out_frame[6] [0]), .C(CLK_c), 
           .D(n28659));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i50 (.Q(\data_out_frame[6] [1]), .C(CLK_c), 
           .D(n28658));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i51 (.Q(\data_out_frame[6] [2]), .C(CLK_c), 
           .D(n28657));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i52 (.Q(\data_out_frame[6] [3]), .C(CLK_c), 
           .D(n28656));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i53 (.Q(\data_out_frame[6] [4]), .C(CLK_c), 
           .D(n28655));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i54 (.Q(\data_out_frame[6] [5]), .C(CLK_c), 
           .D(n28654));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i55 (.Q(\data_out_frame[6] [6]), .C(CLK_c), 
           .D(n28653));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i56 (.Q(\data_out_frame[6] [7]), .C(CLK_c), 
           .D(n28652));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i57 (.Q(\data_out_frame[7] [0]), .C(CLK_c), 
           .D(n28651));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i58 (.Q(\data_out_frame[7] [1]), .C(CLK_c), 
           .D(n28650));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i59 (.Q(\data_out_frame[7] [2]), .C(CLK_c), 
           .D(n28649));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i60 (.Q(\data_out_frame[7] [3]), .C(CLK_c), 
           .D(n28648));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i61 (.Q(\data_out_frame[7] [4]), .C(CLK_c), 
           .D(n28647));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i62 (.Q(\data_out_frame[7] [5]), .C(CLK_c), 
           .D(n28646));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i63 (.Q(\data_out_frame[7] [6]), .C(CLK_c), 
           .D(n28645));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i64 (.Q(\data_out_frame[7] [7]), .C(CLK_c), 
           .D(n28644));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i65 (.Q(\data_out_frame[8] [0]), .C(CLK_c), 
           .D(n28643));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i66 (.Q(\data_out_frame[8] [1]), .C(CLK_c), 
           .D(n28642));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i67 (.Q(\data_out_frame[8] [2]), .C(CLK_c), 
           .D(n28641));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i68 (.Q(\data_out_frame[8] [3]), .C(CLK_c), 
           .D(n28640));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i69 (.Q(\data_out_frame[8] [4]), .C(CLK_c), 
           .D(n28639));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1147 (.I0(\data_in_frame[8] [0]), .I1(\data_in_frame[7] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n44615));
    defparam i1_2_lut_adj_1147.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i70 (.Q(\data_out_frame[8] [5]), .C(CLK_c), 
           .D(n28638));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i71 (.Q(\data_out_frame[8] [6]), .C(CLK_c), 
           .D(n28637));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i72 (.Q(\data_out_frame[8] [7]), .C(CLK_c), 
           .D(n28636));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i73 (.Q(\data_out_frame[9] [0]), .C(CLK_c), 
           .D(n28635));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i74 (.Q(\data_out_frame[9] [1]), .C(CLK_c), 
           .D(n28634));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i75 (.Q(\data_out_frame[9] [2]), .C(CLK_c), 
           .D(n28633));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i76 (.Q(\data_out_frame[9] [3]), .C(CLK_c), 
           .D(n28632));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i77 (.Q(\data_out_frame[9] [4]), .C(CLK_c), 
           .D(n28631));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i78 (.Q(\data_out_frame[9] [5]), .C(CLK_c), 
           .D(n28630));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i79 (.Q(\data_out_frame[9] [6]), .C(CLK_c), 
           .D(n28629));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i80 (.Q(\data_out_frame[9] [7]), .C(CLK_c), 
           .D(n28628));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i81 (.Q(\data_out_frame[10] [0]), .C(CLK_c), 
           .D(n28627));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i82 (.Q(\data_out_frame[10] [1]), .C(CLK_c), 
           .D(n28626));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i83 (.Q(\data_out_frame[10] [2]), .C(CLK_c), 
           .D(n28625));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i84 (.Q(\data_out_frame[10] [3]), .C(CLK_c), 
           .D(n28624));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i85 (.Q(\data_out_frame[10] [4]), .C(CLK_c), 
           .D(n28623));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i86 (.Q(\data_out_frame[10] [5]), .C(CLK_c), 
           .D(n28622));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i87 (.Q(\data_out_frame[10] [6]), .C(CLK_c), 
           .D(n28621));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i88 (.Q(\data_out_frame[10] [7]), .C(CLK_c), 
           .D(n28620));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i89 (.Q(\data_out_frame[11] [0]), .C(CLK_c), 
           .D(n28619));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i90 (.Q(\data_out_frame[11] [1]), .C(CLK_c), 
           .D(n28618));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i91 (.Q(\data_out_frame[11] [2]), .C(CLK_c), 
           .D(n28617));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i92 (.Q(\data_out_frame[11] [3]), .C(CLK_c), 
           .D(n28616));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i93 (.Q(\data_out_frame[11] [4]), .C(CLK_c), 
           .D(n28615));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i94 (.Q(\data_out_frame[11] [5]), .C(CLK_c), 
           .D(n28614));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i95 (.Q(\data_out_frame[11] [6]), .C(CLK_c), 
           .D(n28613));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i96 (.Q(\data_out_frame[11] [7]), .C(CLK_c), 
           .D(n28612));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i97 (.Q(\data_out_frame[12] [0]), .C(CLK_c), 
           .D(n28611));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i98 (.Q(\data_out_frame[12] [1]), .C(CLK_c), 
           .D(n28610));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i99 (.Q(\data_out_frame[12] [2]), .C(CLK_c), 
           .D(n28609));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1148 (.I0(n44615), .I1(n44161), .I2(\data_in_frame[9] [7]), 
            .I3(n44642), .O(n10_adj_4263));
    defparam i4_4_lut_adj_1148.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_adj_1149 (.I0(n44307), .I1(n10_adj_4263), .I2(\data_in_frame[5] [5]), 
            .I3(GND_net), .O(n42133));
    defparam i5_3_lut_adj_1149.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1150 (.I0(\data_in_frame[11] [4]), .I1(n44648), 
            .I2(\data_in_frame[17] [7]), .I3(\data_in_frame[17] [6]), .O(n6_adj_4248));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1150.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1151 (.I0(\data_in_frame[12] [3]), .I1(n42133), 
            .I2(\data_in_frame[12] [4]), .I3(GND_net), .O(n45701));
    defparam i2_3_lut_adj_1151.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1152 (.I0(\data_out_frame[5] [7]), .I1(\data_out_frame[5] [6]), 
            .I2(\data_out_frame[10] [7]), .I3(\data_out_frame[10] [0]), 
            .O(n14_adj_4130));   // verilog/coms.v(71[16:27])
    defparam i5_3_lut_4_lut_adj_1152.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1153 (.I0(n25836), .I1(\data_in_frame[2] [7]), 
            .I2(\data_in_frame[7] [4]), .I3(n10_adj_4264), .O(n44282));
    defparam i5_3_lut_4_lut_adj_1153.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1154 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [7]), 
            .I2(n27356), .I3(GND_net), .O(n6_adj_4265));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1154.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1155 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[1] [7]), 
            .I2(\data_in_frame[1] [5]), .I3(GND_net), .O(n26866));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_3_lut_adj_1155.LUT_INIT = 16'h9696;
    SB_LUT4 i4_4_lut_adj_1156 (.I0(n45701), .I1(n26857), .I2(\data_in_frame[17] [1]), 
            .I3(n44439), .O(n10_adj_4266));
    defparam i4_4_lut_adj_1156.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1157 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(\data_in_frame[1] [4]), .I3(\data_in_frame[5] [6]), .O(n27660));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_4_lut_adj_1157.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1158 (.I0(\data_in_frame[5] [5]), .I1(n44674), 
            .I2(n27063), .I3(\data_in_frame[7] [6]), .O(n27010));
    defparam i2_3_lut_4_lut_adj_1158.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1159 (.I0(\FRAME_MATCHER.state_c [9]), .I1(\FRAME_MATCHER.state_c [8]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4267));
    defparam i2_2_lut_adj_1159.LUT_INIT = 16'heeee;
    SB_LUT4 i5_3_lut_adj_1160 (.I0(\data_in_frame[10] [1]), .I1(n10_adj_4266), 
            .I2(\data_in_frame[16] [7]), .I3(GND_net), .O(n44665));
    defparam i5_3_lut_adj_1160.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1161 (.I0(\data_in_frame[5] [5]), .I1(n44674), 
            .I2(n48361), .I3(n44251), .O(n41468));
    defparam i1_3_lut_4_lut_adj_1161.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1162 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[0] [7]), .I3(\data_in_frame[1] [6]), .O(n22_adj_4132));   // verilog/coms.v(70[16:27])
    defparam i5_3_lut_4_lut_adj_1162.LUT_INIT = 16'h9600;
    SB_LUT4 i2_3_lut_4_lut_adj_1163 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[3] [0]), .I3(Kp_23__N_888), .O(n27579));   // verilog/coms.v(70[16:27])
    defparam i2_3_lut_4_lut_adj_1163.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1164 (.I0(\data_in_frame[8] [6]), .I1(\data_in_frame[11] [0]), 
            .I2(\data_in_frame[10] [7]), .I3(GND_net), .O(n44742));
    defparam i2_3_lut_adj_1164.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1165 (.I0(\FRAME_MATCHER.state_c [10]), .I1(\FRAME_MATCHER.state_c [14]), 
            .I2(\FRAME_MATCHER.state_c [12]), .I3(\FRAME_MATCHER.state_c [15]), 
            .O(n14_adj_4268));
    defparam i6_4_lut_adj_1165.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1166 (.I0(Kp_23__N_1095), .I1(n27425), .I2(GND_net), 
            .I3(GND_net), .O(n26746));
    defparam i1_2_lut_adj_1166.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1167 (.I0(\data_in_frame[15] [2]), .I1(n44742), 
            .I2(\data_in_frame[12] [6]), .I3(GND_net), .O(n44327));
    defparam i2_3_lut_adj_1167.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1168 (.I0(\data_in_frame[0] [6]), .I1(\data_in_frame[1] [0]), 
            .I2(\data_in_frame[3] [2]), .I3(\data_in_frame[1] [1]), .O(n44454));   // verilog/coms.v(70[16:27])
    defparam i1_3_lut_4_lut_adj_1168.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1169 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[3] [5]), .I3(GND_net), .O(n44234));   // verilog/coms.v(75[16:27])
    defparam i1_2_lut_3_lut_adj_1169.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1170 (.I0(\data_in_frame[8] [1]), .I1(n27530), 
            .I2(GND_net), .I3(GND_net), .O(n44730));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1170.LUT_INIT = 16'h6666;
    SB_LUT4 i1_3_lut_4_lut_adj_1171 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[1] [3]), 
            .I2(\data_in_frame[3] [5]), .I3(\data_in_frame[3] [7]), .O(n44556));   // verilog/coms.v(78[16:27])
    defparam i1_3_lut_4_lut_adj_1171.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1172 (.I0(n26966), .I1(n27411), .I2(n41445), 
            .I3(n27414), .O(n41723));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_3_lut_4_lut_adj_1172.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1173 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[1] [3]), 
            .I2(n10_adj_4269), .I3(n44301), .O(n25051));   // verilog/coms.v(75[16:27])
    defparam i5_3_lut_4_lut_adj_1173.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1174 (.I0(n26996), .I1(n27425), .I2(\data_in_frame[12] [7]), 
            .I3(GND_net), .O(n44751));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1174.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1175 (.I0(\data_in_frame[13] [0]), .I1(n44439), 
            .I2(\data_in_frame[12] [4]), .I3(\data_in_frame[14] [6]), .O(n44668));
    defparam i1_2_lut_3_lut_4_lut_adj_1175.LUT_INIT = 16'h6996;
    SB_LUT4 i5_3_lut_4_lut_adj_1176 (.I0(\data_in_frame[1] [1]), .I1(n44310), 
            .I2(\data_in_frame[7] [6]), .I3(n10_adj_4270), .O(n41451));   // verilog/coms.v(73[16:34])
    defparam i5_3_lut_4_lut_adj_1176.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1177 (.I0(\data_in_frame[1] [1]), .I1(n44310), 
            .I2(n27063), .I3(\data_in_frame[5] [5]), .O(n27530));   // verilog/coms.v(73[16:34])
    defparam i2_3_lut_4_lut_adj_1177.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1178 (.I0(n44339), .I1(\data_in_frame[1] [2]), 
            .I2(\data_in_frame[3] [4]), .I3(n44627), .O(n10_adj_4269));
    defparam i4_4_lut_adj_1178.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1179 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(n44282), .I3(\data_in_frame[2] [6]), .O(n27023));
    defparam i2_3_lut_4_lut_adj_1179.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1180 (.I0(\data_in_frame[2] [6]), .I1(Kp_23__N_881), 
            .I2(n26770), .I3(\data_in_frame[5] [0]), .O(n44594));
    defparam i1_2_lut_4_lut_adj_1180.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1181 (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[12] [7]), 
            .I2(\data_in_frame[13] [1]), .I3(GND_net), .O(n44624));
    defparam i2_3_lut_adj_1181.LUT_INIT = 16'h9696;
    SB_LUT4 i5_3_lut_4_lut_adj_1182 (.I0(\data_in_frame[4] [6]), .I1(n10_adj_4271), 
            .I2(\data_in_frame[2] [3]), .I3(n44142), .O(n26966));   // verilog/coms.v(236[9:81])
    defparam i5_3_lut_4_lut_adj_1182.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i100 (.Q(\data_out_frame[12] [3]), .C(CLK_c), 
           .D(n28608));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_4_lut_adj_1183 (.I0(n44327), .I1(n7_adj_4272), .I2(n26746), 
            .I3(n8_adj_4273), .O(n27459));
    defparam i5_4_lut_adj_1183.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1184 (.I0(\data_in_frame[1] [1]), .I1(n44310), 
            .I2(n44307), .I3(GND_net), .O(n41474));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_3_lut_adj_1184.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1185 (.I0(\data_in_frame[8] [5]), .I1(n44760), 
            .I2(n48599), .I3(n26770), .O(n48603));   // verilog/coms.v(75[16:43])
    defparam i1_3_lut_4_lut_adj_1185.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1186 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[8] [2]), 
            .I2(\data_out_frame[10] [3]), .I3(\data_out_frame[10] [2]), 
            .O(n44582));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut_adj_1186.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1187 (.I0(\data_in_frame[8] [5]), .I1(n44760), 
            .I2(\data_in_frame[6] [3]), .I3(n44345), .O(n27425));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1187.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1188 (.I0(n44227), .I1(n44668), .I2(\data_in_frame[17] [2]), 
            .I3(\data_in_frame[10] [6]), .O(n12_adj_4274));
    defparam i5_4_lut_adj_1188.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1189 (.I0(\data_in_frame[15] [1]), .I1(n12_adj_4274), 
            .I2(n44751), .I3(\data_in_frame[12] [5]), .O(n42126));
    defparam i6_4_lut_adj_1189.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1190 (.I0(\data_in_frame[14] [5]), .I1(n44665), 
            .I2(n42126), .I3(GND_net), .O(Kp_23__N_1647));
    defparam i2_3_lut_adj_1190.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1191 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[14] [7]), 
            .I2(\data_in_frame[10] [5]), .I3(GND_net), .O(n26857));
    defparam i1_2_lut_3_lut_adj_1191.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1192 (.I0(n44398), .I1(n44412), .I2(n44161), 
            .I3(n27465), .O(n44736));
    defparam i1_4_lut_adj_1192.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1193 (.I0(n44674), .I1(\data_in_frame[8] [1]), 
            .I2(n41569), .I3(n44736), .O(n10_adj_4270));
    defparam i4_4_lut_adj_1193.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1194 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(n27394), .I3(\data_in_frame[8] [4]), .O(n4_adj_4250));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1194.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1195 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[8] [2]), 
            .I2(\data_out_frame[5] [6]), .I3(GND_net), .O(n10_adj_4126));   // verilog/coms.v(85[17:70])
    defparam i2_2_lut_3_lut_adj_1195.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i101 (.Q(\data_out_frame[12] [4]), .C(CLK_c), 
           .D(n28607));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1196 (.I0(\data_in_frame[10] [2]), .I1(n41451), 
            .I2(GND_net), .I3(GND_net), .O(n44227));
    defparam i1_2_lut_adj_1196.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1197 (.I0(\data_in_frame[12] [5]), .I1(\data_in_frame[14] [7]), 
            .I2(n25051), .I3(\data_in_frame[10] [3]), .O(n8_adj_4273));
    defparam i2_3_lut_4_lut_adj_1197.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1198 (.I0(n27058), .I1(\data_in_frame[10] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44353));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1198.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i102 (.Q(\data_out_frame[12] [5]), .C(CLK_c), 
           .D(n28606));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i103 (.Q(\data_out_frame[12] [6]), .C(CLK_c), 
           .D(n28605));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1199 (.I0(n26996), .I1(n4_adj_4250), .I2(\data_in_frame[12] [6]), 
            .I3(\data_in_frame[15] [0]), .O(n44439));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_4_lut_adj_1199.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1200 (.I0(n26996), .I1(n44353), .I2(\data_in_frame[17] [0]), 
            .I3(n44227), .O(n44769));   // verilog/coms.v(74[16:43])
    defparam i3_4_lut_adj_1200.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1201 (.I0(n26996), .I1(n4_adj_4250), .I2(n27058), 
            .I3(GND_net), .O(n48447));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1201.LUT_INIT = 16'h9696;
    SB_DFF data_out_frame_0___i104 (.Q(\data_out_frame[12] [7]), .C(CLK_c), 
           .D(n28604));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1202 (.I0(\data_in_frame[12] [4]), .I1(\data_in_frame[14] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44772));
    defparam i1_2_lut_adj_1202.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i105 (.Q(\data_out_frame[13] [0]), .C(CLK_c), 
           .D(n28603));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i106 (.Q(\data_out_frame[13] [1]), .C(CLK_c), 
           .D(n28602));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i107 (.Q(\data_out_frame[13] [2]), .C(CLK_c), 
           .D(n28601));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i108 (.Q(\data_out_frame[13] [3]), .C(CLK_c), 
           .D(n28600));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i109 (.Q(\data_out_frame[13] [4]), .C(CLK_c), 
           .D(n28599));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i110 (.Q(\data_out_frame[13] [5]), .C(CLK_c), 
           .D(n28598));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i111 (.Q(\data_out_frame[13] [6]), .C(CLK_c), 
           .D(n28597));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i112 (.Q(\data_out_frame[13] [7]), .C(CLK_c), 
           .D(n28596));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i113 (.Q(\data_out_frame[14] [0]), .C(CLK_c), 
           .D(n28595));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i114 (.Q(\data_out_frame[14] [1]), .C(CLK_c), 
           .D(n28594));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i115 (.Q(\data_out_frame[14] [2]), .C(CLK_c), 
           .D(n28593));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i116 (.Q(\data_out_frame[14] [3]), .C(CLK_c), 
           .D(n28592));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 data_in_frame_16__7__I_0_3896_2_lut (.I0(\data_in_frame[16] [7]), 
            .I1(\data_in_frame[16] [6]), .I2(GND_net), .I3(GND_net), .O(Kp_23__N_1402));   // verilog/coms.v(78[16:27])
    defparam data_in_frame_16__7__I_0_3896_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_out_frame_0___i117 (.Q(\data_out_frame[14] [4]), .C(CLK_c), 
           .D(n28591));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i29945_2_lut_3_lut_4_lut (.I0(\FRAME_MATCHER.state_c [2]), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(n33308), .I3(\FRAME_MATCHER.state[0] ), .O(n61));   // verilog/coms.v(127[12] 300[6])
    defparam i29945_2_lut_3_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i3_4_lut_adj_1203 (.I0(Kp_23__N_1402), .I1(n44772), .I2(n44769), 
            .I3(\data_in_frame[12] [5]), .O(n44464));
    defparam i3_4_lut_adj_1203.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i118 (.Q(\data_out_frame[14] [5]), .C(CLK_c), 
           .D(n28590));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i119 (.Q(\data_out_frame[14] [6]), .C(CLK_c), 
           .D(n28589));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i120 (.Q(\data_out_frame[14] [7]), .C(CLK_c), 
           .D(n28588));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i121 (.Q(\data_out_frame[15] [0]), .C(CLK_c), 
           .D(n28587));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i122 (.Q(\data_out_frame[15] [1]), .C(CLK_c), 
           .D(n28586));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i123 (.Q(\data_out_frame[15] [2]), .C(CLK_c), 
           .D(n28585));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i124 (.Q(\data_out_frame[15] [3]), .C(CLK_c), 
           .D(n28584));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i125 (.Q(\data_out_frame[15] [4]), .C(CLK_c), 
           .D(n28583));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i126 (.Q(\data_out_frame[15] [5]), .C(CLK_c), 
           .D(n28582));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i127 (.Q(\data_out_frame[15] [6]), .C(CLK_c), 
           .D(n28581));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i128 (.Q(\data_out_frame[15] [7]), .C(CLK_c), 
           .D(n28580));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i129 (.Q(\data_out_frame[16] [0]), .C(CLK_c), 
           .D(n28579));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i130 (.Q(\data_out_frame[16] [1]), .C(CLK_c), 
           .D(n28578));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i131 (.Q(\data_out_frame[16] [2]), .C(CLK_c), 
           .D(n28577));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i132 (.Q(\data_out_frame[16] [3]), .C(CLK_c), 
           .D(n28576));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i133 (.Q(\data_out_frame[16] [4]), .C(CLK_c), 
           .D(n28575));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i134 (.Q(\data_out_frame[16] [5]), .C(CLK_c), 
           .D(n28574));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i135 (.Q(\data_out_frame[16] [6]), .C(CLK_c), 
           .D(n28573));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i136 (.Q(\data_out_frame[16] [7]), .C(CLK_c), 
           .D(n28572));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i137 (.Q(\data_out_frame[17] [0]), .C(CLK_c), 
           .D(n28571));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i138 (.Q(\data_out_frame[17] [1]), .C(CLK_c), 
           .D(n28570));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i139 (.Q(\data_out_frame[17] [2]), .C(CLK_c), 
           .D(n28569));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i140 (.Q(\data_out_frame[17] [3]), .C(CLK_c), 
           .D(n28568));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i141 (.Q(\data_out_frame[17] [4]), .C(CLK_c), 
           .D(n28567));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i142 (.Q(\data_out_frame[17] [5]), .C(CLK_c), 
           .D(n28566));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i143 (.Q(\data_out_frame[17] [6]), .C(CLK_c), 
           .D(n28565));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i144 (.Q(\data_out_frame[17] [7]), .C(CLK_c), 
           .D(n28564));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i145 (.Q(\data_out_frame[18][0] ), .C(CLK_c), 
           .D(n28563));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i146 (.Q(\data_out_frame[18]_c [1]), .C(CLK_c), 
           .D(n28562));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i147 (.Q(\data_out_frame[18][2] ), .C(CLK_c), 
           .D(n28561));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i148 (.Q(\data_out_frame[18] [3]), .C(CLK_c), 
           .D(n28560));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i149 (.Q(\data_out_frame[18] [4]), .C(CLK_c), 
           .D(n28559));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i150 (.Q(\data_out_frame[18] [5]), .C(CLK_c), 
           .D(n28558));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i151 (.Q(\data_out_frame[18] [6]), .C(CLK_c), 
           .D(n28557));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i152 (.Q(\data_out_frame[18] [7]), .C(CLK_c), 
           .D(n28556));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i153 (.Q(\data_out_frame[19] [0]), .C(CLK_c), 
           .D(n28555));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i154 (.Q(\data_out_frame[19] [1]), .C(CLK_c), 
           .D(n28554));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i155 (.Q(\data_out_frame[19] [2]), .C(CLK_c), 
           .D(n28553));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i156 (.Q(\data_out_frame[19] [3]), .C(CLK_c), 
           .D(n28552));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i157 (.Q(\data_out_frame[19] [4]), .C(CLK_c), 
           .D(n28551));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i158 (.Q(\data_out_frame[19] [5]), .C(CLK_c), 
           .D(n28550));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i159 (.Q(\data_out_frame[19] [6]), .C(CLK_c), 
           .D(n28549));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i160 (.Q(\data_out_frame[19] [7]), .C(CLK_c), 
           .D(n28548));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i161 (.Q(\data_out_frame[20] [0]), .C(CLK_c), 
           .D(n28547));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i162 (.Q(\data_out_frame[20] [1]), .C(CLK_c), 
           .D(n28546));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i163 (.Q(\data_out_frame[20] [2]), .C(CLK_c), 
           .D(n28545));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i164 (.Q(\data_out_frame[20] [3]), .C(CLK_c), 
           .D(n28544));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i165 (.Q(\data_out_frame[20] [4]), .C(CLK_c), 
           .D(n28543));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i166 (.Q(\data_out_frame[20] [5]), .C(CLK_c), 
           .D(n28542));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i167 (.Q(\data_out_frame[20] [6]), .C(CLK_c), 
           .D(n28541));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i168 (.Q(\data_out_frame[20] [7]), .C(CLK_c), 
           .D(n28540));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i185 (.Q(\data_out_frame[23] [0]), .C(CLK_c), 
           .D(n28539));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i186 (.Q(\data_out_frame[23] [1]), .C(CLK_c), 
           .D(n28538));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i187 (.Q(\data_out_frame[23] [2]), .C(CLK_c), 
           .D(n28537));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i188 (.Q(\data_out_frame[23] [3]), .C(CLK_c), 
           .D(n28536));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i189 (.Q(\data_out_frame[23] [4]), .C(CLK_c), 
           .D(n28535));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i190 (.Q(\data_out_frame[23] [5]), .C(CLK_c), 
           .D(n28534));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i191 (.Q(\data_out_frame[23] [6]), .C(CLK_c), 
           .D(n28533));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i192 (.Q(\data_out_frame[23] [7]), .C(CLK_c), 
           .D(n28532));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i193 (.Q(\data_out_frame[24] [0]), .C(CLK_c), 
           .D(n28531));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i194 (.Q(\data_out_frame[24] [1]), .C(CLK_c), 
           .D(n28530));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i195 (.Q(\data_out_frame[24] [2]), .C(CLK_c), 
           .D(n28529));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i196 (.Q(\data_out_frame[24] [3]), .C(CLK_c), 
           .D(n28528));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1204 (.I0(\data_in_frame[9] [5]), .I1(n44148), 
            .I2(n44207), .I3(n41474), .O(n41956));   // verilog/coms.v(85[17:28])
    defparam i1_3_lut_4_lut_adj_1204.LUT_INIT = 16'h6996;
    SB_DFF data_out_frame_0___i197 (.Q(\data_out_frame[24] [4]), .C(CLK_c), 
           .D(n28527));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i198 (.Q(\data_out_frame[24] [5]), .C(CLK_c), 
           .D(n28526));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i199 (.Q(\data_out_frame[24] [6]), .C(CLK_c), 
           .D(n28525));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i200 (.Q(\data_out_frame[24] [7]), .C(CLK_c), 
           .D(n28524));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i201 (.Q(\data_out_frame[25] [0]), .C(CLK_c), 
           .D(n28523));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i202 (.Q(\data_out_frame[25] [1]), .C(CLK_c), 
           .D(n28522));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1205 (.I0(Kp_23__N_1114), .I1(\data_in_frame[8] [7]), 
            .I2(\data_in_frame[8] [6]), .I3(n44603), .O(n27606));
    defparam i1_2_lut_4_lut_adj_1205.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1206 (.I0(Kp_23__N_1114), .I1(\data_in_frame[8] [7]), 
            .I2(\data_in_frame[8] [6]), .I3(n26966), .O(n27650));
    defparam i1_2_lut_4_lut_adj_1206.LUT_INIT = 16'h6996;
    SB_DFF IntegralLimit_i0_i0 (.Q(IntegralLimit[0]), .C(CLK_c), .D(n28189));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i171 (.Q(\data_in_frame[21] [2]), .C(CLK_c), 
           .D(n28321));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i203 (.Q(\data_out_frame[25] [2]), .C(CLK_c), 
           .D(n28521));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i204 (.Q(\data_out_frame[25] [3]), .C(CLK_c), 
           .D(n28520));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i205 (.Q(\data_out_frame[25] [4]), .C(CLK_c), 
           .D(n28519));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i206 (.Q(\data_out_frame[25] [5]), .C(CLK_c), 
           .D(n28518));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i207 (.Q(\data_out_frame[25] [6]), .C(CLK_c), 
           .D(n28517));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_out_frame_0___i208 (.Q(\data_out_frame[25] [7]), .C(CLK_c), 
           .D(n28516));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i1 (.Q(neopxl_color[1]), .C(CLK_c), .D(n28515));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i2 (.Q(neopxl_color[2]), .C(CLK_c), .D(n28514));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1207 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [3]), 
            .I2(\data_in_frame[11] [3]), .I3(Kp_23__N_1233), .O(n44648));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_4_lut_adj_1207.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1208 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(\data_out_frame[8] [3]), .I3(n27288), .O(n44524));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_4_lut_adj_1208.LUT_INIT = 16'h6996;
    SB_DFF neopxl_color_i0_i3 (.Q(neopxl_color[3]), .C(CLK_c), .D(n28513));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i4 (.Q(neopxl_color[4]), .C(CLK_c), .D(n28512));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i5 (.Q(neopxl_color[5]), .C(CLK_c), .D(n28511));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i6 (.Q(neopxl_color[6]), .C(CLK_c), .D(n28510));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i7 (.Q(neopxl_color[7]), .C(CLK_c), .D(n28509));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i8 (.Q(neopxl_color[8]), .C(CLK_c), .D(n28508));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i9 (.Q(neopxl_color[9]), .C(CLK_c), .D(n28507));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i10 (.Q(neopxl_color[10]), .C(CLK_c), .D(n28506));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i11 (.Q(neopxl_color[11]), .C(CLK_c), .D(n28505));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i12 (.Q(neopxl_color[12]), .C(CLK_c), .D(n28504));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i13 (.Q(neopxl_color[13]), .C(CLK_c), .D(n28503));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i14 (.Q(neopxl_color[14]), .C(CLK_c), .D(n28502));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i15 (.Q(neopxl_color[15]), .C(CLK_c), .D(n28501));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i16 (.Q(neopxl_color[16]), .C(CLK_c), .D(n28500));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i17 (.Q(neopxl_color[17]), .C(CLK_c), .D(n28499));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i18 (.Q(neopxl_color[18]), .C(CLK_c), .D(n28498));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i19 (.Q(neopxl_color[19]), .C(CLK_c), .D(n28497));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i20 (.Q(neopxl_color[20]), .C(CLK_c), .D(n28496));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i21 (.Q(neopxl_color[21]), .C(CLK_c), .D(n28495));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i22 (.Q(neopxl_color[22]), .C(CLK_c), .D(n28494));   // verilog/coms.v(127[12] 300[6])
    SB_DFF neopxl_color_i0_i23 (.Q(neopxl_color[23]), .C(CLK_c), .D(n28493));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i2 (.Q(\data_in_frame[0] [1]), .C(CLK_c), .D(n28492));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i3 (.Q(\data_in_frame[0] [2]), .C(CLK_c), .D(n28491));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i4 (.Q(\data_in_frame[0] [3]), .C(CLK_c), .D(n28490));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i5 (.Q(\data_in_frame[0] [4]), .C(CLK_c), .D(n28489));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i6 (.Q(\data_in_frame[0] [5]), .C(CLK_c), .D(n28488));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i7 (.Q(\data_in_frame[0] [6]), .C(CLK_c), .D(n28485));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i8 (.Q(\data_in_frame[0] [7]), .C(CLK_c), .D(n28484));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i9 (.Q(\data_in_frame[1] [0]), .C(CLK_c), .D(n28483));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i10 (.Q(\data_in_frame[1] [1]), .C(CLK_c), .D(n28482));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i11 (.Q(\data_in_frame[1] [2]), .C(CLK_c), .D(n28481));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i12 (.Q(\data_in_frame[1] [3]), .C(CLK_c), .D(n28480));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i13 (.Q(\data_in_frame[1] [4]), .C(CLK_c), .D(n28479));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i14 (.Q(\data_in_frame[1] [5]), .C(CLK_c), .D(n28478));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i15 (.Q(\data_in_frame[1] [6]), .C(CLK_c), .D(n28477));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1209 (.I0(\data_in_frame[6] [3]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n26938));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1209.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i16 (.Q(\data_in_frame[1] [7]), .C(CLK_c), .D(n28476));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i17 (.Q(\data_in_frame[2] [0]), .C(CLK_c), .D(n28475));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i18 (.Q(\data_in_frame[2] [1]), .C(CLK_c), .D(n28474));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i19 (.Q(\data_in_frame[2] [2]), .C(CLK_c), .D(n28473));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i20 (.Q(\data_in_frame[2] [3]), .C(CLK_c), .D(n28472));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i21 (.Q(\data_in_frame[2] [4]), .C(CLK_c), .D(n28471));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i22 (.Q(\data_in_frame[2] [5]), .C(CLK_c), .D(n28470));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i23 (.Q(\data_in_frame[2] [6]), .C(CLK_c), .D(n28469));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i24 (.Q(\data_in_frame[2] [7]), .C(CLK_c), .D(n28468));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i25 (.Q(\data_in_frame[3] [0]), .C(CLK_c), .D(n28467));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1210 (.I0(n26866), .I1(n44190), .I2(GND_net), 
            .I3(GND_net), .O(n44760));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1210.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i26 (.Q(\data_in_frame[3] [1]), .C(CLK_c), .D(n28466));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i27 (.Q(\data_in_frame[3] [2]), .C(CLK_c), .D(n28465));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_4_lut_adj_1211 (.I0(\data_in_frame[8] [2]), .I1(n44398), 
            .I2(n44642), .I3(\data_in_frame[6] [1]), .O(n44339));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_4_lut_adj_1211.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1212 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[7] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44591));   // verilog/coms.v(70[16:27])
    defparam i1_2_lut_adj_1212.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i28 (.Q(\data_in_frame[3] [3]), .C(CLK_c), .D(n28464));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i29 (.Q(\data_in_frame[3] [4]), .C(CLK_c), .D(n28463));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i30 (.Q(\data_in_frame[3] [5]), .C(CLK_c), .D(n28462));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i31 (.Q(\data_in_frame[3] [6]), .C(CLK_c), .D(n28461));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i32 (.Q(\data_in_frame[3] [7]), .C(CLK_c), .D(n28460));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i33 (.Q(\data_in_frame[4] [0]), .C(CLK_c), .D(n28459));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i34 (.Q(\data_in_frame[4] [1]), .C(CLK_c), .D(n28458));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i35 (.Q(\data_in_frame[4] [2]), .C(CLK_c), .D(n28457));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i36 (.Q(\data_in_frame[4] [3]), .C(CLK_c), .D(n28456));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1213 (.I0(\data_in_frame[3] [6]), .I1(\data_in_frame[6] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n27465));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1213.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i37 (.Q(\data_in_frame[4] [4]), .C(CLK_c), .D(n28455));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i38 (.Q(\data_in_frame[4] [5]), .C(CLK_c), .D(n28454));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i39 (.Q(\data_in_frame[4] [6]), .C(CLK_c), .D(n28453));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1214 (.I0(Kp_23__N_836), .I1(n44339), .I2(n27465), 
            .I3(n27063), .O(n27058));   // verilog/coms.v(76[16:43])
    defparam i3_4_lut_adj_1214.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i40 (.Q(\data_in_frame[4] [7]), .C(CLK_c), .D(n28452));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_4_lut_adj_1215 (.I0(n27584), .I1(n44594), .I2(n44591), 
            .I3(\data_in_frame[6] [7]), .O(n27411));   // verilog/coms.v(70[16:27])
    defparam i3_4_lut_adj_1215.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i41 (.Q(\data_in_frame[5] [0]), .C(CLK_c), .D(n28451));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i42 (.Q(\data_in_frame[5] [1]), .C(CLK_c), .D(n28450));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i43 (.Q(\data_in_frame[5] [2]), .C(CLK_c), .D(n28449));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i44 (.Q(\data_in_frame[5] [3]), .C(CLK_c), .D(n28448));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1216 (.I0(\data_in_frame[9] [1]), .I1(\data_in_frame[9] [3]), 
            .I2(\data_in_frame[9] [2]), .I3(\data_in_frame[9] [4]), .O(n27597));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_3_lut_4_lut_adj_1216.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i45 (.Q(\data_in_frame[5] [4]), .C(CLK_c), .D(n28447));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i46 (.Q(\data_in_frame[5] [5]), .C(CLK_c), .D(n28446));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i47 (.Q(\data_in_frame[5] [6]), .C(CLK_c), .D(n28445));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i48 (.Q(\data_in_frame[5] [7]), .C(CLK_c), .D(n28444));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1217 (.I0(\data_in_frame[6] [1]), .I1(\data_in_frame[6] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44706));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1217.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i49 (.Q(\data_in_frame[6] [0]), .C(CLK_c), .D(n28443));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i50 (.Q(\data_in_frame[6] [1]), .C(CLK_c), .D(n28442));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1218 (.I0(\data_in_frame[9] [5]), .I1(\data_in_frame[9] [7]), 
            .I2(\data_in_frame[9] [6]), .I3(n44677), .O(n48461));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_4_lut_adj_1218.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i51 (.Q(\data_in_frame[6] [2]), .C(CLK_c), .D(n28441));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1219 (.I0(n26770), .I1(\data_in_frame[6] [6]), 
            .I2(\data_in_frame[7] [0]), .I3(n44294), .O(n10_adj_4271));   // verilog/coms.v(236[9:81])
    defparam i4_4_lut_adj_1219.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i52 (.Q(\data_in_frame[6] [3]), .C(CLK_c), .D(n28440));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i53 (.Q(\data_in_frame[6] [4]), .C(CLK_c), .D(n28439));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i54 (.Q(\data_in_frame[6] [5]), .C(CLK_c), .D(n28438));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i55 (.Q(\data_in_frame[6] [6]), .C(CLK_c), .D(n28437));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i56 (.Q(\data_in_frame[6] [7]), .C(CLK_c), .D(n28436));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_4_lut_adj_1220 (.I0(\data_in_frame[5] [7]), .I1(n44556), 
            .I2(\data_in_frame[8] [3]), .I3(\data_in_frame[4] [1]), .O(n12_adj_4275));   // verilog/coms.v(78[16:27])
    defparam i5_4_lut_adj_1220.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1221 (.I0(\data_in_frame[2] [0]), .I1(n12_adj_4275), 
            .I2(n44706), .I3(\data_in_frame[1] [7]), .O(n26996));   // verilog/coms.v(78[16:27])
    defparam i6_4_lut_adj_1221.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1222 (.I0(\data_in_frame[5] [2]), .I1(n27579), 
            .I2(\data_in_frame[5] [3]), .I3(n44454), .O(n10_adj_4264));
    defparam i4_4_lut_adj_1222.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i57 (.Q(\data_in_frame[7] [0]), .C(CLK_c), .D(n28435));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1223 (.I0(\FRAME_MATCHER.state_c [2]), 
            .I1(\FRAME_MATCHER.state_c [1]), .I2(\FRAME_MATCHER.state[0] ), 
            .I3(n33308), .O(\FRAME_MATCHER.i_31__N_2524 ));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_4_lut_adj_1223.LUT_INIT = 16'h0020;
    SB_LUT4 i1_2_lut_adj_1224 (.I0(\data_in_frame[6] [6]), .I1(\data_in_frame[6] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26978));   // verilog/coms.v(77[16:43])
    defparam i1_2_lut_adj_1224.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i58 (.Q(\data_in_frame[7] [1]), .C(CLK_c), .D(n28434));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i59 (.Q(\data_in_frame[7] [2]), .C(CLK_c), .D(n28433));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1225 (.I0(n27334), .I1(n44360), .I2(n26978), 
            .I3(GND_net), .O(Kp_23__N_1114));
    defparam i2_3_lut_adj_1225.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i60 (.Q(\data_in_frame[7] [3]), .C(CLK_c), .D(n28432));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1226 (.I0(\data_in_frame[7] [5]), .I1(\data_in_frame[3] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4276));
    defparam i1_2_lut_adj_1226.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i61 (.Q(\data_in_frame[7] [4]), .C(CLK_c), .D(n28431));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1227 (.I0(\data_in_frame[5] [3]), .I1(\data_in_frame[5] [4]), 
            .I2(n27198), .I3(n6_adj_4276), .O(n44307));
    defparam i4_4_lut_adj_1227.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i62 (.Q(\data_in_frame[7] [5]), .C(CLK_c), .D(n28430));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i63 (.Q(\data_in_frame[7] [6]), .C(CLK_c), .D(n28429));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i64 (.Q(\data_in_frame[7] [7]), .C(CLK_c), .D(n28428));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i65 (.Q(\data_in_frame[8] [0]), .C(CLK_c), .D(n28427));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i66 (.Q(\data_in_frame[8] [1]), .C(CLK_c), .D(n28426));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i67 (.Q(\data_in_frame[8] [2]), .C(CLK_c), .D(n28425));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i68 (.Q(\data_in_frame[8] [3]), .C(CLK_c), .D(n28424));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1228 (.I0(\data_in_frame[14] [5]), .I1(n44665), 
            .I2(n27459), .I3(GND_net), .O(n44378));
    defparam i1_3_lut_4_lut_adj_1228.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i69 (.Q(\data_in_frame[8] [4]), .C(CLK_c), .D(n28423));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 n51453_bdd_4_lut (.I0(n51453), .I1(\data_out_frame[17] [7]), 
            .I2(\data_out_frame[16] [7]), .I3(byte_transmit_counter[1]), 
            .O(n51456));
    defparam n51453_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_DFF data_in_frame_0__i70 (.Q(\data_in_frame[8] [5]), .C(CLK_c), .D(n28422));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1229 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(\FRAME_MATCHER.state_c [2]), .I3(GND_net), .O(n44035));
    defparam i1_2_lut_3_lut_adj_1229.LUT_INIT = 16'h8080;
    SB_DFF data_in_frame_0__i71 (.Q(\data_in_frame[8] [6]), .C(CLK_c), .D(n28421));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i5_4_lut_adj_1230 (.I0(n27579), .I1(n44594), .I2(\data_in_frame[7] [2]), 
            .I3(n26834), .O(n12_adj_4277));
    defparam i5_4_lut_adj_1230.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1231 (.I0(\data_in_frame[5] [1]), .I1(n12_adj_4277), 
            .I2(n44709), .I3(n25836), .O(n27414));
    defparam i6_4_lut_adj_1231.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i72 (.Q(\data_in_frame[8] [7]), .C(CLK_c), .D(n28420));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i73 (.Q(\data_in_frame[9] [0]), .C(CLK_c), .D(n28419));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i74 (.Q(\data_in_frame[9] [1]), .C(CLK_c), .D(n28418));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 equal_1544_i8_2_lut (.I0(Kp_23__N_1114), .I1(\data_in_frame[8] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n8_adj_4278));   // verilog/coms.v(236[9:81])
    defparam equal_1544_i8_2_lut.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i75 (.Q(\data_in_frame[9] [2]), .C(CLK_c), .D(n28417));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i76 (.Q(\data_in_frame[9] [3]), .C(CLK_c), .D(n28416));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i77 (.Q(\data_in_frame[9] [4]), .C(CLK_c), .D(n28415));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1232 (.I0(\data_in_frame[15] [1]), .I1(\data_in_frame[12] [7]), 
            .I2(\data_in_frame[13] [1]), .I3(\data_in_frame[17] [3]), .O(n7_adj_4272));
    defparam i1_2_lut_4_lut_adj_1232.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1233 (.I0(\data_in_frame[1] [6]), .I1(\data_in_frame[4] [0]), 
            .I2(\data_in_frame[3] [7]), .I3(GND_net), .O(n44301));
    defparam i2_3_lut_adj_1233.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i78 (.Q(\data_in_frame[9] [5]), .C(CLK_c), .D(n28414));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i79 (.Q(\data_in_frame[9] [6]), .C(CLK_c), .D(n28413));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i3_3_lut_4_lut (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(\FRAME_MATCHER.state_c [2]), .I3(n33308), .O(\FRAME_MATCHER.i_31__N_2526 ));
    defparam i3_3_lut_4_lut.LUT_INIT = 16'h0008;
    SB_DFF data_in_frame_0__i80 (.Q(\data_in_frame[9] [7]), .C(CLK_c), .D(n28412));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i81 (.Q(\data_in_frame[10] [0]), .C(CLK_c), 
           .D(n28411));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i82 (.Q(\data_in_frame[10] [1]), .C(CLK_c), 
           .D(n28410));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i83 (.Q(\data_in_frame[10] [2]), .C(CLK_c), 
           .D(n28409));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i84 (.Q(\data_in_frame[10] [3]), .C(CLK_c), 
           .D(n28408));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i85 (.Q(\data_in_frame[10] [4]), .C(CLK_c), 
           .D(n28407));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i86 (.Q(\data_in_frame[10] [5]), .C(CLK_c), 
           .D(n28406));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i87 (.Q(\data_in_frame[10] [6]), .C(CLK_c), 
           .D(n28405));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i88 (.Q(\data_in_frame[10] [7]), .C(CLK_c), 
           .D(n28404));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i89 (.Q(\data_in_frame[11] [0]), .C(CLK_c), 
           .D(n28403));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1234 (.I0(\data_out_frame[12] [7]), .I1(\data_out_frame[12] [6]), 
            .I2(\data_out_frame[12] [0]), .I3(GND_net), .O(n44543));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_adj_1234.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i90 (.Q(\data_in_frame[11] [1]), .C(CLK_c), 
           .D(n28402));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i91 (.Q(\data_in_frame[11] [2]), .C(CLK_c), 
           .D(n28401));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i92 (.Q(\data_in_frame[11] [3]), .C(CLK_c), 
           .D(n28400));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i93 (.Q(\data_in_frame[11] [4]), .C(CLK_c), 
           .D(n28399));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i94 (.Q(\data_in_frame[11] [5]), .C(CLK_c), 
           .D(n28398));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i95 (.Q(\data_in_frame[11] [6]), .C(CLK_c), 
           .D(n28397));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i96 (.Q(\data_in_frame[11] [7]), .C(CLK_c), 
           .D(n28396));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i97 (.Q(\data_in_frame[12] [0]), .C(CLK_c), 
           .D(n28395));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i98 (.Q(\data_in_frame[12] [1]), .C(CLK_c), 
           .D(n28394));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i99 (.Q(\data_in_frame[12] [2]), .C(CLK_c), 
           .D(n28393));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i100 (.Q(\data_in_frame[12] [3]), .C(CLK_c), 
           .D(n28392));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i101 (.Q(\data_in_frame[12] [4]), .C(CLK_c), 
           .D(n28391));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i102 (.Q(\data_in_frame[12] [5]), .C(CLK_c), 
           .D(n28390));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i103 (.Q(\data_in_frame[12] [6]), .C(CLK_c), 
           .D(n28389));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i104 (.Q(\data_in_frame[12] [7]), .C(CLK_c), 
           .D(n28388));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i105 (.Q(\data_in_frame[13] [0]), .C(CLK_c), 
           .D(n28387));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i106 (.Q(\data_in_frame[13] [1]), .C(CLK_c), 
           .D(n28386));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i107 (.Q(\data_in_frame[13] [2]), .C(CLK_c), 
           .D(n28385));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i108 (.Q(\data_in_frame[13] [3]), .C(CLK_c), 
           .D(n28384));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i109 (.Q(\data_in_frame[13] [4]), .C(CLK_c), 
           .D(n28383));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i110 (.Q(\data_in_frame[13] [5]), .C(CLK_c), 
           .D(n28382));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1235 (.I0(Kp_23__N_996), .I1(n41468), .I2(GND_net), 
            .I3(GND_net), .O(n44639));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1235.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i111 (.Q(\data_in_frame[13] [6]), .C(CLK_c), 
           .D(n28381));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1236 (.I0(n44301), .I1(n44398), .I2(n44234), 
            .I3(GND_net), .O(Kp_23__N_836));   // verilog/coms.v(78[16:27])
    defparam i2_3_lut_adj_1236.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i112 (.Q(\data_in_frame[13] [7]), .C(CLK_c), 
           .D(n28380));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i4_4_lut_adj_1237 (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[2] [0]), 
            .I2(\data_in_frame[4] [3]), .I3(n6_adj_4265), .O(Kp_23__N_996));   // verilog/coms.v(73[16:42])
    defparam i4_4_lut_adj_1237.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i113 (.Q(\data_in_frame[14] [0]), .C(CLK_c), 
           .D(n28379));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1238 (.I0(\data_in_frame[7] [7]), .I1(\data_in_frame[8] [1]), 
            .I2(n27530), .I3(GND_net), .O(n44627));
    defparam i1_2_lut_3_lut_adj_1238.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i114 (.Q(\data_in_frame[14] [1]), .C(CLK_c), 
           .D(n28378));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1239 (.I0(Kp_23__N_996), .I1(\data_in_frame[6] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44345));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1239.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i115 (.Q(\data_in_frame[14] [2]), .C(CLK_c), 
           .D(n28377));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i116 (.Q(\data_in_frame[14] [3]), .C(CLK_c), 
           .D(n28376));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1240 (.I0(n27530), .I1(n44170), .I2(GND_net), 
            .I3(GND_net), .O(n41569));
    defparam i1_2_lut_adj_1240.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i117 (.Q(\data_in_frame[14] [4]), .C(CLK_c), 
           .D(n28375));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i118 (.Q(\data_in_frame[14] [5]), .C(CLK_c), 
           .D(n28374));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i119 (.Q(\data_in_frame[14] [6]), .C(CLK_c), 
           .D(n28373));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i120 (.Q(\data_in_frame[14] [7]), .C(CLK_c), 
           .D(n28372));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i121 (.Q(\data_in_frame[15] [0]), .C(CLK_c), 
           .D(n28371));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i122 (.Q(\data_in_frame[15] [1]), .C(CLK_c), 
           .D(n28370));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i123 (.Q(\data_in_frame[15] [2]), .C(CLK_c), 
           .D(n28369));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i124 (.Q(\data_in_frame[15] [3]), .C(CLK_c), 
           .D(n28368));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i125 (.Q(\data_in_frame[15] [4]), .C(CLK_c), 
           .D(n28367));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i126 (.Q(\data_in_frame[15] [5]), .C(CLK_c), 
           .D(n28366));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i127 (.Q(\data_in_frame[15] [6]), .C(CLK_c), 
           .D(n28365));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i128 (.Q(\data_in_frame[15] [7]), .C(CLK_c), 
           .D(n28364));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i129 (.Q(\data_in_frame[16] [0]), .C(CLK_c), 
           .D(n28363));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1241 (.I0(Kp_23__N_999), .I1(n44345), .I2(\data_in_frame[6] [5]), 
            .I3(GND_net), .O(Kp_23__N_1095));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1241.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i130 (.Q(\data_in_frame[16] [1]), .C(CLK_c), 
           .D(n28362));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1242 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44261));   // verilog/coms.v(166[9:87])
    defparam i1_2_lut_adj_1242.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1243 (.I0(n44464), .I1(\data_in_frame[14] [5]), 
            .I2(n27297), .I3(n44665), .O(Kp_23__N_1644));
    defparam i1_2_lut_4_lut_adj_1243.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i131 (.Q(\data_in_frame[16] [2]), .C(CLK_c), 
           .D(n28361));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_2_lut_4_lut_adj_1244 (.I0(n44307), .I1(n10_adj_4263), .I2(\data_in_frame[5] [5]), 
            .I3(\data_in_frame[10] [1]), .O(n10_adj_4262));
    defparam i2_2_lut_4_lut_adj_1244.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i132 (.Q(\data_in_frame[16] [3]), .C(CLK_c), 
           .D(n28360));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1245 (.I0(\data_in_frame[1] [4]), .I1(\data_in_frame[5] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44642));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1245.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i133 (.Q(\data_in_frame[16] [4]), .C(CLK_c), 
           .D(n28359));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1246 (.I0(\data_in_frame[1] [5]), .I1(\data_in_frame[5] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n44398));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_adj_1246.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i134 (.Q(\data_in_frame[16] [5]), .C(CLK_c), 
           .D(n28358));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i135 (.Q(\data_in_frame[16] [6]), .C(CLK_c), 
           .D(n28357));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1247 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[3] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n44161));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1247.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i136 (.Q(\data_in_frame[16] [7]), .C(CLK_c), 
           .D(n28356));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i137 (.Q(\data_in_frame[17] [0]), .C(CLK_c), 
           .D(n28355));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i138 (.Q(\data_in_frame[17] [1]), .C(CLK_c), 
           .D(n28354));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i139 (.Q(\data_in_frame[17] [2]), .C(CLK_c), 
           .D(n28353));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i140 (.Q(\data_in_frame[17] [3]), .C(CLK_c), 
           .D(n28352));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i141 (.Q(\data_in_frame[17] [4]), .C(CLK_c), 
           .D(n28351));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i142 (.Q(\data_in_frame[17] [5]), .C(CLK_c), 
           .D(n28350));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i143 (.Q(\data_in_frame[17] [6]), .C(CLK_c), 
           .D(n28349));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i144 (.Q(\data_in_frame[17] [7]), .C(CLK_c), 
           .D(n28348));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i145 (.Q(\data_in_frame[18] [0]), .C(CLK_c), 
           .D(n28347));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i146 (.Q(\data_in_frame[18] [1]), .C(CLK_c), 
           .D(n28346));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i147 (.Q(\data_in_frame[18] [2]), .C(CLK_c), 
           .D(n28345));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i148 (.Q(\data_in_frame[18] [3]), .C(CLK_c), 
           .D(n28344));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_adj_1248 (.I0(\data_in_frame[1] [2]), .I1(\data_in_frame[0] [7]), 
            .I2(\data_in_frame[3] [3]), .I3(GND_net), .O(n44310));   // verilog/coms.v(73[16:34])
    defparam i1_3_lut_adj_1248.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i149 (.Q(\data_in_frame[18] [4]), .C(CLK_c), 
           .D(n28343));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_3_lut_4_lut_adj_1249 (.I0(n41445), .I1(n27023), .I2(n44458), 
            .I3(Kp_23__N_1233), .O(n42348));
    defparam i1_3_lut_4_lut_adj_1249.LUT_INIT = 16'h6996;
    SB_DFF data_in_frame_0__i150 (.Q(\data_in_frame[18] [5]), .C(CLK_c), 
           .D(n28342));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i151 (.Q(\data_in_frame[18] [6]), .C(CLK_c), 
           .D(n28341));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_4_lut_adj_1250 (.I0(\data_in_frame[13] [5]), .I1(n26966), 
            .I2(Kp_23__N_1114), .I3(\data_in_frame[8] [7]), .O(n44549));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1250.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1251 (.I0(\data_in_frame[5] [4]), .I1(n44454), 
            .I2(GND_net), .I3(GND_net), .O(n44674));
    defparam i1_2_lut_adj_1251.LUT_INIT = 16'h6666;
    SB_DFF data_in_frame_0__i152 (.Q(\data_in_frame[18] [7]), .C(CLK_c), 
           .D(n28340));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_3_lut_adj_1252 (.I0(\data_in_frame[9] [4]), .I1(n41445), 
            .I2(n27414), .I3(GND_net), .O(n41580));
    defparam i1_2_lut_3_lut_adj_1252.LUT_INIT = 16'h9696;
    SB_DFF data_in_frame_0__i153 (.Q(\data_in_frame[19] [0]), .C(CLK_c), 
           .D(n28339));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i154 (.Q(\data_in_frame[19] [1]), .C(CLK_c), 
           .D(n28338));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i155 (.Q(\data_in_frame[19] [2]), .C(CLK_c), 
           .D(n28337));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i156 (.Q(\data_in_frame[19] [3]), .C(CLK_c), 
           .D(n28336));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i157 (.Q(\data_in_frame[19] [4]), .C(CLK_c), 
           .D(n28335));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i7_4_lut_adj_1253 (.I0(\FRAME_MATCHER.state_c [11]), .I1(n14_adj_4268), 
            .I2(n10_adj_4267), .I3(\FRAME_MATCHER.state_c [13]), .O(n34549));
    defparam i7_4_lut_adj_1253.LUT_INIT = 16'hfffe;
    SB_DFF data_in_frame_0__i158 (.Q(\data_in_frame[19] [5]), .C(CLK_c), 
           .D(n28334));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i159 (.Q(\data_in_frame[19] [6]), .C(CLK_c), 
           .D(n28333));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i160 (.Q(\data_in_frame[19] [7]), .C(CLK_c), 
           .D(n28332));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i161 (.Q(\data_in_frame[20] [0]), .C(CLK_c), 
           .D(n28331));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i162 (.Q(\data_in_frame[20] [1]), .C(CLK_c), 
           .D(n28330));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i163 (.Q(\data_in_frame[20] [2]), .C(CLK_c), 
           .D(n28329));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i164 (.Q(\data_in_frame[20] [3]), .C(CLK_c), 
           .D(n28328));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i165 (.Q(\data_in_frame[20] [4]), .C(CLK_c), 
           .D(n28327));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i166 (.Q(\data_in_frame[20] [5]), .C(CLK_c), 
           .D(n28326));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i167 (.Q(\data_in_frame[20] [6]), .C(CLK_c), 
           .D(n28325));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i168 (.Q(\data_in_frame[20] [7]), .C(CLK_c), 
           .D(n28324));   // verilog/coms.v(127[12] 300[6])
    SB_DFF data_in_frame_0__i169 (.Q(\data_in_frame[21] [0]), .C(CLK_c), 
           .D(n28323));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i1_2_lut_adj_1254 (.I0(\data_in_frame[2] [7]), .I1(\data_in_frame[4] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44709));   // verilog/coms.v(73[16:42])
    defparam i1_2_lut_adj_1254.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1255 (.I0(\data_in_frame[4] [2]), .I1(\data_in_frame[3] [0]), 
            .I2(\data_in_frame[5] [3]), .I3(\data_in_frame[0] [4]), .O(n48339));   // verilog/coms.v(78[16:27])
    defparam i1_4_lut_adj_1255.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1256 (.I0(\data_in_frame[2] [0]), .I1(\data_in_frame[3] [4]), 
            .I2(\data_in_frame[1] [5]), .I3(\data_in_frame[2] [2]), .O(n48341));   // verilog/coms.v(78[16:27])
    defparam i1_4_lut_adj_1256.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1257 (.I0(n26966), .I1(n27411), .I2(\data_in_frame[9] [2]), 
            .I3(GND_net), .O(n27347));   // verilog/coms.v(72[16:41])
    defparam i1_2_lut_3_lut_adj_1257.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_adj_1258 (.I0(n48341), .I1(n44709), .I2(n48339), 
            .I3(GND_net), .O(n48347));   // verilog/coms.v(78[16:27])
    defparam i1_3_lut_adj_1258.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1259 (.I0(\data_in_frame[18] [1]), .I1(n46232), 
            .I2(\data_in_frame[20] [3]), .I3(n44656), .O(n45653));
    defparam i2_3_lut_4_lut_adj_1259.LUT_INIT = 16'h9669;
    SB_LUT4 i2_2_lut_3_lut_adj_1260 (.I0(n26966), .I1(Kp_23__N_1114), .I2(\data_in_frame[8] [7]), 
            .I3(GND_net), .O(Kp_23__N_1221));   // verilog/coms.v(85[17:70])
    defparam i2_2_lut_3_lut_adj_1260.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1261 (.I0(n44310), .I1(n48351), .I2(n48347), 
            .I3(n44363), .O(n48355));   // verilog/coms.v(78[16:27])
    defparam i1_4_lut_adj_1261.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1262 (.I0(\data_in_frame[18] [1]), .I1(n46232), 
            .I2(\data_in_frame[20] [2]), .I3(n44659), .O(n45673));
    defparam i2_3_lut_4_lut_adj_1262.LUT_INIT = 16'h9669;
    SB_LUT4 i1_3_lut_4_lut_adj_1263 (.I0(\data_in_frame[13] [4]), .I1(n44357), 
            .I2(n44406), .I3(\data_in_frame[15] [5]), .O(n41435));   // verilog/coms.v(76[16:43])
    defparam i1_3_lut_4_lut_adj_1263.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_4_lut_adj_1264 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(n44662), .I3(n41478), .O(n44395));   // verilog/coms.v(71[16:27])
    defparam i2_3_lut_4_lut_adj_1264.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1265 (.I0(\data_in_frame[13] [4]), .I1(n44357), 
            .I2(\data_in_frame[15] [6]), .I3(\data_in_frame[18] [0]), .O(n44230));   // verilog/coms.v(76[16:43])
    defparam i2_3_lut_4_lut_adj_1265.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1266 (.I0(n48355), .I1(n27660), .I2(n44556), 
            .I3(n26866), .O(n48361));   // verilog/coms.v(78[16:27])
    defparam i1_4_lut_adj_1266.LUT_INIT = 16'h6996;
    SB_LUT4 i1361_2_lut_3_lut (.I0(n31_adj_4279), .I1(n24120), .I2(\FRAME_MATCHER.state_c [1]), 
            .I3(GND_net), .O(n5785));
    defparam i1361_2_lut_3_lut.LUT_INIT = 16'h1010;
    SB_LUT4 i2_3_lut_4_lut_adj_1267 (.I0(n31_adj_4279), .I1(n24120), .I2(n33307), 
            .I3(\FRAME_MATCHER.state_c [2]), .O(n46360));
    defparam i2_3_lut_4_lut_adj_1267.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_3_lut_adj_1268 (.I0(\data_in_frame[14] [2]), .I1(\data_in_frame[16] [4]), 
            .I2(n41494), .I3(GND_net), .O(n44680));
    defparam i1_2_lut_3_lut_adj_1268.LUT_INIT = 16'h6969;
    SB_LUT4 i15301_3_lut_4_lut (.I0(n34417), .I1(n44095), .I2(rx_data[7]), 
            .I3(\data_in_frame[15] [7]), .O(n28364));
    defparam i15301_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1269 (.I0(\data_in_frame[6] [0]), .I1(\data_in_frame[6] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n48453));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_adj_1269.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1270 (.I0(n27584), .I1(n41468), .I2(n44336), 
            .I3(n48453), .O(n44170));   // verilog/coms.v(85[17:28])
    defparam i1_4_lut_adj_1270.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1271 (.I0(n26996), .I1(n27425), .I2(\data_in_frame[12] [7]), 
            .I3(n44754), .O(n44527));
    defparam i1_2_lut_4_lut_adj_1271.LUT_INIT = 16'h6996;
    SB_LUT4 i15302_3_lut_4_lut (.I0(n34417), .I1(n44095), .I2(rx_data[6]), 
            .I3(\data_in_frame[15] [6]), .O(n28365));
    defparam i15302_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_DFF data_in_frame_0__i170 (.Q(\data_in_frame[21] [1]), .C(CLK_c), 
           .D(n28322));   // verilog/coms.v(127[12] 300[6])
    SB_LUT4 i2_3_lut_adj_1272 (.I0(\data_in_frame[1] [0]), .I1(Kp_23__N_888), 
            .I2(\data_in_frame[0] [5]), .I3(GND_net), .O(n25836));   // verilog/coms.v(77[16:27])
    defparam i2_3_lut_adj_1272.LUT_INIT = 16'h9696;
    SB_LUT4 add_3971_9_lut (.I0(GND_net), .I1(byte_transmit_counter[7]), 
            .I2(GND_net), .I3(n39112), .O(n8825[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1_2_lut_adj_1273 (.I0(\data_in_frame[1] [3]), .I1(\data_in_frame[1] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44184));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_adj_1273.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1274 (.I0(\data_in_frame[19] [6]), .I1(n42281), 
            .I2(n46677), .I3(GND_net), .O(n44291));   // verilog/coms.v(268[9:85])
    defparam i1_2_lut_3_lut_adj_1274.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1275 (.I0(n26866), .I1(n44184), .I2(\data_in_frame[1] [1]), 
            .I3(\data_in_frame[1] [4]), .O(Kp_23__N_888));   // verilog/coms.v(73[16:34])
    defparam i3_4_lut_adj_1275.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1276 (.I0(\data_out_frame[16] [4]), .I1(\data_out_frame[18] [5]), 
            .I2(\data_out_frame[16] [2]), .I3(\data_out_frame[18] [4]), 
            .O(n26809));   // verilog/coms.v(85[17:28])
    defparam i1_2_lut_3_lut_4_lut_adj_1276.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1277 (.I0(\data_in_frame[4] [7]), .I1(\data_in_frame[3] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n48617));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1277.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1278 (.I0(\data_in_frame[5] [2]), .I1(n48617), 
            .I2(\data_in_frame[2] [6]), .I3(\data_in_frame[5] [1]), .O(n44243));   // verilog/coms.v(85[17:70])
    defparam i1_4_lut_adj_1278.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1279 (.I0(\data_in_frame[15] [7]), .I1(n44648), 
            .I2(\data_in_frame[17] [7]), .I3(GND_net), .O(n48653));
    defparam i1_2_lut_3_lut_adj_1279.LUT_INIT = 16'h9696;
    SB_LUT4 add_3971_8_lut (.I0(GND_net), .I1(byte_transmit_counter[6]), 
            .I2(GND_net), .I3(n39111), .O(n8825[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 data_in_frame_0__5__I_0_2_lut (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(GND_net), .I3(GND_net), .O(Kp_23__N_881));   // verilog/coms.v(76[16:27])
    defparam data_in_frame_0__5__I_0_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1280 (.I0(n27198), .I1(n44243), .I2(GND_net), 
            .I3(GND_net), .O(n6_adj_4280));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_adj_1280.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1281 (.I0(\data_in_frame[7] [3]), .I1(n26770), 
            .I2(Kp_23__N_881), .I3(n6_adj_4280), .O(n41445));   // verilog/coms.v(85[17:70])
    defparam i4_4_lut_adj_1281.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1282 (.I0(\data_in_frame[8] [0]), .I1(n48477), 
            .I2(n44170), .I3(n27063), .O(n44412));
    defparam i1_4_lut_adj_1282.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1283 (.I0(\data_in_frame[0] [2]), .I1(\data_in_frame[0] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n44142));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_adj_1283.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1284 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[4] [4]), 
            .I2(\data_in_frame[2] [1]), .I3(\data_in_frame[4] [3]), .O(n44363));   // verilog/coms.v(74[16:43])
    defparam i1_4_lut_adj_1284.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1285 (.I0(n27337), .I1(n44363), .I2(\data_in_frame[1] [7]), 
            .I3(GND_net), .O(Kp_23__N_999));   // verilog/coms.v(74[16:43])
    defparam i2_3_lut_adj_1285.LUT_INIT = 16'h9696;
    SB_CARRY add_3971_8 (.CI(n39111), .I0(byte_transmit_counter[6]), .I1(GND_net), 
            .CO(n39112));
    SB_LUT4 i1_2_lut_adj_1286 (.I0(\data_in_frame[4] [1]), .I1(\data_in_frame[4] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n27360));
    defparam i1_2_lut_adj_1286.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1287 (.I0(\data_in_frame[11] [5]), .I1(\data_in_frame[9] [2]), 
            .I2(\data_in_frame[9] [4]), .I3(GND_net), .O(n27312));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1287.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1288 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [0]), 
            .I2(\data_in_frame[2] [2]), .I3(GND_net), .O(n27356));   // verilog/coms.v(73[16:42])
    defparam i2_3_lut_adj_1288.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1289 (.I0(\data_in_frame[11] [3]), .I1(n27347), 
            .I2(n27606), .I3(GND_net), .O(n44357));   // verilog/coms.v(76[16:43])
    defparam i1_2_lut_3_lut_adj_1289.LUT_INIT = 16'h9696;
    SB_LUT4 i3_2_lut_3_lut_4_lut (.I0(\data_out_frame[20] [2]), .I1(n27138), 
            .I2(n2206), .I3(\data_out_frame[17] [6]), .O(n11_adj_4281));
    defparam i3_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1290 (.I0(n26834), .I1(n27356), .I2(\data_in_frame[4] [4]), 
            .I3(GND_net), .O(n27334));   // verilog/coms.v(75[16:43])
    defparam i2_3_lut_adj_1290.LUT_INIT = 16'h9696;
    SB_LUT4 i1_3_lut_4_lut_adj_1291 (.I0(\FRAME_MATCHER.state[0] ), .I1(n33308), 
            .I2(n73), .I3(n2482), .O(n26472));   // verilog/coms.v(127[12] 300[6])
    defparam i1_3_lut_4_lut_adj_1291.LUT_INIT = 16'hff10;
    SB_LUT4 add_3971_7_lut (.I0(GND_net), .I1(byte_transmit_counter[5]), 
            .I2(GND_net), .I3(n39110), .O(n8825[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_3971_7 (.CI(n39110), .I0(byte_transmit_counter[5]), .I1(GND_net), 
            .CO(n39111));
    SB_LUT4 i1_2_lut_adj_1292 (.I0(\data_in_frame[2] [1]), .I1(\data_in_frame[3] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4282));   // verilog/coms.v(70[16:69])
    defparam i1_2_lut_adj_1292.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1293 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[4] [1]), 
            .I2(\data_in_frame[4] [2]), .I3(n6_adj_4282), .O(n44190));   // verilog/coms.v(70[16:69])
    defparam i4_4_lut_adj_1293.LUT_INIT = 16'h6996;
    SB_LUT4 i15303_3_lut_4_lut (.I0(n34417), .I1(n44095), .I2(rx_data[5]), 
            .I3(\data_in_frame[15] [5]), .O(n28366));
    defparam i15303_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i1_2_lut_adj_1294 (.I0(\data_in_frame[2] [0]), .I1(n44190), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4283));   // verilog/coms.v(78[16:27])
    defparam i1_2_lut_adj_1294.LUT_INIT = 16'h6666;
    SB_LUT4 i15304_3_lut_4_lut (.I0(n34417), .I1(n44095), .I2(rx_data[4]), 
            .I3(\data_in_frame[15] [4]), .O(n28367));
    defparam i15304_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i4_4_lut_adj_1295 (.I0(\data_in_frame[3] [6]), .I1(n27360), 
            .I2(\data_in_frame[1] [4]), .I3(n6_adj_4283), .O(n27394));   // verilog/coms.v(78[16:27])
    defparam i4_4_lut_adj_1295.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1296 (.I0(\data_in_frame[6] [1]), .I1(n26938), 
            .I2(n26978), .I3(\data_in_frame[6] [4]), .O(n44336));   // verilog/coms.v(85[17:28])
    defparam i3_4_lut_adj_1296.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1297 (.I0(Kp_23__N_1095), .I1(n41569), .I2(\data_in_frame[8] [6]), 
            .I3(\data_in_frame[7] [7]), .O(n24_adj_4284));
    defparam i8_4_lut_adj_1297.LUT_INIT = 16'hde7b;
    SB_LUT4 i5_4_lut_adj_1298 (.I0(n44336), .I1(n44360), .I2(n27394), 
            .I3(n44294), .O(n12_adj_4285));   // verilog/coms.v(85[17:28])
    defparam i5_4_lut_adj_1298.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1299 (.I0(Kp_23__N_836), .I1(n12_adj_4285), .I2(n44639), 
            .I3(\data_in_frame[8] [1]), .O(n45516));   // verilog/coms.v(85[17:28])
    defparam i6_4_lut_adj_1299.LUT_INIT = 16'h6996;
    SB_LUT4 i12_3_lut (.I0(n44412), .I1(n24_adj_4284), .I2(n41445), .I3(GND_net), 
            .O(n28_adj_4286));
    defparam i12_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i10_4_lut_adj_1300 (.I0(n41474), .I1(n8_adj_4278), .I2(n27023), 
            .I3(n27414), .O(n26_adj_4287));
    defparam i10_4_lut_adj_1300.LUT_INIT = 16'hffef;
    SB_LUT4 i11_4_lut (.I0(n26996), .I1(n45516), .I2(n26966), .I3(n27010), 
            .O(n27_adj_4288));
    defparam i11_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i9_4_lut_adj_1301 (.I0(n27425), .I1(n4_adj_4250), .I2(n27411), 
            .I3(n27058), .O(n25_adj_4289));
    defparam i9_4_lut_adj_1301.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut_adj_1302 (.I0(n25_adj_4289), .I1(n27_adj_4288), .I2(n26_adj_4287), 
            .I3(n28_adj_4286), .O(n31_adj_4279));
    defparam i15_4_lut_adj_1302.LUT_INIT = 16'hfffe;
    SB_LUT4 add_3971_6_lut (.I0(GND_net), .I1(byte_transmit_counter[4]), 
            .I2(GND_net), .I3(n39109), .O(n8825[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_3971_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i5_4_lut_adj_1303 (.I0(\data_in_frame[18] [6]), .I1(n44464), 
            .I2(\data_in_frame[21] [2]), .I3(\data_in_frame[19] [1]), .O(n12_adj_4290));
    defparam i5_4_lut_adj_1303.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1304 (.I0(\data_in_frame[19] [2]), .I1(Kp_23__N_1644), 
            .I2(\data_in_frame[19] [3]), .I3(GND_net), .O(n6_adj_4291));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_1304.LUT_INIT = 16'h9696;
    SB_LUT4 i3_4_lut_adj_1305 (.I0(\data_in_frame[21] [5]), .I1(n44378), 
            .I2(\data_in_frame[19] [4]), .I3(\data_in_frame[19] [3]), .O(n45393));
    defparam i3_4_lut_adj_1305.LUT_INIT = 16'h6996;
    SB_LUT4 i3_3_lut_adj_1306 (.I0(Kp_23__N_1644), .I1(\data_in_frame[21] [3]), 
            .I2(n42418), .I3(GND_net), .O(n8_adj_4292));
    defparam i3_3_lut_adj_1306.LUT_INIT = 16'h6969;
    SB_LUT4 i1_4_lut_adj_1307 (.I0(n45393), .I1(\data_in_frame[21] [4]), 
            .I2(n6_adj_4291), .I3(Kp_23__N_1647), .O(n48487));
    defparam i1_4_lut_adj_1307.LUT_INIT = 16'hd77d;
    SB_LUT4 i1_4_lut_adj_1308 (.I0(\data_in_frame[19] [2]), .I1(n48487), 
            .I2(n8_adj_4292), .I3(\data_in_frame[19] [1]), .O(n48489));
    defparam i1_4_lut_adj_1308.LUT_INIT = 16'hdeed;
    SB_LUT4 i1_4_lut_adj_1309 (.I0(n48489), .I1(\data_in_frame[20] [4]), 
            .I2(n44483), .I3(n44656), .O(n48491));
    defparam i1_4_lut_adj_1309.LUT_INIT = 16'hebbe;
    SB_LUT4 i1_3_lut_adj_1310 (.I0(\data_in_frame[20] [6]), .I1(n44500), 
            .I2(n44691), .I3(GND_net), .O(n44159));
    defparam i1_3_lut_adj_1310.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1311 (.I0(\data_in_frame[19] [0]), .I1(n12_adj_4290), 
            .I2(n44680), .I3(\data_in_frame[16] [5]), .O(n45788));
    defparam i6_4_lut_adj_1311.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1312 (.I0(n44483), .I1(n44691), .I2(\data_in_frame[20] [5]), 
            .I3(GND_net), .O(n45839));
    defparam i2_3_lut_adj_1312.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1313 (.I0(\data_in_frame[19] [4]), .I1(\data_in_frame[21] [6]), 
            .I2(\data_in_frame[19] [5]), .I3(GND_net), .O(n6_adj_4293));
    defparam i2_3_lut_adj_1313.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1314 (.I0(n45839), .I1(n45788), .I2(n44159), 
            .I3(n48491), .O(n48497));
    defparam i1_4_lut_adj_1314.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_3_lut_adj_1315 (.I0(Kp_23__N_761), .I1(\data_in_frame[19] [0]), 
            .I2(\data_in_frame[20] [7]), .I3(GND_net), .O(n48545));
    defparam i1_3_lut_adj_1315.LUT_INIT = 16'h9696;
    SB_LUT4 i1_4_lut_adj_1316 (.I0(n46677), .I1(n48497), .I2(n6_adj_4293), 
            .I3(n42126), .O(n48499));
    defparam i1_4_lut_adj_1316.LUT_INIT = 16'hedde;
    SB_LUT4 i3_4_lut_adj_1317 (.I0(Kp_23__N_1653), .I1(n44291), .I2(\data_in_frame[19] [5]), 
            .I3(\data_in_frame[21] [7]), .O(n46067));   // verilog/coms.v(268[9:85])
    defparam i3_4_lut_adj_1317.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1318 (.I0(\data_out_frame[20] [2]), .I1(n27138), 
            .I2(n2206), .I3(n46491), .O(n44683));
    defparam i1_2_lut_3_lut_4_lut_adj_1318.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1319 (.I0(n45653), .I1(n45673), .I2(n46067), 
            .I3(n48499), .O(n48505));
    defparam i1_4_lut_adj_1319.LUT_INIT = 16'hfff7;
    SB_LUT4 i1_2_lut_adj_1320 (.I0(\data_in_frame[21] [1]), .I1(n44418), 
            .I2(GND_net), .I3(GND_net), .O(n44419));
    defparam i1_2_lut_adj_1320.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1321 (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[21] [0]), 
            .I2(GND_net), .I3(GND_net), .O(n48529));
    defparam i1_2_lut_adj_1321.LUT_INIT = 16'h6666;
    SB_LUT4 i1_4_lut_adj_1322 (.I0(n27297), .I1(n26749), .I2(n26890), 
            .I3(n48529), .O(n48535));
    defparam i1_4_lut_adj_1322.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1323 (.I0(n42281), .I1(n42322), .I2(n44500), 
            .I3(n48545), .O(n46266));
    defparam i1_4_lut_adj_1323.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1324 (.I0(\data_in_frame[20] [1]), .I1(n44419), 
            .I2(n44537), .I3(n48505), .O(n48509));
    defparam i1_4_lut_adj_1324.LUT_INIT = 16'hffde;
    SB_LUT4 i1_4_lut_adj_1325 (.I0(n44291), .I1(n44537), .I2(n44659), 
            .I3(\data_in_frame[20] [0]), .O(n45684));
    defparam i1_4_lut_adj_1325.LUT_INIT = 16'h6996;
    SB_LUT4 i1_4_lut_adj_1326 (.I0(n42442), .I1(n44418), .I2(n44636), 
            .I3(n48535), .O(n45508));
    defparam i1_4_lut_adj_1326.LUT_INIT = 16'h9669;
    SB_LUT4 i1_4_lut_adj_1327 (.I0(n45508), .I1(n45684), .I2(n48509), 
            .I3(n46266), .O(n31_adj_4185));
    defparam i1_4_lut_adj_1327.LUT_INIT = 16'hf7ff;
    SB_LUT4 i15305_3_lut_4_lut (.I0(n34417), .I1(n44095), .I2(rx_data[3]), 
            .I3(\data_in_frame[15] [3]), .O(n28368));
    defparam i15305_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15306_3_lut_4_lut (.I0(n34417), .I1(n44095), .I2(rx_data[2]), 
            .I3(\data_in_frame[15] [2]), .O(n28369));
    defparam i15306_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15421_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44104), .I2(rx_data[7]), 
            .I3(\data_in_frame[0] [7]), .O(n28484));
    defparam i15421_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15422_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44104), .I2(rx_data[6]), 
            .I3(\data_in_frame[0] [6]), .O(n28485));
    defparam i15422_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15307_3_lut_4_lut (.I0(n34417), .I1(n44095), .I2(rx_data[1]), 
            .I3(\data_in_frame[15] [1]), .O(n28370));
    defparam i15307_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i15425_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44104), .I2(rx_data[5]), 
            .I3(\data_in_frame[0] [5]), .O(n28488));
    defparam i15425_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15426_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44104), .I2(rx_data[4]), 
            .I3(\data_in_frame[0] [4]), .O(n28489));
    defparam i15426_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15427_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44104), .I2(rx_data[3]), 
            .I3(\data_in_frame[0] [3]), .O(n28490));
    defparam i15427_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15428_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44104), .I2(rx_data[2]), 
            .I3(\data_in_frame[0] [2]), .O(n28491));
    defparam i15428_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i7390_3_lut (.I0(n31_adj_4185), .I1(n31_adj_4279), .I2(\FRAME_MATCHER.state_c [1]), 
            .I3(GND_net), .O(n23701));   // verilog/coms.v(145[4] 299[11])
    defparam i7390_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15429_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44104), .I2(rx_data[1]), 
            .I3(\data_in_frame[0] [1]), .O(n28492));
    defparam i15429_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i4_4_lut_adj_1328 (.I0(\data_in_frame[0] [4]), .I1(\data_in_frame[0] [6]), 
            .I2(ID[4]), .I3(ID[6]), .O(n12_adj_4294));   // verilog/coms.v(238[12:32])
    defparam i4_4_lut_adj_1328.LUT_INIT = 16'h7bde;
    SB_LUT4 i15149_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44104), .I2(rx_data[0]), 
            .I3(\data_in_frame[0] [0]), .O(n28212));
    defparam i15149_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_4_lut_adj_1329 (.I0(\data_in_frame[0] [1]), .I1(\data_in_frame[0] [2]), 
            .I2(ID[1]), .I3(ID[2]), .O(n10_adj_4295));   // verilog/coms.v(238[12:32])
    defparam i2_4_lut_adj_1329.LUT_INIT = 16'h7bde;
    SB_LUT4 i2_3_lut_4_lut_adj_1330 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n33565), .O(n44095));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1330.LUT_INIT = 16'hefff;
    SB_LUT4 i2_3_lut_4_lut_adj_1331 (.I0(\FRAME_MATCHER.i [4]), .I1(\FRAME_MATCHER.i [5]), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n33565), .O(n44104));   // verilog/coms.v(154[7:23])
    defparam i2_3_lut_4_lut_adj_1331.LUT_INIT = 16'hfeff;
    SB_LUT4 i15308_3_lut_4_lut (.I0(n34417), .I1(n44095), .I2(rx_data[0]), 
            .I3(\data_in_frame[15] [0]), .O(n28371));
    defparam i15308_3_lut_4_lut.LUT_INIT = 16'hfd20;
    SB_LUT4 i3_4_lut_adj_1332 (.I0(\data_in_frame[0] [7]), .I1(\data_in_frame[0] [5]), 
            .I2(ID[7]), .I3(ID[5]), .O(n11_adj_4296));   // verilog/coms.v(238[12:32])
    defparam i3_4_lut_adj_1332.LUT_INIT = 16'h7bde;
    SB_LUT4 i1_4_lut_adj_1333 (.I0(\data_in_frame[0] [0]), .I1(\data_in_frame[0] [3]), 
            .I2(ID[0]), .I3(ID[3]), .O(n9_adj_4297));   // verilog/coms.v(238[12:32])
    defparam i1_4_lut_adj_1333.LUT_INIT = 16'h7bde;
    SB_LUT4 i7_4_lut_adj_1334 (.I0(n9_adj_4297), .I1(n11_adj_4296), .I2(n10_adj_4295), 
            .I3(n12_adj_4294), .O(n24120));   // verilog/coms.v(238[12:32])
    defparam i7_4_lut_adj_1334.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_adj_1335 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state [3]), 
            .I2(GND_net), .I3(GND_net), .O(n48623));
    defparam i1_2_lut_adj_1335.LUT_INIT = 16'heeee;
    SB_LUT4 i1_4_lut_adj_1336 (.I0(\FRAME_MATCHER.state_c [2]), .I1(n34355), 
            .I2(n34549), .I3(n48623), .O(n48629));
    defparam i1_4_lut_adj_1336.LUT_INIT = 16'hfffd;
    SB_LUT4 i35744_4_lut (.I0(n24120), .I1(n23701), .I2(n34685), .I3(n48629), 
            .O(n27781));
    defparam i35744_4_lut.LUT_INIT = 16'h0001;
    SB_LUT4 mux_1361_i1_3_lut (.I0(\data_in_frame[19] [0]), .I1(\data_in_frame[3] [0]), 
            .I2(n5785), .I3(GND_net), .O(n5786));
    defparam mux_1361_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i5_3_lut_4_lut_adj_1337 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(n10_adj_4124), .I3(n27269), .O(n44304));   // verilog/coms.v(85[17:70])
    defparam i5_3_lut_4_lut_adj_1337.LUT_INIT = 16'h6996;
    SB_LUT4 i1_3_lut_4_lut_adj_1338 (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(n26770), .I3(\data_in_frame[5] [0]), .O(n44251));
    defparam i1_3_lut_4_lut_adj_1338.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1339 (.I0(\data_out_frame[7] [7]), .I1(\data_out_frame[7] [6]), 
            .I2(\data_out_frame[8] [0]), .I3(GND_net), .O(n44606));   // verilog/coms.v(85[17:70])
    defparam i1_2_lut_3_lut_adj_1339.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1340 (.I0(n44439), .I1(\data_in_frame[12] [4]), 
            .I2(\data_in_frame[14] [6]), .I3(GND_net), .O(n44763));
    defparam i1_2_lut_3_lut_adj_1340.LUT_INIT = 16'h9696;
    SB_LUT4 i15293_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44085), .I2(rx_data[7]), 
            .I3(\data_in_frame[16] [7]), .O(n28356));
    defparam i15293_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15294_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44085), .I2(rx_data[6]), 
            .I3(\data_in_frame[16] [6]), .O(n28357));
    defparam i15294_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_3_lut_4_lut_adj_1341 (.I0(n23831), .I1(n2482), .I2(n61), 
            .I3(n76), .O(n43975));
    defparam i2_3_lut_4_lut_adj_1341.LUT_INIT = 16'h0200;
    SB_LUT4 i2_3_lut_4_lut_adj_1342 (.I0(n23831), .I1(n2482), .I2(n33302), 
            .I3(n76), .O(n44042));
    defparam i2_3_lut_4_lut_adj_1342.LUT_INIT = 16'h2000;
    SB_LUT4 i30097_2_lut_3_lut (.I0(n34823), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n44977), .I3(GND_net), .O(n44989));
    defparam i30097_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i35851_2_lut_3_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state_c [2]), 
            .I2(\FRAME_MATCHER.state[0] ), .I3(GND_net), .O(n44_adj_4244));
    defparam i35851_2_lut_3_lut.LUT_INIT = 16'h0e0e;
    SB_LUT4 i1_2_lut_3_lut_adj_1343 (.I0(n63_adj_4138), .I1(n63_c), .I2(\FRAME_MATCHER.state_c [1]), 
            .I3(GND_net), .O(n39));   // verilog/coms.v(136[7:86])
    defparam i1_2_lut_3_lut_adj_1343.LUT_INIT = 16'h8080;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36494 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18] [3]), .I2(\data_out_frame[19] [3]), 
            .I3(byte_transmit_counter[1]), .O(n51447));
    defparam byte_transmit_counter_0__bdd_4_lut_36494.LUT_INIT = 16'he4aa;
    SB_LUT4 i1_2_lut_3_lut_adj_1344 (.I0(n63_adj_4138), .I1(n63_c), .I2(n63), 
            .I3(GND_net), .O(n23831));   // verilog/coms.v(136[7:86])
    defparam i1_2_lut_3_lut_adj_1344.LUT_INIT = 16'h8080;
    SB_LUT4 i2_3_lut_4_lut_adj_1345 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(\FRAME_MATCHER.state_c [2]), .I3(n67), .O(n69));
    defparam i2_3_lut_4_lut_adj_1345.LUT_INIT = 16'h5400;
    SB_LUT4 n51447_bdd_4_lut (.I0(n51447), .I1(\data_out_frame[17] [3]), 
            .I2(\data_out_frame[16] [3]), .I3(byte_transmit_counter[1]), 
            .O(n51450));
    defparam n51447_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i3_4_lut_adj_1346 (.I0(\FRAME_MATCHER.state_c [7]), .I1(\FRAME_MATCHER.state_c [6]), 
            .I2(\FRAME_MATCHER.state_c [4]), .I3(\FRAME_MATCHER.state_c [5]), 
            .O(n34355));
    defparam i3_4_lut_adj_1346.LUT_INIT = 16'hfffe;
    SB_LUT4 i15295_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44085), .I2(rx_data[5]), 
            .I3(\data_in_frame[16] [5]), .O(n28358));
    defparam i15295_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15296_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44085), .I2(rx_data[4]), 
            .I3(\data_in_frame[16] [4]), .O(n28359));
    defparam i15296_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15297_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44085), .I2(rx_data[3]), 
            .I3(\data_in_frame[16] [3]), .O(n28360));
    defparam i15297_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15298_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44085), .I2(rx_data[2]), 
            .I3(\data_in_frame[16] [2]), .O(n28361));
    defparam i15298_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1347 (.I0(\FRAME_MATCHER.i [4]), .I1(n26686), 
            .I2(\FRAME_MATCHER.i [1]), .I3(\FRAME_MATCHER.i [0]), .O(n5_adj_4150));   // verilog/coms.v(154[7:23])
    defparam i1_3_lut_4_lut_adj_1347.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_3_lut_4_lut_adj_1348 (.I0(\FRAME_MATCHER.i [4]), .I1(n26686), 
            .I2(\FRAME_MATCHER.i [3]), .I3(n8_adj_4134), .O(n26489));   // verilog/coms.v(154[7:23])
    defparam i1_3_lut_4_lut_adj_1348.LUT_INIT = 16'hfeee;
    SB_LUT4 equal_124_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4141));   // verilog/coms.v(154[7:23])
    defparam equal_124_i8_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i2_2_lut_3_lut_adj_1349 (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4134));   // verilog/coms.v(154[7:23])
    defparam i2_2_lut_3_lut_adj_1349.LUT_INIT = 16'hfefe;
    SB_LUT4 i8_4_lut_adj_1350 (.I0(\FRAME_MATCHER.state_c [16]), .I1(\FRAME_MATCHER.state_c [17]), 
            .I2(\FRAME_MATCHER.state_c [26]), .I3(\FRAME_MATCHER.state_c [18]), 
            .O(n20_adj_4299));   // verilog/coms.v(231[5:23])
    defparam i8_4_lut_adj_1350.LUT_INIT = 16'hfffe;
    SB_LUT4 i15299_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44085), .I2(rx_data[1]), 
            .I3(\data_in_frame[16] [1]), .O(n28362));
    defparam i15299_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1351 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [4]), 
            .I3(GND_net), .O(n43589));
    defparam i1_2_lut_3_lut_adj_1351.LUT_INIT = 16'he0e0;
    SB_LUT4 i15300_3_lut_4_lut (.I0(n8_adj_4134), .I1(n44085), .I2(rx_data[0]), 
            .I3(\data_in_frame[16] [0]), .O(n28363));
    defparam i15300_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1352 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [5]), 
            .I3(GND_net), .O(n43591));
    defparam i1_2_lut_3_lut_adj_1352.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1353 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [6]), 
            .I3(GND_net), .O(n43593));
    defparam i1_2_lut_3_lut_adj_1353.LUT_INIT = 16'he0e0;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36489 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18][2] ), .I2(\data_out_frame[19] [2]), 
            .I3(byte_transmit_counter[1]), .O(n51441));
    defparam byte_transmit_counter_0__bdd_4_lut_36489.LUT_INIT = 16'he4aa;
    SB_LUT4 i2_3_lut_adj_1354 (.I0(byte_transmit_counter[7]), .I1(byte_transmit_counter[6]), 
            .I2(byte_transmit_counter[5]), .I3(GND_net), .O(n6_adj_4242));
    defparam i2_3_lut_adj_1354.LUT_INIT = 16'hfefe;
    SB_LUT4 i21348_2_lut (.I0(\byte_transmit_counter[0] ), .I1(byte_transmit_counter[1]), 
            .I2(GND_net), .I3(GND_net), .O(n34409));
    defparam i21348_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i2_4_lut_adj_1355 (.I0(byte_transmit_counter[3]), .I1(byte_transmit_counter[4]), 
            .I2(n34409), .I3(\byte_transmit_counter[2] ), .O(n34527));
    defparam i2_4_lut_adj_1355.LUT_INIT = 16'h8880;
    SB_LUT4 i1_2_lut_3_lut_adj_1356 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [7]), 
            .I3(GND_net), .O(n43595));
    defparam i1_2_lut_3_lut_adj_1356.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1357 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [8]), 
            .I3(GND_net), .O(n43597));
    defparam i1_2_lut_3_lut_adj_1357.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1358 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [9]), 
            .I3(GND_net), .O(n43599));
    defparam i1_2_lut_3_lut_adj_1358.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_adj_1359 (.I0(n34355), .I1(n34685), .I2(n34549), 
            .I3(GND_net), .O(n44929));
    defparam i2_3_lut_adj_1359.LUT_INIT = 16'hfefe;
    SB_LUT4 i30087_3_lut (.I0(\FRAME_MATCHER.state [3]), .I1(n44929), .I2(n34047), 
            .I3(GND_net), .O(n44977));
    defparam i30087_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 n51441_bdd_4_lut (.I0(n51441), .I1(\data_out_frame[17] [2]), 
            .I2(\data_out_frame[16] [2]), .I3(byte_transmit_counter[1]), 
            .O(n51444));
    defparam n51441_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_adj_1360 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [10]), 
            .I3(GND_net), .O(n43601));
    defparam i1_2_lut_3_lut_adj_1360.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1361 (.I0(\data_out_frame[8] [5]), .I1(n26712), 
            .I2(\data_out_frame[8] [6]), .I3(GND_net), .O(n44570));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1361.LUT_INIT = 16'h9696;
    SB_LUT4 i7_4_lut_adj_1362 (.I0(\FRAME_MATCHER.state_c [28]), .I1(\FRAME_MATCHER.state_c [22]), 
            .I2(\FRAME_MATCHER.state_c [21]), .I3(\FRAME_MATCHER.state_c [20]), 
            .O(n19_adj_4300));   // verilog/coms.v(231[5:23])
    defparam i7_4_lut_adj_1362.LUT_INIT = 16'hfffe;
    SB_LUT4 i3_4_lut_adj_1363 (.I0(n34527), .I1(n6_adj_4242), .I2(n40), 
            .I3(n44035), .O(n46506));
    defparam i3_4_lut_adj_1363.LUT_INIT = 16'hfeff;
    SB_LUT4 mux_870_i1_3_lut (.I0(n46506), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n34823), .I3(GND_net), .O(n3912[0]));   // verilog/coms.v(145[4] 299[11])
    defparam mux_870_i1_3_lut.LUT_INIT = 16'h5c5c;
    SB_LUT4 i1_2_lut_3_lut_adj_1364 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [11]), 
            .I3(GND_net), .O(n43603));
    defparam i1_2_lut_3_lut_adj_1364.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1365 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [12]), 
            .I3(GND_net), .O(n43605));
    defparam i1_2_lut_3_lut_adj_1365.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1366 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [13]), 
            .I3(GND_net), .O(n43607));
    defparam i1_2_lut_3_lut_adj_1366.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1367 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [14]), 
            .I3(GND_net), .O(n43609));
    defparam i1_2_lut_3_lut_adj_1367.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_2_lut_3_lut_adj_1368 (.I0(\data_out_frame[8] [5]), .I1(n26712), 
            .I2(n27407), .I3(GND_net), .O(n27403));   // verilog/coms.v(75[16:43])
    defparam i2_2_lut_3_lut_adj_1368.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1369 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [15]), 
            .I3(GND_net), .O(n43611));
    defparam i1_2_lut_3_lut_adj_1369.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1370 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [16]), 
            .I3(GND_net), .O(n43613));
    defparam i1_2_lut_3_lut_adj_1370.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_2_lut_3_lut_4_lut (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(\data_out_frame[9] [7]), .I3(\data_out_frame[4] [7]), .O(n10_adj_4120));   // verilog/coms.v(73[16:34])
    defparam i2_2_lut_3_lut_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1371 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [17]), 
            .I3(GND_net), .O(n43615));
    defparam i1_2_lut_3_lut_adj_1371.LUT_INIT = 16'he0e0;
    SB_LUT4 i33980_3_lut (.I0(\data_out_frame[6] [3]), .I1(\data_out_frame[7] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48932));
    defparam i33980_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1372 (.I0(n33298), .I1(\FRAME_MATCHER.state [3]), 
            .I2(n44055), .I3(GND_net), .O(n4_adj_4169));
    defparam i1_2_lut_3_lut_adj_1372.LUT_INIT = 16'h1010;
    SB_LUT4 i33981_4_lut (.I0(n48932), .I1(byte_transmit_counter[1]), .I2(\byte_transmit_counter[2] ), 
            .I3(\byte_transmit_counter[0] ), .O(n48933));
    defparam i33981_4_lut.LUT_INIT = 16'hafa3;
    SB_LUT4 i1_2_lut_3_lut_adj_1373 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [18]), 
            .I3(GND_net), .O(n43617));
    defparam i1_2_lut_3_lut_adj_1373.LUT_INIT = 16'he0e0;
    SB_LUT4 i33979_3_lut (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[5] [3]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48931));
    defparam i33979_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i20522_2_lut_3_lut (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [19]), 
            .I3(GND_net), .O(n33568));
    defparam i20522_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1374 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [20]), 
            .I3(GND_net), .O(n43619));
    defparam i1_2_lut_3_lut_adj_1374.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_3_lut_4_lut_adj_1375 (.I0(n26489), .I1(\FRAME_MATCHER.i[31] ), 
            .I2(\FRAME_MATCHER.i_31__N_2524 ), .I3(n23831), .O(n4_c));
    defparam i1_3_lut_4_lut_adj_1375.LUT_INIT = 16'hd000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_1376 (.I0(\data_out_frame[5] [2]), .I1(\data_out_frame[5] [1]), 
            .I2(n44712), .I3(\data_out_frame[4] [7]), .O(n6_adj_4114));   // verilog/coms.v(73[16:34])
    defparam i1_2_lut_3_lut_4_lut_adj_1376.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1377 (.I0(\FRAME_MATCHER.state_c [27]), .I1(\FRAME_MATCHER.state_c [30]), 
            .I2(\FRAME_MATCHER.state_c [29]), .I3(\FRAME_MATCHER.state_c [23]), 
            .O(n42170));   // verilog/coms.v(127[12] 300[6])
    defparam i3_4_lut_adj_1377.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_3_lut_adj_1378 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [21]), 
            .I3(GND_net), .O(n7_adj_4189));
    defparam i1_2_lut_3_lut_adj_1378.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1379 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [22]), 
            .I3(GND_net), .O(n7_adj_4187));
    defparam i1_2_lut_3_lut_adj_1379.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1380 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [23]), 
            .I3(GND_net), .O(n43621));
    defparam i1_2_lut_3_lut_adj_1380.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut_adj_1381 (.I0(\FRAME_MATCHER.state[0] ), .I1(\FRAME_MATCHER.state_c [1]), 
            .I2(n33298), .I3(\FRAME_MATCHER.state [3]), .O(n33307));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_4_lut_adj_1381.LUT_INIT = 16'hfffb;
    SB_LUT4 i1_2_lut_3_lut_adj_1382 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [24]), 
            .I3(GND_net), .O(n43623));
    defparam i1_2_lut_3_lut_adj_1382.LUT_INIT = 16'he0e0;
    SB_LUT4 i20524_2_lut_3_lut (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [25]), 
            .I3(GND_net), .O(n33572));
    defparam i20524_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_3_lut_adj_1383 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [26]), 
            .I3(GND_net), .O(n43625));
    defparam i1_2_lut_3_lut_adj_1383.LUT_INIT = 16'he0e0;
    SB_LUT4 i20525_2_lut_3_lut (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [27]), 
            .I3(GND_net), .O(n33574));
    defparam i20525_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i15285_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44085), .I2(rx_data[7]), 
            .I3(\data_in_frame[17] [7]), .O(n28348));
    defparam i15285_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1384 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [28]), 
            .I3(GND_net), .O(n43627));
    defparam i1_2_lut_3_lut_adj_1384.LUT_INIT = 16'he0e0;
    SB_LUT4 i15286_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44085), .I2(rx_data[6]), 
            .I3(\data_in_frame[17] [6]), .O(n28349));
    defparam i15286_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_4_lut_adj_1385 (.I0(\FRAME_MATCHER.state_c [31]), .I1(\FRAME_MATCHER.state_c [19]), 
            .I2(\FRAME_MATCHER.state_c [24]), .I3(\FRAME_MATCHER.state_c [25]), 
            .O(n21_adj_4301));   // verilog/coms.v(231[5:23])
    defparam i9_4_lut_adj_1385.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_4_lut_adj_1386 (.I0(n21_adj_4301), .I1(n42170), .I2(n19_adj_4300), 
            .I3(n20_adj_4299), .O(n34685));
    defparam i1_4_lut_adj_1386.LUT_INIT = 16'hfffe;
    SB_LUT4 i20526_2_lut_3_lut (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [29]), 
            .I3(GND_net), .O(n33576));
    defparam i20526_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_3_lut_4_lut_adj_1387 (.I0(n26687), .I1(\FRAME_MATCHER.i[31] ), 
            .I2(\FRAME_MATCHER.i_31__N_2526 ), .I3(n23831), .O(n72));   // verilog/coms.v(254[5:25])
    defparam i1_3_lut_4_lut_adj_1387.LUT_INIT = 16'hd000;
    SB_LUT4 i1_2_lut_3_lut_adj_1388 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [30]), 
            .I3(GND_net), .O(n7_adj_4183));
    defparam i1_2_lut_3_lut_adj_1388.LUT_INIT = 16'he0e0;
    SB_LUT4 i2_3_lut_4_lut_adj_1389 (.I0(n46253), .I1(n42300), .I2(\data_out_frame[23] [0]), 
            .I3(\data_out_frame[23] [1]), .O(n44518));
    defparam i2_3_lut_4_lut_adj_1389.LUT_INIT = 16'h9669;
    SB_LUT4 i330_2_lut_4_lut (.I0(n34527), .I1(n6_adj_4242), .I2(r_SM_Main_2__N_3516[0]), 
            .I3(tx_active), .O(n1476));   // verilog/coms.v(213[6] 220[9])
    defparam i330_2_lut_4_lut.LUT_INIT = 16'hfff1;
    SB_LUT4 i15287_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44085), .I2(rx_data[5]), 
            .I3(\data_in_frame[17] [5]), .O(n28350));
    defparam i15287_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1390 (.I0(n68), .I1(n72), .I2(\FRAME_MATCHER.state_c [31]), 
            .I3(GND_net), .O(n43587));
    defparam i1_2_lut_3_lut_adj_1390.LUT_INIT = 16'he0e0;
    SB_LUT4 i15288_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44085), .I2(rx_data[4]), 
            .I3(\data_in_frame[17] [4]), .O(n28351));
    defparam i15288_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i35045_2_lut (.I0(n51564), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n49808));
    defparam i35045_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i33947_4_lut (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[23] [3]), 
            .I2(byte_transmit_counter[1]), .I3(\byte_transmit_counter[0] ), 
            .O(n48899));
    defparam i33947_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i35346_3_lut (.I0(n51450), .I1(n48899), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n50299));
    defparam i35346_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_adj_1391 (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n6014));
    defparam i1_2_lut_3_lut_adj_1391.LUT_INIT = 16'h0202;
    SB_LUT4 i1_2_lut_adj_1392 (.I0(n33298), .I1(\FRAME_MATCHER.state [3]), 
            .I2(GND_net), .I3(GND_net), .O(n33308));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_adj_1392.LUT_INIT = 16'heeee;
    SB_LUT4 i33974_3_lut (.I0(\data_out_frame[6] [2]), .I1(\data_out_frame[7] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48926));
    defparam i33974_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i33975_4_lut (.I0(n48926), .I1(\byte_transmit_counter[0] ), 
            .I2(\byte_transmit_counter[2] ), .I3(byte_transmit_counter[1]), 
            .O(n48927));
    defparam i33975_4_lut.LUT_INIT = 16'ha0a3;
    SB_LUT4 i35966_2_lut (.I0(\FRAME_MATCHER.state_c [1]), .I1(\FRAME_MATCHER.state_c [2]), 
            .I2(GND_net), .I3(GND_net), .O(n73));
    defparam i35966_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 i33973_3_lut (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[5] [2]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48925));
    defparam i33973_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35043_2_lut (.I0(n51570), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n49811));
    defparam i35043_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15289_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44085), .I2(rx_data[3]), 
            .I3(\data_in_frame[17] [3]), .O(n28352));
    defparam i15289_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15290_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44085), .I2(rx_data[2]), 
            .I3(\data_in_frame[17] [2]), .O(n28353));
    defparam i15290_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1393 (.I0(n46253), .I1(n42300), .I2(\data_out_frame[24] [7]), 
            .I3(GND_net), .O(n42438));
    defparam i1_2_lut_3_lut_adj_1393.LUT_INIT = 16'h6969;
    SB_LUT4 i15291_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44085), .I2(rx_data[1]), 
            .I3(\data_in_frame[17] [1]), .O(n28354));
    defparam i15291_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15292_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44085), .I2(rx_data[0]), 
            .I3(\data_in_frame[17] [0]), .O(n28355));
    defparam i15292_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i33944_4_lut (.I0(\data_out_frame[20] [2]), .I1(\data_out_frame[23] [2]), 
            .I2(byte_transmit_counter[1]), .I3(\byte_transmit_counter[0] ), 
            .O(n48896));
    defparam i33944_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i35350_3_lut (.I0(n51444), .I1(n48896), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n50303));
    defparam i35350_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15277_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44085), .I2(rx_data[7]), 
            .I3(\data_in_frame[18] [7]), .O(n28340));
    defparam i15277_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i35987_3_lut_4_lut (.I0(n33302), .I1(n76), .I2(r_SM_Main_2__N_3516[0]), 
            .I3(tx_active), .O(n27787));
    defparam i35987_3_lut_4_lut.LUT_INIT = 16'h3337;
    SB_LUT4 i1_2_lut_3_lut_adj_1394 (.I0(n44035), .I1(n33298), .I2(\FRAME_MATCHER.state [3]), 
            .I3(GND_net), .O(n33302));   // verilog/coms.v(127[12] 300[6])
    defparam i1_2_lut_3_lut_adj_1394.LUT_INIT = 16'hfdfd;
    SB_LUT4 i33966_4_lut (.I0(\data_out_frame[6] [1]), .I1(\byte_transmit_counter[0] ), 
            .I2(\byte_transmit_counter[2] ), .I3(\data_out_frame[7] [1]), 
            .O(n48918));
    defparam i33966_4_lut.LUT_INIT = 16'hec2c;
    SB_LUT4 i33964_3_lut (.I0(\data_out_frame[4] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(\byte_transmit_counter[0] ), .I3(GND_net), .O(n48916));
    defparam i33964_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35040_2_lut (.I0(n51576), .I1(\byte_transmit_counter[2] ), 
            .I2(GND_net), .I3(GND_net), .O(n49814));
    defparam i35040_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i33941_4_lut (.I0(\data_out_frame[20] [1]), .I1(\data_out_frame[23] [1]), 
            .I2(byte_transmit_counter[1]), .I3(\byte_transmit_counter[0] ), 
            .O(n48893));
    defparam i33941_4_lut.LUT_INIT = 16'hc00a;
    SB_LUT4 i35352_3_lut (.I0(n51438), .I1(n48893), .I2(\byte_transmit_counter[2] ), 
            .I3(GND_net), .O(n50305));
    defparam i35352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i15278_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44085), .I2(rx_data[6]), 
            .I3(\data_in_frame[18] [6]), .O(n28341));
    defparam i15278_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36484 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18]_c [1]), .I2(\data_out_frame[19] [1]), 
            .I3(byte_transmit_counter[1]), .O(n51435));
    defparam byte_transmit_counter_0__bdd_4_lut_36484.LUT_INIT = 16'he4aa;
    SB_LUT4 i15279_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44085), .I2(rx_data[5]), 
            .I3(\data_in_frame[18] [5]), .O(n28342));
    defparam i15279_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_3_lut_4_lut_adj_1395 (.I0(\FRAME_MATCHER.state_c [30]), .I1(n6_adj_4135), 
            .I2(n4_c), .I3(n1), .O(n43477));
    defparam i1_3_lut_4_lut_adj_1395.LUT_INIT = 16'haaa8;
    SB_LUT4 i15280_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44085), .I2(rx_data[4]), 
            .I3(\data_in_frame[18] [4]), .O(n28343));
    defparam i15280_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i86_3_lut_4_lut (.I0(n68), .I1(\FRAME_MATCHER.state [3]), .I2(n4_c), 
            .I3(n1), .O(n81));
    defparam i86_3_lut_4_lut.LUT_INIT = 16'hccc8;
    SB_LUT4 equal_1543_i7_2_lut_3_lut (.I0(\data_in_frame[0] [5]), .I1(\data_in_frame[0] [4]), 
            .I2(\data_in_frame[2] [6]), .I3(GND_net), .O(n7_c));   // verilog/coms.v(166[9:87])
    defparam equal_1543_i7_2_lut_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i15413_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44104), .I2(rx_data[7]), 
            .I3(\data_in_frame[1] [7]), .O(n28476));
    defparam i15413_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15414_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44104), .I2(rx_data[6]), 
            .I3(\data_in_frame[1] [6]), .O(n28477));
    defparam i15414_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15281_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44085), .I2(rx_data[3]), 
            .I3(\data_in_frame[18] [3]), .O(n28344));
    defparam i15281_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15415_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44104), .I2(rx_data[5]), 
            .I3(\data_in_frame[1] [5]), .O(n28478));
    defparam i15415_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15416_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44104), .I2(rx_data[4]), 
            .I3(\data_in_frame[1] [4]), .O(n28479));
    defparam i15416_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 n51435_bdd_4_lut (.I0(n51435), .I1(\data_out_frame[17] [1]), 
            .I2(\data_out_frame[16] [1]), .I3(byte_transmit_counter[1]), 
            .O(n51438));
    defparam n51435_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i15417_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44104), .I2(rx_data[3]), 
            .I3(\data_in_frame[1] [3]), .O(n28480));
    defparam i15417_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15418_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44104), .I2(rx_data[2]), 
            .I3(\data_in_frame[1] [2]), .O(n28481));
    defparam i15418_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15419_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44104), .I2(rx_data[1]), 
            .I3(\data_in_frame[1] [1]), .O(n28482));
    defparam i15419_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15420_3_lut_4_lut (.I0(n8_adj_4141), .I1(n44104), .I2(rx_data[0]), 
            .I3(\data_in_frame[1] [0]), .O(n28483));
    defparam i15420_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15282_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44085), .I2(rx_data[2]), 
            .I3(\data_in_frame[18] [2]), .O(n28345));
    defparam i15282_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i21305_2_lut_3_lut (.I0(n58), .I1(n44113), .I2(\FRAME_MATCHER.state_c [19]), 
            .I3(GND_net), .O(n34362));
    defparam i21305_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i21306_2_lut_3_lut (.I0(n58), .I1(n44113), .I2(\FRAME_MATCHER.state_c [25]), 
            .I3(GND_net), .O(n34364));
    defparam i21306_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i21307_2_lut_3_lut (.I0(n58), .I1(n44113), .I2(\FRAME_MATCHER.state_c [27]), 
            .I3(GND_net), .O(n34366));
    defparam i21307_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i21308_2_lut_3_lut (.I0(n58), .I1(n44113), .I2(\FRAME_MATCHER.state_c [29]), 
            .I3(GND_net), .O(n34368));
    defparam i21308_2_lut_3_lut.LUT_INIT = 16'he0e0;
    SB_LUT4 i1_2_lut_4_lut_adj_1396 (.I0(n26473), .I1(n44079), .I2(n44055), 
            .I3(\FRAME_MATCHER.state_c [4]), .O(n43491));
    defparam i1_2_lut_4_lut_adj_1396.LUT_INIT = 16'hdc00;
    SB_LUT4 i15283_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44085), .I2(rx_data[1]), 
            .I3(\data_in_frame[18] [1]), .O(n28346));
    defparam i15283_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1397 (.I0(n26473), .I1(n44079), .I2(n44055), 
            .I3(\FRAME_MATCHER.state_c [24]), .O(n43515));
    defparam i1_2_lut_4_lut_adj_1397.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1398 (.I0(n26473), .I1(n44079), .I2(n44055), 
            .I3(\FRAME_MATCHER.state_c [26]), .O(n43513));
    defparam i1_2_lut_4_lut_adj_1398.LUT_INIT = 16'hdc00;
    SB_LUT4 i1_2_lut_4_lut_adj_1399 (.I0(n26473), .I1(n44079), .I2(n44055), 
            .I3(\FRAME_MATCHER.state_c [28]), .O(n43511));
    defparam i1_2_lut_4_lut_adj_1399.LUT_INIT = 16'hdc00;
    SB_LUT4 i15405_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44104), .I2(rx_data[7]), 
            .I3(\data_in_frame[2] [7]), .O(n28468));
    defparam i15405_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15406_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44104), .I2(rx_data[6]), 
            .I3(\data_in_frame[2] [6]), .O(n28469));
    defparam i15406_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15407_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44104), .I2(rx_data[5]), 
            .I3(\data_in_frame[2] [5]), .O(n28470));
    defparam i15407_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15408_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44104), .I2(rx_data[4]), 
            .I3(\data_in_frame[2] [4]), .O(n28471));
    defparam i15408_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15284_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44085), .I2(rx_data[0]), 
            .I3(\data_in_frame[18] [0]), .O(n28347));
    defparam i15284_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 equal_127_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(GND_net), .O(n8_adj_4232));   // verilog/coms.v(154[7:23])
    defparam equal_127_i8_2_lut_3_lut.LUT_INIT = 16'hbfbf;
    SB_LUT4 i15409_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44104), .I2(rx_data[3]), 
            .I3(\data_in_frame[2] [3]), .O(n28472));
    defparam i15409_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15410_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44104), .I2(rx_data[2]), 
            .I3(\data_in_frame[2] [2]), .O(n28473));
    defparam i15410_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1400 (.I0(n44255), .I1(\data_out_frame[14] [4]), 
            .I2(\data_out_frame[12] [2]), .I3(n41455), .O(n41486));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1400.LUT_INIT = 16'h6996;
    SB_LUT4 i15411_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44104), .I2(rx_data[1]), 
            .I3(\data_in_frame[2] [1]), .O(n28474));
    defparam i15411_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1401 (.I0(n44255), .I1(\data_out_frame[14] [4]), 
            .I2(\data_out_frame[12] [2]), .I3(n27220), .O(n1794));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1401.LUT_INIT = 16'h6996;
    SB_LUT4 i15412_3_lut_4_lut (.I0(n8_adj_4142), .I1(n44104), .I2(rx_data[0]), 
            .I3(\data_in_frame[2] [0]), .O(n28475));
    defparam i15412_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i20523_2_lut_4_lut (.I0(n1), .I1(n58), .I2(n4_c), .I3(\FRAME_MATCHER.state_c [21]), 
            .O(n33570));   // verilog/coms.v(115[11:12])
    defparam i20523_2_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 i21356_2_lut_3_lut (.I0(\FRAME_MATCHER.i [0]), .I1(\FRAME_MATCHER.i [1]), 
            .I2(\FRAME_MATCHER.i [2]), .I3(GND_net), .O(n34417));
    defparam i21356_2_lut_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_4_lut_adj_1402 (.I0(n1), .I1(n58), .I2(n4_c), .I3(\FRAME_MATCHER.state_c [22]), 
            .O(n8_adj_4188));   // verilog/coms.v(115[11:12])
    defparam i1_2_lut_4_lut_adj_1402.LUT_INIT = 16'hfe00;
    SB_LUT4 i1_2_lut_adj_1403 (.I0(\FRAME_MATCHER.i_31__N_2524 ), .I1(n74), 
            .I2(GND_net), .I3(GND_net), .O(n44092));
    defparam i1_2_lut_adj_1403.LUT_INIT = 16'hbbbb;
    SB_LUT4 equal_131_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4142));   // verilog/coms.v(154[7:23])
    defparam equal_131_i8_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 equal_122_i8_2_lut_3_lut (.I0(\FRAME_MATCHER.i [1]), .I1(\FRAME_MATCHER.i [2]), 
            .I2(\FRAME_MATCHER.i [0]), .I3(GND_net), .O(n8_adj_4147));   // verilog/coms.v(154[7:23])
    defparam equal_122_i8_2_lut_3_lut.LUT_INIT = 16'hdfdf;
    SB_LUT4 i15397_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44104), .I2(rx_data[7]), 
            .I3(\data_in_frame[3] [7]), .O(n28460));
    defparam i15397_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_4_lut_adj_1404 (.I0(n44255), .I1(\data_out_frame[14] [4]), 
            .I2(\data_out_frame[12] [2]), .I3(\data_out_frame[17] [1]), 
            .O(n44688));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_4_lut_adj_1404.LUT_INIT = 16'h6996;
    SB_LUT4 i15398_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44104), .I2(rx_data[6]), 
            .I3(\data_in_frame[3] [6]), .O(n28461));
    defparam i15398_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15399_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44104), .I2(rx_data[5]), 
            .I3(\data_in_frame[3] [5]), .O(n28462));
    defparam i15399_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1405 (.I0(\data_out_frame[19] [1]), .I1(n41589), 
            .I2(n42393), .I3(GND_net), .O(n27152));
    defparam i1_2_lut_3_lut_adj_1405.LUT_INIT = 16'h9696;
    SB_LUT4 i15400_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44104), .I2(rx_data[4]), 
            .I3(\data_in_frame[3] [4]), .O(n28463));
    defparam i15400_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1406 (.I0(\data_out_frame[19] [1]), .I1(n41589), 
            .I2(n41571), .I3(GND_net), .O(n2122));
    defparam i1_2_lut_3_lut_adj_1406.LUT_INIT = 16'h9696;
    SB_LUT4 i15401_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44104), .I2(rx_data[3]), 
            .I3(\data_in_frame[3] [3]), .O(n28464));
    defparam i15401_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15402_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44104), .I2(rx_data[2]), 
            .I3(\data_in_frame[3] [2]), .O(n28465));
    defparam i15402_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15403_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44104), .I2(rx_data[1]), 
            .I3(\data_in_frame[3] [1]), .O(n28466));
    defparam i15403_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15404_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44104), .I2(rx_data[0]), 
            .I3(\data_in_frame[3] [0]), .O(n28467));
    defparam i15404_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15389_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44104), .I2(rx_data[7]), 
            .I3(\data_in_frame[4] [7]), .O(n28452));
    defparam i15389_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1407 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[4] [1]), 
            .I2(\data_out_frame[6] [3]), .I3(GND_net), .O(n26712));   // verilog/coms.v(75[16:43])
    defparam i1_2_lut_3_lut_adj_1407.LUT_INIT = 16'h9696;
    SB_LUT4 i15390_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44104), .I2(rx_data[6]), 
            .I3(\data_in_frame[4] [6]), .O(n28453));
    defparam i15390_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i5_3_lut_4_lut_adj_1408 (.I0(\data_out_frame[6] [0]), .I1(\data_out_frame[8] [1]), 
            .I2(n10_adj_4128), .I3(\data_out_frame[5] [5]), .O(n1519));   // verilog/coms.v(72[16:27])
    defparam i5_3_lut_4_lut_adj_1408.LUT_INIT = 16'h6996;
    SB_LUT4 i15391_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44104), .I2(rx_data[5]), 
            .I3(\data_in_frame[4] [5]), .O(n28454));
    defparam i15391_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_2_lut (.I0(rx_data_ready), .I1(\FRAME_MATCHER.rx_data_ready_prev ), 
            .I2(GND_net), .I3(GND_net), .O(n161));   // verilog/coms.v(153[9:50])
    defparam i14_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15392_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44104), .I2(rx_data[4]), 
            .I3(\data_in_frame[4] [4]), .O(n28455));
    defparam i15392_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_427_Select_1_i3_2_lut (.I0(\FRAME_MATCHER.i [1]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4230));
    defparam select_427_Select_1_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1409 (.I0(\data_out_frame[12] [5]), .I1(\data_out_frame[12] [4]), 
            .I2(n1516), .I3(GND_net), .O(n44201));
    defparam i1_2_lut_3_lut_adj_1409.LUT_INIT = 16'h9696;
    SB_LUT4 i15393_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44104), .I2(rx_data[3]), 
            .I3(\data_in_frame[4] [3]), .O(n28456));
    defparam i15393_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_427_Select_2_i3_2_lut (.I0(\FRAME_MATCHER.i [2]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4228));
    defparam select_427_Select_2_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_3_i3_2_lut (.I0(\FRAME_MATCHER.i [3]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4226));
    defparam select_427_Select_3_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_4_i3_2_lut (.I0(\FRAME_MATCHER.i [4]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4224));
    defparam select_427_Select_4_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_5_i3_2_lut (.I0(\FRAME_MATCHER.i [5]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4223));
    defparam select_427_Select_5_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_6_i3_2_lut (.I0(\FRAME_MATCHER.i [6]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4222));
    defparam select_427_Select_6_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15394_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44104), .I2(rx_data[2]), 
            .I3(\data_in_frame[4] [2]), .O(n28457));
    defparam i15394_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_427_Select_7_i3_2_lut (.I0(\FRAME_MATCHER.i [7]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4221));
    defparam select_427_Select_7_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_2_lut_3_lut_adj_1410 (.I0(\data_out_frame[5] [3]), .I1(\data_out_frame[9] [4]), 
            .I2(\data_out_frame[9] [5]), .I3(GND_net), .O(n44258));
    defparam i1_2_lut_3_lut_adj_1410.LUT_INIT = 16'h9696;
    SB_LUT4 i15395_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44104), .I2(rx_data[1]), 
            .I3(\data_in_frame[4] [1]), .O(n28458));
    defparam i15395_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15396_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44104), .I2(rx_data[0]), 
            .I3(\data_in_frame[4] [0]), .O(n28459));
    defparam i15396_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15381_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44104), .I2(rx_data[7]), 
            .I3(\data_in_frame[5] [7]), .O(n28444));
    defparam i15381_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1411 (.I0(n33565), .I1(\FRAME_MATCHER.i [5]), .I2(\FRAME_MATCHER.i [4]), 
            .I3(\FRAME_MATCHER.i [3]), .O(n44085));   // verilog/coms.v(154[7:23])
    defparam i3_4_lut_adj_1411.LUT_INIT = 16'hffdf;
    SB_LUT4 i15382_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44104), .I2(rx_data[6]), 
            .I3(\data_in_frame[5] [6]), .O(n28445));
    defparam i15382_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_427_Select_8_i3_2_lut (.I0(\FRAME_MATCHER.i [8]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4220));
    defparam select_427_Select_8_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_9_i3_2_lut (.I0(\FRAME_MATCHER.i [9]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4219));
    defparam select_427_Select_9_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_10_i3_2_lut (.I0(\FRAME_MATCHER.i [10]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4218));
    defparam select_427_Select_10_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_11_i3_2_lut (.I0(\FRAME_MATCHER.i [11]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4217));
    defparam select_427_Select_11_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_12_i3_2_lut (.I0(\FRAME_MATCHER.i [12]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4216));
    defparam select_427_Select_12_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15383_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44104), .I2(rx_data[5]), 
            .I3(\data_in_frame[5] [5]), .O(n28446));
    defparam i15383_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_427_Select_13_i3_2_lut (.I0(\FRAME_MATCHER.i [13]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4215));
    defparam select_427_Select_13_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15384_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44104), .I2(rx_data[4]), 
            .I3(\data_in_frame[5] [4]), .O(n28447));
    defparam i15384_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_3_lut_adj_1412 (.I0(\data_out_frame[4] [2]), .I1(\data_out_frame[6] [4]), 
            .I2(\data_out_frame[4] [3]), .I3(GND_net), .O(n27407));
    defparam i1_2_lut_3_lut_adj_1412.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1413 (.I0(\data_out_frame[5] [5]), .I1(\data_out_frame[5] [4]), 
            .I2(n44573), .I3(\data_out_frame[5] [3]), .O(n1168));   // verilog/coms.v(71[16:62])
    defparam i2_3_lut_4_lut_adj_1413.LUT_INIT = 16'h6996;
    SB_LUT4 select_427_Select_14_i3_2_lut (.I0(\FRAME_MATCHER.i [14]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4214));
    defparam select_427_Select_14_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i2_3_lut_4_lut_adj_1414 (.I0(\data_out_frame[4] [6]), .I1(\data_out_frame[5] [0]), 
            .I2(n1168), .I3(\data_out_frame[7] [0]), .O(n27666));   // verilog/coms.v(85[17:70])
    defparam i2_3_lut_4_lut_adj_1414.LUT_INIT = 16'h6996;
    SB_LUT4 select_427_Select_15_i3_2_lut (.I0(\FRAME_MATCHER.i [15]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4213));
    defparam select_427_Select_15_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15385_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44104), .I2(rx_data[3]), 
            .I3(\data_in_frame[5] [3]), .O(n28448));
    defparam i15385_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_427_Select_16_i3_2_lut (.I0(\FRAME_MATCHER.i [16]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4212));
    defparam select_427_Select_16_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_17_i3_2_lut (.I0(\FRAME_MATCHER.i [17]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4211));
    defparam select_427_Select_17_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_18_i3_2_lut (.I0(\FRAME_MATCHER.i [18]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4210));
    defparam select_427_Select_18_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_19_i3_2_lut (.I0(\FRAME_MATCHER.i [19]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4209));
    defparam select_427_Select_19_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_20_i3_2_lut (.I0(\FRAME_MATCHER.i [20]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4208));
    defparam select_427_Select_20_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_21_i3_2_lut (.I0(\FRAME_MATCHER.i [21]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4207));
    defparam select_427_Select_21_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_22_i3_2_lut (.I0(\FRAME_MATCHER.i [22]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4206));
    defparam select_427_Select_22_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_23_i3_2_lut (.I0(\FRAME_MATCHER.i [23]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4205));
    defparam select_427_Select_23_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15386_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44104), .I2(rx_data[2]), 
            .I3(\data_in_frame[5] [2]), .O(n28449));
    defparam i15386_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15269_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44085), .I2(rx_data[7]), 
            .I3(\data_in_frame[19] [7]), .O(n28332));
    defparam i15269_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_427_Select_24_i3_2_lut (.I0(\FRAME_MATCHER.i [24]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4204));
    defparam select_427_Select_24_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_25_i3_2_lut (.I0(\FRAME_MATCHER.i [25]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4203));
    defparam select_427_Select_25_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_26_i3_2_lut (.I0(\FRAME_MATCHER.i [26]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4202));
    defparam select_427_Select_26_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_27_i3_2_lut (.I0(\FRAME_MATCHER.i [27]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4201));
    defparam select_427_Select_27_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15387_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44104), .I2(rx_data[1]), 
            .I3(\data_in_frame[5] [1]), .O(n28450));
    defparam i15387_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 select_427_Select_28_i3_2_lut (.I0(\FRAME_MATCHER.i [28]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4200));
    defparam select_427_Select_28_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_29_i3_2_lut (.I0(\FRAME_MATCHER.i [29]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4199));
    defparam select_427_Select_29_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_30_i3_2_lut (.I0(\FRAME_MATCHER.i [30]), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4198));
    defparam select_427_Select_30_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 select_427_Select_31_i3_2_lut (.I0(\FRAME_MATCHER.i[31] ), .I1(n26472), 
            .I2(GND_net), .I3(GND_net), .O(n3_adj_4197));
    defparam select_427_Select_31_i3_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i15388_3_lut_4_lut (.I0(n8_adj_4177), .I1(n44104), .I2(rx_data[0]), 
            .I3(\data_in_frame[5] [0]), .O(n28451));
    defparam i15388_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15373_3_lut_4_lut (.I0(n8_adj_4232), .I1(n44104), .I2(rx_data[7]), 
            .I3(\data_in_frame[6] [7]), .O(n28436));
    defparam i15373_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15374_3_lut_4_lut (.I0(n8_adj_4232), .I1(n44104), .I2(rx_data[6]), 
            .I3(\data_in_frame[6] [6]), .O(n28437));
    defparam i15374_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15270_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44085), .I2(rx_data[6]), 
            .I3(\data_in_frame[19] [6]), .O(n28333));
    defparam i15270_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15375_3_lut_4_lut (.I0(n8_adj_4232), .I1(n44104), .I2(rx_data[5]), 
            .I3(\data_in_frame[6] [5]), .O(n28438));
    defparam i15375_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15376_3_lut_4_lut (.I0(n8_adj_4232), .I1(n44104), .I2(rx_data[4]), 
            .I3(\data_in_frame[6] [4]), .O(n28439));
    defparam i15376_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1415 (.I0(\data_out_frame[25] [6]), .I1(n44486), 
            .I2(n42339), .I3(n41597), .O(n46095));
    defparam i3_4_lut_adj_1415.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1416 (.I0(\data_out_frame[25] [7]), .I1(n42333), 
            .I2(\data_out_frame[23] [6]), .I3(GND_net), .O(n44486));
    defparam i2_3_lut_adj_1416.LUT_INIT = 16'h6969;
    SB_LUT4 i5_4_lut_adj_1417 (.I0(n44494), .I1(n44531), .I2(n41846), 
            .I3(n44486), .O(n12_adj_4302));
    defparam i5_4_lut_adj_1417.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1418 (.I0(n42407), .I1(n12_adj_4302), .I2(n44540), 
            .I3(n44381), .O(n45401));
    defparam i6_4_lut_adj_1418.LUT_INIT = 16'h6996;
    SB_LUT4 i4_2_lut_adj_1419 (.I0(\data_out_frame[24] [0]), .I1(n42393), 
            .I2(GND_net), .I3(GND_net), .O(n12_adj_4303));   // verilog/coms.v(71[16:27])
    defparam i4_2_lut_adj_1419.LUT_INIT = 16'h9999;
    SB_LUT4 i5_4_lut_adj_1420 (.I0(\data_out_frame[24] [1]), .I1(n44237), 
            .I2(n27497), .I3(\data_out_frame[23] [6]), .O(n13));   // verilog/coms.v(71[16:27])
    defparam i5_4_lut_adj_1420.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1421 (.I0(n13), .I1(n44436), .I2(n12_adj_4303), 
            .I3(n44687), .O(n45555));   // verilog/coms.v(71[16:27])
    defparam i7_4_lut_adj_1421.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1422 (.I0(n44683), .I1(n44685), .I2(GND_net), 
            .I3(GND_net), .O(n44687));
    defparam i1_2_lut_adj_1422.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1423 (.I0(\data_out_frame[10] [1]), .I1(\data_out_frame[7] [7]), 
            .I2(\data_out_frame[7] [6]), .I3(\data_out_frame[8] [0]), .O(n6_adj_4123));   // verilog/coms.v(74[16:27])
    defparam i1_2_lut_4_lut_adj_1423.LUT_INIT = 16'h6996;
    SB_LUT4 i15377_3_lut_4_lut (.I0(n8_adj_4232), .I1(n44104), .I2(rx_data[3]), 
            .I3(\data_in_frame[6] [3]), .O(n28440));
    defparam i15377_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1424 (.I0(\data_out_frame[23] [7]), .I1(n44381), 
            .I2(n42407), .I3(n42333), .O(n45867));
    defparam i3_4_lut_adj_1424.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1425 (.I0(n42378), .I1(n27497), .I2(GND_net), 
            .I3(GND_net), .O(n42487));
    defparam i1_2_lut_adj_1425.LUT_INIT = 16'h6666;
    SB_LUT4 i15378_3_lut_4_lut (.I0(n8_adj_4232), .I1(n44104), .I2(rx_data[2]), 
            .I3(\data_in_frame[6] [2]), .O(n28441));
    defparam i15378_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1426 (.I0(n41521), .I1(\data_out_frame[19] [4]), 
            .I2(n42487), .I3(n42407), .O(n41437));
    defparam i3_4_lut_adj_1426.LUT_INIT = 16'h9669;
    SB_LUT4 i2_3_lut_adj_1427 (.I0(\data_out_frame[24] [2]), .I1(n44390), 
            .I2(n41437), .I3(GND_net), .O(n46700));
    defparam i2_3_lut_adj_1427.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_4_lut_adj_1428 (.I0(\data_out_frame[7] [5]), .I1(\data_out_frame[7] [4]), 
            .I2(\data_out_frame[5] [2]), .I3(\data_out_frame[10] [0]), .O(n44285));   // verilog/coms.v(74[16:27])
    defparam i2_3_lut_4_lut_adj_1428.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1429 (.I0(\data_out_frame[24] [3]), .I1(n42363), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4304));
    defparam i1_2_lut_adj_1429.LUT_INIT = 16'h9999;
    SB_LUT4 i4_4_lut_adj_1430 (.I0(\data_out_frame[20] [5]), .I1(n42407), 
            .I2(n44683), .I3(n6_adj_4304), .O(n44390));
    defparam i4_4_lut_adj_1430.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1431 (.I0(n1794), .I1(n27321), .I2(\data_out_frame[18] [7]), 
            .I3(\data_out_frame[16] [5]), .O(n6_adj_4121));
    defparam i1_2_lut_4_lut_adj_1431.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1432 (.I0(\data_out_frame[17] [6]), .I1(\data_out_frame[19] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n44237));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1432.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1433 (.I0(\data_out_frame[20] [0]), .I1(\data_out_frame[19] [7]), 
            .I2(n44240), .I3(n6_adj_4245), .O(n42407));
    defparam i4_4_lut_adj_1433.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_4_lut_adj_1434 (.I0(\data_out_frame[12] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(n44727), .I3(\data_out_frame[11] [6]), .O(n44576));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_4_lut_adj_1434.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_3_lut_adj_1435 (.I0(\data_out_frame[5] [1]), .I1(n44727), 
            .I2(\data_out_frame[11] [6]), .I3(GND_net), .O(n44597));
    defparam i1_2_lut_3_lut_adj_1435.LUT_INIT = 16'h9696;
    SB_LUT4 i15379_3_lut_4_lut (.I0(n8_adj_4232), .I1(n44104), .I2(rx_data[1]), 
            .I3(\data_in_frame[6] [1]), .O(n28442));
    defparam i15379_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1436 (.I0(\data_out_frame[24] [5]), .I1(n42350), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4305));
    defparam i1_2_lut_adj_1436.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1437 (.I0(n42444), .I1(n41565), .I2(\data_out_frame[24] [6]), 
            .I3(n6_adj_4305), .O(n45769));
    defparam i4_4_lut_adj_1437.LUT_INIT = 16'h6996;
    SB_LUT4 i15380_3_lut_4_lut (.I0(n8_adj_4232), .I1(n44104), .I2(rx_data[0]), 
            .I3(\data_in_frame[6] [0]), .O(n28443));
    defparam i15380_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1438 (.I0(n45752), .I1(n27163), .I2(GND_net), 
            .I3(GND_net), .O(n41565));
    defparam i1_2_lut_adj_1438.LUT_INIT = 16'h9999;
    SB_LUT4 i1_2_lut_4_lut_adj_1439 (.I0(\data_out_frame[20] [7]), .I1(n41486), 
            .I2(n41571), .I3(\data_out_frame[16] [5]), .O(n6_adj_4118));
    defparam i1_2_lut_4_lut_adj_1439.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1440 (.I0(\data_out_frame[7] [1]), .I1(n1168), 
            .I2(\data_out_frame[4] [7]), .I3(\data_out_frame[9] [3]), .O(n44612));
    defparam i1_2_lut_4_lut_adj_1440.LUT_INIT = 16'h6996;
    SB_LUT4 i4_4_lut_adj_1441 (.I0(n44662), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[19] [7]), .I3(n44748), .O(n10_adj_4243));
    defparam i4_4_lut_adj_1441.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1442 (.I0(\data_out_frame[19] [7]), .I1(\data_out_frame[19] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n26881));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_adj_1442.LUT_INIT = 16'h6666;
    SB_LUT4 i7_4_lut_adj_1443 (.I0(\data_out_frame[8] [3]), .I1(n27687), 
            .I2(n27212), .I3(\data_out_frame[13] [1]), .O(n18_adj_4306));
    defparam i7_4_lut_adj_1443.LUT_INIT = 16'h6996;
    SB_LUT4 i5_2_lut_adj_1444 (.I0(\data_out_frame[11] [0]), .I1(n42387), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4307));
    defparam i5_2_lut_adj_1444.LUT_INIT = 16'h6666;
    SB_LUT4 i15271_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44085), .I2(rx_data[5]), 
            .I3(\data_in_frame[19] [5]), .O(n28334));
    defparam i15271_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15272_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44085), .I2(rx_data[4]), 
            .I3(\data_in_frame[19] [4]), .O(n28335));
    defparam i15272_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i9_4_lut_adj_1445 (.I0(\data_out_frame[12] [7]), .I1(n18_adj_4306), 
            .I2(n42387), .I3(n44570), .O(n20_adj_4308));
    defparam i9_4_lut_adj_1445.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_1446 (.I0(n44342), .I1(n20_adj_4308), .I2(n16_adj_4307), 
            .I3(\data_out_frame[8] [4]), .O(n41525));
    defparam i10_4_lut_adj_1446.LUT_INIT = 16'h6996;
    SB_LUT4 i3_4_lut_adj_1447 (.I0(n41525), .I1(n44421), .I2(n41480), 
            .I3(\data_out_frame[15] [1]), .O(n27497));
    defparam i3_4_lut_adj_1447.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_adj_1448 (.I0(n42365), .I1(n27244), .I2(\data_out_frame[17] [4]), 
            .I3(GND_net), .O(n44506));
    defparam i2_3_lut_adj_1448.LUT_INIT = 16'h9696;
    SB_LUT4 i2_3_lut_adj_1449 (.I0(n27546), .I1(n44506), .I2(n27497), 
            .I3(GND_net), .O(n46294));
    defparam i2_3_lut_adj_1449.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1450 (.I0(\data_out_frame[15] [2]), .I1(\data_out_frame[17] [3]), 
            .I2(GND_net), .I3(GND_net), .O(n44421));
    defparam i1_2_lut_adj_1450.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1451 (.I0(\data_out_frame[19] [3]), .I1(\data_out_frame[19] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n44480));
    defparam i1_2_lut_adj_1451.LUT_INIT = 16'h6666;
    SB_LUT4 i15273_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44085), .I2(rx_data[3]), 
            .I3(\data_in_frame[19] [3]), .O(n28336));
    defparam i15273_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1452 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[17] [5]), 
            .I2(GND_net), .I3(GND_net), .O(n44433));
    defparam i1_2_lut_adj_1452.LUT_INIT = 16'h6666;
    SB_LUT4 i11_4_lut_adj_1453 (.I0(n44688), .I1(\data_out_frame[18] [3]), 
            .I2(\data_out_frame[16] [1]), .I3(n44433), .O(n30_adj_4309));
    defparam i11_4_lut_adj_1453.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1454 (.I0(\data_out_frame[17] [4]), .I1(n30_adj_4309), 
            .I2(\data_out_frame[17] [2]), .I3(n44409), .O(n34_adj_4310));
    defparam i15_4_lut_adj_1454.LUT_INIT = 16'h6996;
    SB_LUT4 i13_4_lut_adj_1455 (.I0(n44480), .I1(n44395), .I2(n44421), 
            .I3(n44195), .O(n32));
    defparam i13_4_lut_adj_1455.LUT_INIT = 16'h6996;
    SB_LUT4 i15274_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44085), .I2(rx_data[2]), 
            .I3(\data_in_frame[19] [2]), .O(n28337));
    defparam i15274_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15275_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44085), .I2(rx_data[1]), 
            .I3(\data_in_frame[19] [1]), .O(n28338));
    defparam i15275_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i15276_3_lut_4_lut (.I0(n8_adj_4147), .I1(n44085), .I2(rx_data[0]), 
            .I3(\data_in_frame[19] [0]), .O(n28339));
    defparam i15276_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_4_lut_adj_1456 (.I0(n26881), .I1(\data_out_frame[19] [2]), 
            .I2(\data_out_frame[19] [6]), .I3(\data_out_frame[16] [3]), 
            .O(n33));
    defparam i14_4_lut_adj_1456.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1457 (.I0(n44333), .I1(\data_out_frame[16] [0]), 
            .I2(\data_out_frame[18] [6]), .I3(\data_out_frame[19] [1]), 
            .O(n31_adj_4311));
    defparam i12_4_lut_adj_1457.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1458 (.I0(n31_adj_4311), .I1(n33), .I2(n32), 
            .I3(n34_adj_4310), .O(n45838));
    defparam i18_4_lut_adj_1458.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1459 (.I0(n41589), .I1(n41571), .I2(n44518), 
            .I3(n41521), .O(n16_adj_4312));
    defparam i6_4_lut_adj_1459.LUT_INIT = 16'h6996;
    SB_LUT4 i2_3_lut_4_lut_adj_1460 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[11] [4]), 
            .I2(n24830), .I3(n26380), .O(n27110));
    defparam i2_3_lut_4_lut_adj_1460.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_0__bdd_4_lut_36479 (.I0(\byte_transmit_counter[0] ), 
            .I1(\data_out_frame[18][0] ), .I2(\data_out_frame[19] [0]), 
            .I3(byte_transmit_counter[1]), .O(n51429));
    defparam byte_transmit_counter_0__bdd_4_lut_36479.LUT_INIT = 16'he4aa;
    SB_LUT4 n51429_bdd_4_lut (.I0(n51429), .I1(\data_out_frame[17] [0]), 
            .I2(\data_out_frame[16] [0]), .I3(byte_transmit_counter[1]), 
            .O(n51432));
    defparam n51429_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i7_4_lut_adj_1461 (.I0(\data_out_frame[23] [3]), .I1(n45838), 
            .I2(n44534), .I3(n41571), .O(n17_adj_4313));
    defparam i7_4_lut_adj_1461.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1462 (.I0(n17_adj_4313), .I1(n42363), .I2(n16_adj_4312), 
            .I3(n26846), .O(n44494));
    defparam i9_4_lut_adj_1462.LUT_INIT = 16'h9669;
    SB_LUT4 i5_3_lut_4_lut_adj_1463 (.I0(\data_out_frame[11] [5]), .I1(\data_out_frame[11] [4]), 
            .I2(n44524), .I3(n27687), .O(n14_adj_4117));
    defparam i5_3_lut_4_lut_adj_1463.LUT_INIT = 16'h6996;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_36508 (.I0(byte_transmit_counter[1]), 
            .I1(n49818), .I2(n49819), .I3(\byte_transmit_counter[2] ), 
            .O(n51423));
    defparam byte_transmit_counter_1__bdd_4_lut_36508.LUT_INIT = 16'he4aa;
    SB_LUT4 n51423_bdd_4_lut (.I0(n51423), .I1(n17_adj_4314), .I2(n15), 
            .I3(\byte_transmit_counter[2] ), .O(n51426));
    defparam n51423_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_36470 (.I0(byte_transmit_counter[1]), 
            .I1(n49803), .I2(n49804), .I3(\byte_transmit_counter[2] ), 
            .O(n51417));
    defparam byte_transmit_counter_1__bdd_4_lut_36470.LUT_INIT = 16'he4aa;
    SB_LUT4 n51417_bdd_4_lut (.I0(n51417), .I1(n17_adj_4316), .I2(n16_adj_4317), 
            .I3(\byte_transmit_counter[2] ), .O(n51420));
    defparam n51417_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 byte_transmit_counter_1__bdd_4_lut_36465 (.I0(byte_transmit_counter[1]), 
            .I1(n49806), .I2(n49807), .I3(\byte_transmit_counter[2] ), 
            .O(n51411));
    defparam byte_transmit_counter_1__bdd_4_lut_36465.LUT_INIT = 16'he4aa;
    SB_LUT4 n51411_bdd_4_lut (.I0(n51411), .I1(n17_adj_4318), .I2(n16_adj_4319), 
            .I3(\byte_transmit_counter[2] ), .O(n51414));
    defparam n51411_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i5_4_lut_adj_1464 (.I0(n44685), .I1(n44436), .I2(n41525), 
            .I3(\data_out_frame[17] [5]), .O(n13_adj_4320));
    defparam i5_4_lut_adj_1464.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1465 (.I0(n13_adj_4320), .I1(n11_adj_4281), .I2(n46294), 
            .I3(n44451), .O(n46491));
    defparam i7_4_lut_adj_1465.LUT_INIT = 16'h9669;
    SB_LUT4 i15261_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44085), .I2(rx_data[7]), 
            .I3(\data_in_frame[20] [7]), .O(n28324));
    defparam i15261_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i16_3_lut (.I0(\data_out_frame[16] [4]), 
            .I1(\data_out_frame[17] [4]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n16_adj_4319));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_4_i17_3_lut (.I0(\data_out_frame[18] [4]), 
            .I1(\data_out_frame[19] [4]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n17_adj_4318));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_4_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34999_2_lut (.I0(\data_out_frame[23] [4]), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n49807));
    defparam i34999_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35046_2_lut (.I0(\data_out_frame[20] [4]), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n49806));
    defparam i35046_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i16_3_lut (.I0(\data_out_frame[16] [5]), 
            .I1(\data_out_frame[17] [5]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n16_adj_4317));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i16_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1466 (.I0(\data_out_frame[24] [5]), .I1(\data_out_frame[24] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27178));
    defparam i1_2_lut_adj_1466.LUT_INIT = 16'h6666;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_5_i17_3_lut (.I0(\data_out_frame[18] [5]), 
            .I1(\data_out_frame[19] [5]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n17_adj_4316));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_5_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35047_2_lut (.I0(\data_out_frame[23] [5]), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n49804));
    defparam i35047_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i35049_2_lut (.I0(\data_out_frame[20] [5]), .I1(\byte_transmit_counter[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n49803));
    defparam i35049_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 byte_transmit_counter_4__I_0_Mux_6_i17_3_lut (.I0(\data_out_frame[18] [6]), 
            .I1(\data_out_frame[19] [6]), .I2(\byte_transmit_counter[0] ), 
            .I3(GND_net), .O(n17_adj_4314));   // verilog/coms.v(106[34:55])
    defparam byte_transmit_counter_4__I_0_Mux_6_i17_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_adj_1467 (.I0(\data_out_frame[24] [6]), .I1(\data_out_frame[24] [7]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4321));
    defparam i1_2_lut_adj_1467.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1468 (.I0(\data_out_frame[24] [3]), .I1(n42350), 
            .I2(n27178), .I3(n6_adj_4321), .O(n44540));
    defparam i4_4_lut_adj_1468.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1469 (.I0(\data_out_frame[20] [3]), .I1(n42361), 
            .I2(GND_net), .I3(GND_net), .O(n42448));
    defparam i1_2_lut_adj_1469.LUT_INIT = 16'h9999;
    SB_LUT4 i11_4_lut_adj_1470 (.I0(\data_out_frame[23] [6]), .I1(\data_out_frame[23] [5]), 
            .I2(n44540), .I3(n42339), .O(n26_adj_4322));
    defparam i11_4_lut_adj_1470.LUT_INIT = 16'h6996;
    SB_LUT4 i9_4_lut_adj_1471 (.I0(n44694), .I1(n42448), .I2(n27152), 
            .I3(\data_out_frame[20] [5]), .O(n24_adj_4323));
    defparam i9_4_lut_adj_1471.LUT_INIT = 16'h9669;
    SB_LUT4 i10_4_lut_adj_1472 (.I0(n46491), .I1(n44494), .I2(\data_out_frame[23] [7]), 
            .I3(n26249), .O(n25_adj_4324));
    defparam i10_4_lut_adj_1472.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_4_lut_adj_1473 (.I0(n42312), .I1(n2122), .I2(\data_out_frame[23] [3]), 
            .I3(n44534), .O(n42434));
    defparam i1_2_lut_4_lut_adj_1473.LUT_INIT = 16'h6996;
    SB_LUT4 i14_4_lut_adj_1474 (.I0(n23), .I1(n25_adj_4324), .I2(n24_adj_4323), 
            .I3(n26_adj_4322), .O(n41846));
    defparam i14_4_lut_adj_1474.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_adj_1475 (.I0(n44427), .I1(\data_out_frame[25] [1]), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_4325));
    defparam i2_2_lut_adj_1475.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1476 (.I0(n44489), .I1(\data_out_frame[25] [4]), 
            .I2(\data_out_frame[25] [7]), .I3(n41846), .O(n14_adj_4326));
    defparam i6_4_lut_adj_1476.LUT_INIT = 16'h9669;
    SB_LUT4 i7_4_lut_adj_1477 (.I0(n42434), .I1(n14_adj_4326), .I2(n10_adj_4325), 
            .I3(n42339), .O(n27163));
    defparam i7_4_lut_adj_1477.LUT_INIT = 16'h6996;
    SB_LUT4 i15262_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44085), .I2(rx_data[6]), 
            .I3(\data_in_frame[20] [6]), .O(n28325));
    defparam i15262_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1478 (.I0(n46282), .I1(n27163), .I2(GND_net), 
            .I3(GND_net), .O(n42381));
    defparam i1_2_lut_adj_1478.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_adj_1479 (.I0(\data_out_frame[17] [7]), .I1(\data_out_frame[18][0] ), 
            .I2(GND_net), .I3(GND_net), .O(n44748));
    defparam i1_2_lut_adj_1479.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1480 (.I0(\data_out_frame[15] [7]), .I1(\data_out_frame[15] [6]), 
            .I2(\data_out_frame[16] [0]), .I3(GND_net), .O(n27561));   // verilog/coms.v(71[16:27])
    defparam i1_2_lut_3_lut_adj_1480.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1481 (.I0(n44579), .I1(n44621), .I2(\data_out_frame[6] [6]), 
            .I3(n44221), .O(n15_adj_4327));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_1481.LUT_INIT = 16'h6996;
    SB_LUT4 i8_4_lut_adj_1482 (.I0(n15_adj_4327), .I1(\data_out_frame[10] [6]), 
            .I2(n14_adj_4241), .I3(\data_out_frame[4] [0]), .O(n27546));   // verilog/coms.v(74[16:43])
    defparam i8_4_lut_adj_1482.LUT_INIT = 16'h6996;
    SB_LUT4 i5_4_lut_adj_1483 (.I0(\data_out_frame[15] [6]), .I1(n44195), 
            .I2(n46733), .I3(n27546), .O(n12_adj_4328));   // verilog/coms.v(74[16:43])
    defparam i5_4_lut_adj_1483.LUT_INIT = 16'h9669;
    SB_LUT4 i6_4_lut_adj_1484 (.I0(n26226), .I1(n12_adj_4328), .I2(n44564), 
            .I3(n42344), .O(n26249));   // verilog/coms.v(74[16:43])
    defparam i6_4_lut_adj_1484.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1485 (.I0(\data_out_frame[20] [2]), .I1(n26249), 
            .I2(GND_net), .I3(GND_net), .O(n44129));
    defparam i1_2_lut_adj_1485.LUT_INIT = 16'h6666;
    SB_LUT4 i5_4_lut_adj_1486 (.I0(n42438), .I1(n42427), .I2(\data_out_frame[25] [0]), 
            .I3(n45876), .O(n12_adj_4329));
    defparam i5_4_lut_adj_1486.LUT_INIT = 16'h6996;
    SB_LUT4 i6_4_lut_adj_1487 (.I0(n46282), .I1(n12_adj_4329), .I2(\data_out_frame[24] [6]), 
            .I3(n46253), .O(n45752));
    defparam i6_4_lut_adj_1487.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1488 (.I0(\data_out_frame[25] [1]), .I1(n45752), 
            .I2(GND_net), .I3(GND_net), .O(n42395));
    defparam i1_2_lut_adj_1488.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_4_lut_adj_1489 (.I0(\data_out_frame[16] [2]), .I1(\data_out_frame[20] [5]), 
            .I2(\data_out_frame[20] [6]), .I3(n42312), .O(n9));
    defparam i2_3_lut_4_lut_adj_1489.LUT_INIT = 16'h6996;
    SB_LUT4 i2_2_lut_3_lut_adj_1490 (.I0(\data_out_frame[9] [1]), .I1(\data_out_frame[5] [1]), 
            .I2(n44727), .I3(GND_net), .O(n10_adj_4113));
    defparam i2_2_lut_3_lut_adj_1490.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_3_lut_adj_1491 (.I0(\data_out_frame[4] [3]), .I1(\data_out_frame[6] [5]), 
            .I2(\data_out_frame[4] [4]), .I3(GND_net), .O(n27212));
    defparam i1_2_lut_3_lut_adj_1491.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1492 (.I0(\data_out_frame[15] [3]), .I1(\data_out_frame[15] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n27244));
    defparam i1_2_lut_adj_1492.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_4_lut_adj_1493 (.I0(\data_out_frame[18][2] ), .I1(\data_out_frame[16] [4]), 
            .I2(\data_out_frame[18] [5]), .I3(n44318), .O(n44333));
    defparam i1_2_lut_4_lut_adj_1493.LUT_INIT = 16'h6996;
    SB_LUT4 i1_2_lut_adj_1494 (.I0(n41601), .I1(\data_out_frame[13] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n42344));
    defparam i1_2_lut_adj_1494.LUT_INIT = 16'h6666;
    SB_LUT4 i1_2_lut_3_lut_adj_1495 (.I0(\data_out_frame[4] [4]), .I1(\data_out_frame[9] [0]), 
            .I2(\data_out_frame[4] [5]), .I3(GND_net), .O(n27539));   // verilog/coms.v(76[16:27])
    defparam i1_2_lut_3_lut_adj_1495.LUT_INIT = 16'h9696;
    SB_LUT4 i6_4_lut_adj_1496 (.I0(\data_out_frame[11] [1]), .I1(\data_out_frame[11] [2]), 
            .I2(n44570), .I3(n27666), .O(n14_adj_4330));   // verilog/coms.v(85[17:28])
    defparam i6_4_lut_adj_1496.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1497 (.I0(\data_out_frame[15] [4]), .I1(n14_adj_4330), 
            .I2(n10_adj_4240), .I3(n44712), .O(n44564));   // verilog/coms.v(85[17:28])
    defparam i7_4_lut_adj_1497.LUT_INIT = 16'h6996;
    SB_LUT4 i15263_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44085), .I2(rx_data[5]), 
            .I3(\data_in_frame[20] [5]), .O(n28326));
    defparam i15263_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i1_2_lut_adj_1498 (.I0(\data_out_frame[15] [3]), .I1(n44564), 
            .I2(GND_net), .I3(GND_net), .O(n44451));
    defparam i1_2_lut_adj_1498.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut_adj_1499 (.I0(\data_out_frame[10] [7]), .I1(\data_out_frame[13] [3]), 
            .I2(\data_out_frame[8] [7]), .I3(GND_net), .O(n44210));   // verilog/coms.v(85[17:28])
    defparam i2_3_lut_adj_1499.LUT_INIT = 16'h9696;
    SB_LUT4 i1_2_lut_adj_1500 (.I0(\data_out_frame[8] [5]), .I1(\data_out_frame[13] [2]), 
            .I2(GND_net), .I3(GND_net), .O(n44221));   // verilog/coms.v(74[16:43])
    defparam i1_2_lut_adj_1500.LUT_INIT = 16'h6666;
    SB_LUT4 i19_4_lut_adj_1501 (.I0(n44218), .I1(n42075), .I2(\data_out_frame[6] [5]), 
            .I3(\data_out_frame[11] [3]), .O(n46));
    defparam i19_4_lut_adj_1501.LUT_INIT = 16'h6996;
    SB_LUT4 i17_4_lut_adj_1502 (.I0(\data_out_frame[6] [4]), .I1(\data_out_frame[13] [0]), 
            .I2(\data_out_frame[14] [5]), .I3(\data_out_frame[14] [6]), 
            .O(n44_adj_4331));
    defparam i17_4_lut_adj_1502.LUT_INIT = 16'h6996;
    SB_LUT4 i18_4_lut_adj_1503 (.I0(n44700), .I1(n44461), .I2(n44576), 
            .I3(n44304), .O(n45_adj_4332));
    defparam i18_4_lut_adj_1503.LUT_INIT = 16'h6996;
    SB_LUT4 i16_4_lut_adj_1504 (.I0(n27558), .I1(n44543), .I2(\data_out_frame[14] [7]), 
            .I3(n44221), .O(n43_adj_4333));
    defparam i16_4_lut_adj_1504.LUT_INIT = 16'h6996;
    SB_LUT4 i15_4_lut_adj_1505 (.I0(\data_out_frame[14] [3]), .I1(n44612), 
            .I2(\data_out_frame[14] [0]), .I3(n44210), .O(n42_adj_4334));
    defparam i15_4_lut_adj_1505.LUT_INIT = 16'h6996;
    SB_LUT4 i15264_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44085), .I2(rx_data[4]), 
            .I3(\data_in_frame[20] [4]), .O(n28327));
    defparam i15264_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i14_4_lut_adj_1506 (.I0(n27110), .I1(n44366), .I2(n1699), 
            .I3(n44424), .O(n41_adj_4335));
    defparam i14_4_lut_adj_1506.LUT_INIT = 16'h9669;
    SB_LUT4 i25_4_lut_adj_1507 (.I0(n43_adj_4333), .I1(n45_adj_4332), .I2(n44_adj_4331), 
            .I3(n46), .O(n52));
    defparam i25_4_lut_adj_1507.LUT_INIT = 16'h6996;
    SB_LUT4 i20_4_lut_adj_1508 (.I0(\data_out_frame[13] [1]), .I1(\data_out_frame[14] [4]), 
            .I2(n42285), .I3(\data_out_frame[13] [4]), .O(n47));
    defparam i20_4_lut_adj_1508.LUT_INIT = 16'h9669;
    SB_LUT4 i26_4_lut (.I0(n47), .I1(n52), .I2(n41_adj_4335), .I3(n42_adj_4334), 
            .O(n41478));
    defparam i26_4_lut.LUT_INIT = 16'h6996;
    SB_LUT4 i3_2_lut_adj_1509 (.I0(\data_out_frame[15] [2]), .I1(n41478), 
            .I2(GND_net), .I3(GND_net), .O(n16_adj_4336));
    defparam i3_2_lut_adj_1509.LUT_INIT = 16'h6666;
    SB_LUT4 i9_4_lut_adj_1510 (.I0(n44451), .I1(n26226), .I2(n1699), .I3(n41486), 
            .O(n22_adj_4337));
    defparam i9_4_lut_adj_1510.LUT_INIT = 16'h6996;
    SB_LUT4 i7_3_lut (.I0(n42344), .I1(n50676), .I2(n27561), .I3(GND_net), 
            .O(n20_adj_4338));
    defparam i7_3_lut.LUT_INIT = 16'h9696;
    SB_LUT4 i11_4_lut_adj_1511 (.I0(n41540), .I1(n22_adj_4337), .I2(n16_adj_4336), 
            .I3(n44366), .O(n24_adj_4339));
    defparam i11_4_lut_adj_1511.LUT_INIT = 16'h6996;
    SB_LUT4 i15265_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44085), .I2(rx_data[3]), 
            .I3(\data_in_frame[20] [3]), .O(n28328));
    defparam i15265_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1512 (.I0(\data_out_frame[17] [7]), .I1(n44395), 
            .I2(n27220), .I3(n27244), .O(n45357));
    defparam i3_4_lut_adj_1512.LUT_INIT = 16'h6996;
    SB_LUT4 i12_4_lut_adj_1513 (.I0(n45357), .I1(n24_adj_4339), .I2(n20_adj_4338), 
            .I3(n1794), .O(n46733));
    defparam i12_4_lut_adj_1513.LUT_INIT = 16'h9669;
    SB_LUT4 i1_2_lut_adj_1514 (.I0(\data_out_frame[20] [3]), .I1(\data_out_frame[20] [4]), 
            .I2(GND_net), .I3(GND_net), .O(n27138));
    defparam i1_2_lut_adj_1514.LUT_INIT = 16'h6666;
    SB_LUT4 i15266_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44085), .I2(rx_data[2]), 
            .I3(\data_in_frame[20] [2]), .O(n28329));
    defparam i15266_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i2_2_lut_adj_1515 (.I0(\data_out_frame[18][2] ), .I1(\data_out_frame[18]_c [1]), 
            .I2(GND_net), .I3(GND_net), .O(n7_adj_4340));
    defparam i2_2_lut_adj_1515.LUT_INIT = 16'h6666;
    SB_LUT4 i4_4_lut_adj_1516 (.I0(n7_adj_4340), .I1(n41615), .I2(n46733), 
            .I3(n44351), .O(n42361));
    defparam i4_4_lut_adj_1516.LUT_INIT = 16'h9669;
    SB_LUT4 i15267_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44085), .I2(rx_data[1]), 
            .I3(\data_in_frame[20] [1]), .O(n28330));
    defparam i15267_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1517 (.I0(\data_out_frame[18][2] ), .I1(n44697), 
            .I2(n42361), .I3(n27138), .O(n44503));
    defparam i3_4_lut_adj_1517.LUT_INIT = 16'h9669;
    SB_LUT4 i1418_2_lut (.I0(\data_out_frame[20] [7]), .I1(\data_out_frame[20] [6]), 
            .I2(GND_net), .I3(GND_net), .O(n2206));   // verilog/coms.v(78[16:27])
    defparam i1418_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i6_4_lut_adj_1518 (.I0(n41571), .I1(n2206), .I2(n44491), .I3(n44204), 
            .O(n16_adj_4341));
    defparam i6_4_lut_adj_1518.LUT_INIT = 16'h6996;
    SB_LUT4 i7_4_lut_adj_1519 (.I0(\data_out_frame[23] [0]), .I1(n44318), 
            .I2(n44503), .I3(n50676), .O(n17_adj_4342));
    defparam i7_4_lut_adj_1519.LUT_INIT = 16'h9669;
    SB_LUT4 i9_4_lut_adj_1520 (.I0(n17_adj_4342), .I1(n42416), .I2(n16_adj_4341), 
            .I3(n42438), .O(n46282));
    defparam i9_4_lut_adj_1520.LUT_INIT = 16'h9669;
    SB_LUT4 i15268_3_lut_4_lut (.I0(n8_adj_4175), .I1(n44085), .I2(rx_data[0]), 
            .I3(\data_in_frame[20] [0]), .O(n28331));
    defparam i15268_3_lut_4_lut.LUT_INIT = 16'hfe10;
    SB_LUT4 i3_4_lut_adj_1521 (.I0(\data_out_frame[25] [1]), .I1(\data_out_frame[25] [2]), 
            .I2(n46282), .I3(n41225), .O(n45719));
    defparam i3_4_lut_adj_1521.LUT_INIT = 16'h6996;
    uart_tx tx (.CLK_c(CLK_c), .GND_net(GND_net), .tx_o(tx_o), .tx_data({tx_data}), 
            .VCC_net(VCC_net), .tx_active(tx_active), .\r_SM_Main_2__N_3516[0] (r_SM_Main_2__N_3516[0]), 
            .tx_enable(tx_enable)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(107[10:70])
    uart_rx rx (.CLK_c(CLK_c), .r_SM_Main({r_SM_Main}), .\r_SM_Main_2__N_3442[2] (\r_SM_Main_2__N_3442[2] ), 
            .r_Bit_Index({Open_36, Open_37, \r_Bit_Index[0] }), .n26629(n26629), 
            .GND_net(GND_net), .n4(n4), .r_Rx_Data(r_Rx_Data), .RX_N_10(RX_N_10), 
            .n27846(n27846), .VCC_net(VCC_net), .n28246(n28246), .n43659(n43659), 
            .rx_data_ready(rx_data_ready), .n28250(n28250), .rx_data({rx_data}), 
            .n28223(n28223), .n28222(n28222), .n28221(n28221), .n28219(n28219), 
            .n28218(n28218), .n43968(n43968), .n28203(n28203), .n28202(n28202), 
            .n44048(n44048), .n4_adj_8(n4_adj_10), .n4_adj_9(n4_adj_11), 
            .n26624(n26624), .n33765(n33765)) /* synthesis syn_module_defined=1 */ ;   // verilog/coms.v(93[10:44])
    
endmodule
//
// Verilog Description of module uart_tx
//

module uart_tx (CLK_c, GND_net, tx_o, tx_data, VCC_net, tx_active, 
            \r_SM_Main_2__N_3516[0] , tx_enable) /* synthesis syn_module_defined=1 */ ;
    input CLK_c;
    input GND_net;
    output tx_o;
    input [7:0]tx_data;
    input VCC_net;
    output tx_active;
    input \r_SM_Main_2__N_3516[0] ;
    output tx_enable;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [8:0]n41;
    
    wire n1;
    wire [8:0]r_Clock_Count;   // verilog/uart_tx.v(32[16:29])
    
    wire n28121, n27839;
    wire [2:0]r_Bit_Index;   // verilog/uart_tx.v(33[16:27])
    wire [2:0]r_SM_Main;   // verilog/uart_tx.v(31[16:25])
    
    wire n28486, n3, n23923;
    wire [7:0]r_Tx_Data;   // verilog/uart_tx.v(34[16:25])
    
    wire n19902, n38370, n28052;
    wire [2:0]n307;
    
    wire n3_adj_4110, n40467, n40466, n40465, n40464, n40463, n40462, 
        n40461, n40460, n45407, n48973, n48974, n10, n43699, n48980, 
        n48979, n45691;
    wire [2:0]r_SM_Main_2__N_3513;
    
    wire n51519, n51522, n43971, n21, n4, n19244;
    
    SB_DFFESR r_Clock_Count_1552__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(n1), 
            .D(n41[3]), .R(n28121));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1552__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(n1), 
            .D(n41[2]), .R(n28121));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1552__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(n1), 
            .D(n41[0]), .R(n28121));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1552__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(n1), 
            .D(n41[1]), .R(n28121));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i17465_3_lut (.I0(n27839), .I1(r_Bit_Index[0]), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n28486));   // verilog/uart_tx.v(33[16:27])
    defparam i17465_3_lut.LUT_INIT = 16'h6464;
    SB_DFFE o_Tx_Serial_45 (.Q(tx_o), .C(CLK_c), .E(n1), .D(n3));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i0 (.Q(r_Tx_Data[0]), .C(CLK_c), .E(n23923), .D(tx_data[0]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n19902), .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index[1]), .C(CLK_c), .E(n27839), 
            .D(n38370), .R(n28052));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index[2]), .C(CLK_c), .E(n27839), 
            .D(n307[2]), .R(n28052));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n3_adj_4110), 
            .R(r_SM_Main[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i7 (.Q(r_Tx_Data[7]), .C(CLK_c), .E(n23923), .D(tx_data[7]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i6 (.Q(r_Tx_Data[6]), .C(CLK_c), .E(n23923), .D(tx_data[6]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i5 (.Q(r_Tx_Data[5]), .C(CLK_c), .E(n23923), .D(tx_data[5]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i4 (.Q(r_Tx_Data[4]), .C(CLK_c), .E(n23923), .D(tx_data[4]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i3 (.Q(r_Tx_Data[3]), .C(CLK_c), .E(n23923), .D(tx_data[3]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i2 (.Q(r_Tx_Data[2]), .C(CLK_c), .E(n23923), .D(tx_data[2]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFE r_Tx_Data_i1 (.Q(r_Tx_Data[1]), .C(CLK_c), .E(n23923), .D(tx_data[1]));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 r_Clock_Count_1552_add_4_10_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[8]), .I3(n40467), .O(n41[8])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1552_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1552_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n40466), .O(n41[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1552_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1552_add_4_9 (.CI(n40466), .I0(GND_net), .I1(r_Clock_Count[7]), 
            .CO(n40467));
    SB_LUT4 r_Clock_Count_1552_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n40465), .O(n41[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1552_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1552_add_4_8 (.CI(n40465), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n40466));
    SB_LUT4 r_Clock_Count_1552_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n40464), .O(n41[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1552_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1552_add_4_7 (.CI(n40464), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n40465));
    SB_LUT4 r_Clock_Count_1552_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n40463), .O(n41[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1552_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1552_add_4_6 (.CI(n40463), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n40464));
    SB_LUT4 r_Clock_Count_1552_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n40462), .O(n41[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1552_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1552_add_4_5 (.CI(n40462), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n40463));
    SB_LUT4 r_Clock_Count_1552_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n40461), .O(n41[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1552_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1552_add_4_4 (.CI(n40461), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n40462));
    SB_LUT4 r_Clock_Count_1552_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n40460), .O(n41[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1552_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1552_add_4_3 (.CI(n40460), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n40461));
    SB_LUT4 r_Clock_Count_1552_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n41[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1552_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1552_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n40460));
    SB_DFFESR r_Clock_Count_1552__i8 (.Q(r_Clock_Count[8]), .C(CLK_c), .E(n1), 
            .D(n41[8]), .R(n28121));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1552__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .E(n1), 
            .D(n41[7]), .R(n28121));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1552__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(n1), 
            .D(n41[6]), .R(n28121));   // verilog/uart_tx.v(118[34:51])
    SB_DFFESR r_Clock_Count_1552__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(n1), 
            .D(n41[5]), .R(n28121));   // verilog/uart_tx.v(118[34:51])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n45407));   // verilog/uart_tx.v(40[10] 143[8])
    SB_DFFESR r_Clock_Count_1552__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(n1), 
            .D(n41[4]), .R(n28121));   // verilog/uart_tx.v(118[34:51])
    SB_LUT4 i34021_3_lut (.I0(r_Tx_Data[0]), .I1(r_Tx_Data[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n48973));
    defparam i34021_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34022_3_lut (.I0(r_Tx_Data[2]), .I1(r_Tx_Data[3]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n48974));
    defparam i34022_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i4_4_lut (.I0(r_Clock_Count[6]), .I1(r_Clock_Count[4]), .I2(r_Clock_Count[5]), 
            .I3(r_Clock_Count[7]), .O(n10));   // verilog/uart_tx.v(32[16:29])
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF r_Tx_Active_47 (.Q(tx_active), .C(CLK_c), .D(n43699));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i34028_3_lut (.I0(r_Tx_Data[6]), .I1(r_Tx_Data[7]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n48980));
    defparam i34028_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i34027_3_lut (.I0(r_Tx_Data[4]), .I1(r_Tx_Data[5]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n48979));
    defparam i34027_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i35129_3_lut (.I0(r_Bit_Index[2]), .I1(r_Bit_Index[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n307[2]));
    defparam i35129_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i3_4_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[2]), .I2(r_Clock_Count[1]), 
            .I3(r_Clock_Count[0]), .O(n45691));   // verilog/uart_tx.v(32[16:29])
    defparam i3_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(n45691), .I1(n10), .I2(r_Clock_Count[8]), .I3(GND_net), 
            .O(r_SM_Main_2__N_3513[1]));   // verilog/uart_tx.v(32[16:29])
    defparam i5_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i28_2_lut (.I0(r_Bit_Index[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n38370));   // verilog/uart_tx.v(33[16:27])
    defparam i28_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i1_1_lut (.I0(r_SM_Main[2]), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(n1));
    defparam i1_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 r_Bit_Index_1__bdd_4_lut (.I0(r_Bit_Index[1]), .I1(n48979), 
            .I2(n48980), .I3(r_Bit_Index[2]), .O(n51519));
    defparam r_Bit_Index_1__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n51519_bdd_4_lut (.I0(n51519), .I1(n48974), .I2(n48973), .I3(r_Bit_Index[2]), 
            .O(n51522));
    defparam n51519_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_4_lut (.I0(r_Bit_Index[0]), .I1(r_SM_Main_2__N_3513[1]), 
            .I2(r_Bit_Index[1]), .I3(r_Bit_Index[2]), .O(n43971));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i22_3_lut (.I0(\r_SM_Main_2__N_3516[0] ), .I1(n43971), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n21));   // verilog/uart_tx.v(31[16:25])
    defparam i22_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i23_3_lut (.I0(n21), .I1(r_SM_Main_2__N_3513[1]), .I2(r_SM_Main[0]), 
            .I3(GND_net), .O(n19902));   // verilog/uart_tx.v(31[16:25])
    defparam i23_3_lut.LUT_INIT = 16'h3a3a;
    SB_LUT4 i25330_3_lut (.I0(r_SM_Main[0]), .I1(n51522), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // verilog/uart_tx.v(31[16:25])
    defparam i25330_3_lut.LUT_INIT = 16'he5e5;
    SB_LUT4 i1_3_lut_4_lut_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_3513[1]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n4));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_3_lut_4_lut_4_lut.LUT_INIT = 16'h008f;
    SB_LUT4 i2_3_lut_4_lut_4_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_3513[1]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[2]), .O(n45407));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i2_3_lut_4_lut_4_lut.LUT_INIT = 16'h0080;
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(CLK_c), .D(n28486));   // verilog/uart_tx.v(40[10] 143[8])
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(n43971), .O(n28052));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i1_3_lut_4_lut_adj_851 (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main_2__N_3513[1]), .O(n27839));
    defparam i1_3_lut_4_lut_adj_851.LUT_INIT = 16'h1101;
    SB_LUT4 i2_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(\r_SM_Main_2__N_3516[0] ), .O(n23923));
    defparam i2_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_LUT4 i24_2_lut_3_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_3513[1]), 
            .I2(r_SM_Main[1]), .I3(GND_net), .O(n3_adj_4110));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i24_2_lut_3_lut.LUT_INIT = 16'h7878;
    SB_LUT4 i15058_4_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main_2__N_3513[1]), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n28121));   // verilog/uart_tx.v(118[34:51])
    defparam i15058_4_lut_4_lut.LUT_INIT = 16'h4445;
    SB_LUT4 i1_2_lut (.I0(r_SM_Main[0]), .I1(\r_SM_Main_2__N_3516[0] ), 
            .I2(GND_net), .I3(GND_net), .O(n19244));   // verilog/uart_tx.v(40[10] 143[8])
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i12_4_lut (.I0(tx_active), .I1(r_SM_Main[1]), .I2(n19244), 
            .I3(n4), .O(n43699));   // verilog/uart_tx.v(31[16:25])
    defparam i12_4_lut.LUT_INIT = 16'h32aa;
    SB_LUT4 o_Tx_Serial_I_0_1_lut (.I0(tx_o), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(tx_enable));   // verilog/uart_tx.v(38[24:36])
    defparam o_Tx_Serial_I_0_1_lut.LUT_INIT = 16'h5555;
    
endmodule
//
// Verilog Description of module uart_rx
//

module uart_rx (CLK_c, r_SM_Main, \r_SM_Main_2__N_3442[2] , r_Bit_Index, 
            n26629, GND_net, n4, r_Rx_Data, RX_N_10, n27846, VCC_net, 
            n28246, n43659, rx_data_ready, n28250, rx_data, n28223, 
            n28222, n28221, n28219, n28218, n43968, n28203, n28202, 
            n44048, n4_adj_8, n4_adj_9, n26624, n33765) /* synthesis syn_module_defined=1 */ ;
    input CLK_c;
    output [2:0]r_SM_Main;
    output \r_SM_Main_2__N_3442[2] ;
    output [2:0]r_Bit_Index;
    output n26629;
    input GND_net;
    output n4;
    output r_Rx_Data;
    input RX_N_10;
    output n27846;
    input VCC_net;
    input n28246;
    input n43659;
    output rx_data_ready;
    input n28250;
    output [7:0]rx_data;
    input n28223;
    input n28222;
    input n28221;
    input n28219;
    input n28218;
    output n43968;
    input n28203;
    input n28202;
    input n44048;
    output n4_adj_8;
    output n4_adj_9;
    output n26624;
    output n33765;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [7:0]n37;
    
    wire n27913;
    wire [7:0]r_Clock_Count;   // verilog/uart_rx.v(32[17:30])
    
    wire n28119, n26493;
    wire [2:0]r_Bit_Index_c;   // verilog/uart_rx.v(33[17:28])
    
    wire n3, r_Rx_Data_R;
    wire [2:0]n326;
    
    wire n28054, n34535, n40459, n40458, n40457, n40456, n40455, 
        n40454, n40453, n48659, n26485;
    wire [2:0]r_SM_Main_2__N_3448;
    
    wire n6, n49791, n49789, n6_adj_4107, n49770;
    wire [2:0]r_SM_Main_2__N_3445;
    
    wire n34405, n1;
    
    SB_DFFESR r_Clock_Count_1550__i0 (.Q(r_Clock_Count[0]), .C(CLK_c), .E(n27913), 
            .D(n37[0]), .R(n28119));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1550__i7 (.Q(r_Clock_Count[7]), .C(CLK_c), .E(n27913), 
            .D(n37[7]), .R(n28119));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1550__i6 (.Q(r_Clock_Count[6]), .C(CLK_c), .E(n27913), 
            .D(n37[6]), .R(n28119));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1550__i5 (.Q(r_Clock_Count[5]), .C(CLK_c), .E(n27913), 
            .D(n37[5]), .R(n28119));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1550__i4 (.Q(r_Clock_Count[4]), .C(CLK_c), .E(n27913), 
            .D(n37[4]), .R(n28119));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1550__i3 (.Q(r_Clock_Count[3]), .C(CLK_c), .E(n27913), 
            .D(n37[3]), .R(n28119));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1550__i2 (.Q(r_Clock_Count[2]), .C(CLK_c), .E(n27913), 
            .D(n37[2]), .R(n28119));   // verilog/uart_rx.v(120[34:51])
    SB_DFFESR r_Clock_Count_1550__i1 (.Q(r_Clock_Count[1]), .C(CLK_c), .E(n27913), 
            .D(n37[1]), .R(n28119));   // verilog/uart_rx.v(120[34:51])
    SB_LUT4 i3_4_lut (.I0(r_SM_Main[1]), .I1(r_SM_Main[2]), .I2(r_SM_Main[0]), 
            .I3(\r_SM_Main_2__N_3442[2] ), .O(n26493));
    defparam i3_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i1_2_lut (.I0(n26493), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n26629));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 equal_156_i4_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4));   // verilog/uart_rx.v(97[17:39])
    defparam equal_156_i4_2_lut.LUT_INIT = 16'heeee;
    SB_DFFSR r_SM_Main_i0 (.Q(r_SM_Main[0]), .C(CLK_c), .D(n3), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Data_50 (.Q(r_Rx_Data), .C(CLK_c), .D(r_Rx_Data_R));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFF r_Rx_Data_R_49 (.Q(r_Rx_Data_R), .C(CLK_c), .D(RX_N_10));   // verilog/uart_rx.v(41[10] 45[8])
    SB_DFFESR r_Bit_Index_i1 (.Q(r_Bit_Index_c[1]), .C(CLK_c), .E(n27846), 
            .D(n326[1]), .R(n28054));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFESR r_Bit_Index_i2 (.Q(r_Bit_Index_c[2]), .C(CLK_c), .E(n27846), 
            .D(n326[2]), .R(n28054));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFFSR r_SM_Main_i1 (.Q(r_SM_Main[1]), .C(CLK_c), .D(n34535), .R(r_SM_Main[2]));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 r_Clock_Count_1550_add_4_9_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[7]), .I3(n40459), .O(n37[7])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1550_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 r_Clock_Count_1550_add_4_8_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[6]), .I3(n40458), .O(n37[6])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1550_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1550_add_4_8 (.CI(n40458), .I0(GND_net), .I1(r_Clock_Count[6]), 
            .CO(n40459));
    SB_LUT4 r_Clock_Count_1550_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[5]), .I3(n40457), .O(n37[5])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1550_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1550_add_4_7 (.CI(n40457), .I0(GND_net), .I1(r_Clock_Count[5]), 
            .CO(n40458));
    SB_LUT4 r_Clock_Count_1550_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[4]), .I3(n40456), .O(n37[4])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1550_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1550_add_4_6 (.CI(n40456), .I0(GND_net), .I1(r_Clock_Count[4]), 
            .CO(n40457));
    SB_LUT4 r_Clock_Count_1550_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[3]), .I3(n40455), .O(n37[3])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1550_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1550_add_4_5 (.CI(n40455), .I0(GND_net), .I1(r_Clock_Count[3]), 
            .CO(n40456));
    SB_LUT4 r_Clock_Count_1550_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[2]), .I3(n40454), .O(n37[2])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1550_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1550_add_4_4 (.CI(n40454), .I0(GND_net), .I1(r_Clock_Count[2]), 
            .CO(n40455));
    SB_LUT4 r_Clock_Count_1550_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[1]), .I3(n40453), .O(n37[1])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1550_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1550_add_4_3 (.CI(n40453), .I0(GND_net), .I1(r_Clock_Count[1]), 
            .CO(n40454));
    SB_LUT4 r_Clock_Count_1550_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(r_Clock_Count[0]), .I3(VCC_net), .O(n37[0])) /* synthesis syn_instantiated=1 */ ;
    defparam r_Clock_Count_1550_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY r_Clock_Count_1550_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(r_Clock_Count[0]), 
            .CO(n40453));
    SB_LUT4 i33767_2_lut (.I0(r_Clock_Count[0]), .I1(r_Clock_Count[2]), 
            .I2(GND_net), .I3(GND_net), .O(n48659));
    defparam i33767_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i4_4_lut (.I0(n48659), .I1(n26485), .I2(r_Clock_Count[3]), 
            .I3(r_Clock_Count[1]), .O(r_SM_Main_2__N_3448[0]));
    defparam i4_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i2_2_lut (.I0(r_Clock_Count[3]), .I1(r_Clock_Count[2]), .I2(GND_net), 
            .I3(GND_net), .O(n6));
    defparam i2_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i21242_4_lut (.I0(r_Clock_Count[0]), .I1(n26485), .I2(n6), 
            .I3(r_Clock_Count[1]), .O(\r_SM_Main_2__N_3442[2] ));
    defparam i21242_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i3_4_lut_adj_847 (.I0(r_Clock_Count[4]), .I1(r_Clock_Count[7]), 
            .I2(r_Clock_Count[6]), .I3(r_Clock_Count[5]), .O(n26485));   // verilog/uart_rx.v(68[17:52])
    defparam i3_4_lut_adj_847.LUT_INIT = 16'hfffe;
    SB_LUT4 i34964_4_lut (.I0(r_Rx_Data), .I1(r_Clock_Count[1]), .I2(n26485), 
            .I3(r_Clock_Count[3]), .O(n49791));
    defparam i34964_4_lut.LUT_INIT = 16'h0004;
    SB_LUT4 i35090_3_lut (.I0(n49791), .I1(r_SM_Main[0]), .I2(n48659), 
            .I3(GND_net), .O(n49789));
    defparam i35090_3_lut.LUT_INIT = 16'hb3b3;
    SB_LUT4 i1_4_lut (.I0(r_SM_Main[2]), .I1(n49789), .I2(\r_SM_Main_2__N_3442[2] ), 
            .I3(r_SM_Main[1]), .O(n28119));
    defparam i1_4_lut.LUT_INIT = 16'h5044;
    SB_LUT4 i2_2_lut_adj_848 (.I0(r_SM_Main_2__N_3448[0]), .I1(r_SM_Main[0]), 
            .I2(GND_net), .I3(GND_net), .O(n6_adj_4107));
    defparam i2_2_lut_adj_848.LUT_INIT = 16'h4444;
    SB_LUT4 i35747_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[1]), .I2(n6_adj_4107), 
            .I3(r_Rx_Data), .O(n27913));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i35747_4_lut.LUT_INIT = 16'h4555;
    SB_DFF r_Bit_Index_i0 (.Q(r_Bit_Index[0]), .C(CLK_c), .D(n28246));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_DV_52 (.Q(rx_data_ready), .C(CLK_c), .D(n43659));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i0 (.Q(rx_data[0]), .C(CLK_c), .D(n28250));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i34963_3_lut (.I0(r_SM_Main[0]), .I1(r_SM_Main_2__N_3448[0]), 
            .I2(r_Rx_Data), .I3(GND_net), .O(n49770));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i34963_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_1_i3_4_lut (.I0(n49770), .I1(\r_SM_Main_2__N_3442[2] ), 
            .I2(r_SM_Main[1]), .I3(r_SM_Main[0]), .O(n34535));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_1_i3_4_lut.LUT_INIT = 16'h35f5;
    SB_DFF r_Rx_Byte_i7 (.Q(rx_data[7]), .C(CLK_c), .D(n28223));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i6 (.Q(rx_data[6]), .C(CLK_c), .D(n28222));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i5 (.Q(rx_data[5]), .C(CLK_c), .D(n28221));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i4 (.Q(rx_data[4]), .C(CLK_c), .D(n28219));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i3 (.Q(rx_data[3]), .C(CLK_c), .D(n28218));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1669_3_lut (.I0(r_Bit_Index_c[2]), .I1(r_Bit_Index_c[1]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n326[2]));   // verilog/uart_rx.v(102[36:51])
    defparam i1669_3_lut.LUT_INIT = 16'h6a6a;
    SB_LUT4 i1662_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n326[1]));   // verilog/uart_rx.v(102[36:51])
    defparam i1662_2_lut.LUT_INIT = 16'h6666;
    SB_LUT4 i2_3_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), .I2(r_Bit_Index[0]), 
            .I3(GND_net), .O(n43968));
    defparam i2_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i2_3_lut (.I0(r_SM_Main_2__N_3445[0]), 
            .I1(\r_SM_Main_2__N_3442[2] ), .I2(r_SM_Main[0]), .I3(GND_net), 
            .O(n34405));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i2_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i1_3_lut (.I0(r_Rx_Data), .I1(r_SM_Main_2__N_3448[0]), 
            .I2(r_SM_Main[0]), .I3(GND_net), .O(n1));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i1_3_lut.LUT_INIT = 16'hc5c5;
    SB_LUT4 r_SM_Main_2__I_0_56_Mux_0_i3_3_lut (.I0(n1), .I1(n34405), .I2(r_SM_Main[1]), 
            .I3(GND_net), .O(n3));   // verilog/uart_rx.v(52[7] 143[14])
    defparam r_SM_Main_2__I_0_56_Mux_0_i3_3_lut.LUT_INIT = 16'h3a3a;
    SB_DFF r_Rx_Byte_i2 (.Q(rx_data[2]), .C(CLK_c), .D(n28203));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_Rx_Byte_i1 (.Q(rx_data[1]), .C(CLK_c), .D(n28202));   // verilog/uart_rx.v(49[10] 144[8])
    SB_DFF r_SM_Main_i2 (.Q(r_SM_Main[2]), .C(CLK_c), .D(n44048));   // verilog/uart_rx.v(49[10] 144[8])
    SB_LUT4 i1_3_lut_4_lut (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), .I2(r_SM_Main[1]), 
            .I3(r_SM_Main_2__N_3445[0]), .O(n28054));
    defparam i1_3_lut_4_lut.LUT_INIT = 16'h1101;
    SB_LUT4 i1_3_lut_4_lut_adj_849 (.I0(r_SM_Main[2]), .I1(r_SM_Main[0]), 
            .I2(r_SM_Main[1]), .I3(\r_SM_Main_2__N_3442[2] ), .O(n27846));
    defparam i1_3_lut_4_lut_adj_849.LUT_INIT = 16'h1101;
    SB_LUT4 i21414_2_lut_4_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(r_Bit_Index[0]), .I3(\r_SM_Main_2__N_3442[2] ), .O(r_SM_Main_2__N_3445[0]));
    defparam i21414_2_lut_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 equal_154_i4_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_8));   // verilog/uart_rx.v(97[17:39])
    defparam equal_154_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 equal_152_i4_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(GND_net), .I3(GND_net), .O(n4_adj_9));   // verilog/uart_rx.v(97[17:39])
    defparam equal_152_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1_2_lut_adj_850 (.I0(n26493), .I1(r_Bit_Index[0]), .I2(GND_net), 
            .I3(GND_net), .O(n26624));   // verilog/uart_rx.v(52[7] 143[14])
    defparam i1_2_lut_adj_850.LUT_INIT = 16'hbbbb;
    SB_LUT4 i20715_2_lut (.I0(r_Bit_Index_c[1]), .I1(r_Bit_Index_c[2]), 
            .I2(GND_net), .I3(GND_net), .O(n33765));
    defparam i20715_2_lut.LUT_INIT = 16'h8888;
    
endmodule
//
// Verilog Description of module EEPROM
//

module EEPROM (CLK_c, n4226, \state[1] , GND_net, \state[0] , read, 
            \state[2] , n7, \state[3] , n6, n28217, rw, n43797, 
            data_ready, enable_slow_N_4090, n43693, n43685, n44859, 
            n44120, n34334, VCC_net, n5538, n33769, n4, scl_enable, 
            \state_7__N_4003[3] , n6014, \state_7__N_3987[0] , sda_enable, 
            n4_adj_4, \saved_addr[0] , \state[0]_adj_5 , n10, n10_adj_6, 
            n8, n28230, data, n10_adj_7, n28224, scl, sda_out, 
            n28207, n28206, n28205, n28204, n28200, n28199, n28198, 
            n26650, n26645, n49785) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input CLK_c;
    output [0:0]n4226;
    output \state[1] ;
    input GND_net;
    output \state[0] ;
    input read;
    output \state[2] ;
    output n7;
    output \state[3] ;
    output n6;
    input n28217;
    output rw;
    input n43797;
    output data_ready;
    output enable_slow_N_4090;
    input n43693;
    input n43685;
    input n44859;
    output n44120;
    output n34334;
    input VCC_net;
    output n5538;
    output n33769;
    output n4;
    output scl_enable;
    input \state_7__N_4003[3] ;
    input n6014;
    output \state_7__N_3987[0] ;
    output sda_enable;
    output n4_adj_4;
    output \saved_addr[0] ;
    output \state[0]_adj_5 ;
    output n10;
    output n10_adj_6;
    input n8;
    input n28230;
    output [7:0]data;
    input n10_adj_7;
    input n28224;
    output scl;
    output sda_out;
    input n28207;
    input n28206;
    input n28205;
    input n28204;
    input n28200;
    input n28199;
    input n28198;
    output n26650;
    output n26645;
    output n49785;
    
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [15:0]delay_counter_15__N_3889;
    
    wire n27876;
    wire [15:0]delay_counter;   // verilog/eeprom.v(24[12:25])
    
    wire n28073, enable;
    wire [15:0]n3652;
    
    wire n39178, n39177;
    wire [7:0]state;   // verilog/i2c_controller.v(33[12:17])
    
    wire n39176, n39175, n39174, n39173, n39172, n39171, n39170, 
        n26478, n39169, n39168, n39167, n39166, n39165, n39164, 
        n28, n26, n27, n25;
    
    SB_DFFESR delay_counter_i0_i1 (.Q(delay_counter[1]), .C(CLK_c), .E(n27876), 
            .D(delay_counter_15__N_3889[1]), .R(n28073));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i2 (.Q(delay_counter[2]), .C(CLK_c), .E(n27876), 
            .D(delay_counter_15__N_3889[2]), .R(n28073));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i3 (.Q(delay_counter[3]), .C(CLK_c), .E(n27876), 
            .D(delay_counter_15__N_3889[3]), .R(n28073));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i4 (.Q(delay_counter[4]), .C(CLK_c), .E(n27876), 
            .D(delay_counter_15__N_3889[4]), .S(n28073));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i5 (.Q(delay_counter[5]), .C(CLK_c), .E(n27876), 
            .D(delay_counter_15__N_3889[5]), .R(n28073));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i6 (.Q(delay_counter[6]), .C(CLK_c), .E(n27876), 
            .D(delay_counter_15__N_3889[6]), .S(n28073));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i7 (.Q(delay_counter[7]), .C(CLK_c), .E(n27876), 
            .D(delay_counter_15__N_3889[7]), .S(n28073));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i8 (.Q(delay_counter[8]), .C(CLK_c), .E(n27876), 
            .D(delay_counter_15__N_3889[8]), .S(n28073));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i9 (.Q(delay_counter[9]), .C(CLK_c), .E(n27876), 
            .D(delay_counter_15__N_3889[9]), .S(n28073));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESS delay_counter_i0_i10 (.Q(delay_counter[10]), .C(CLK_c), .E(n27876), 
            .D(delay_counter_15__N_3889[10]), .S(n28073));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i11 (.Q(delay_counter[11]), .C(CLK_c), .E(n27876), 
            .D(delay_counter_15__N_3889[11]), .R(n28073));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i12 (.Q(delay_counter[12]), .C(CLK_c), .E(n27876), 
            .D(delay_counter_15__N_3889[12]), .R(n28073));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i13 (.Q(delay_counter[13]), .C(CLK_c), .E(n27876), 
            .D(delay_counter_15__N_3889[13]), .R(n28073));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i14 (.Q(delay_counter[14]), .C(CLK_c), .E(n27876), 
            .D(delay_counter_15__N_3889[14]), .R(n28073));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i15 (.Q(delay_counter[15]), .C(CLK_c), .E(n27876), 
            .D(delay_counter_15__N_3889[15]), .R(n28073));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFSR enable_39 (.Q(enable), .C(CLK_c), .D(n4226[0]), .R(\state[1] ));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 add_714_17_lut (.I0(GND_net), .I1(delay_counter[15]), .I2(n3652[5]), 
            .I3(n39178), .O(delay_counter_15__N_3889[15])) /* synthesis syn_instantiated=1 */ ;
    defparam add_714_17_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i15023_2_lut (.I0(n27876), .I1(\state[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n28073));   // verilog/eeprom.v(26[8] 58[4])
    defparam i15023_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i1_3_lut (.I0(read), .I1(\state[1] ), .I2(\state[0] ), .I3(GND_net), 
            .O(n27876));
    defparam i1_3_lut.LUT_INIT = 16'h3232;
    SB_LUT4 add_714_16_lut (.I0(GND_net), .I1(delay_counter[14]), .I2(n3652[5]), 
            .I3(n39177), .O(delay_counter_15__N_3889[14])) /* synthesis syn_instantiated=1 */ ;
    defparam add_714_16_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_2_lut (.I0(state[1]), .I1(\state[2] ), .I2(GND_net), .I3(GND_net), 
            .O(n7));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_CARRY add_714_16 (.CI(n39177), .I0(delay_counter[14]), .I1(n3652[5]), 
            .CO(n39178));
    SB_LUT4 add_714_15_lut (.I0(GND_net), .I1(delay_counter[13]), .I2(n3652[5]), 
            .I3(n39176), .O(delay_counter_15__N_3889[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_714_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_714_15 (.CI(n39176), .I0(delay_counter[13]), .I1(n3652[5]), 
            .CO(n39177));
    SB_LUT4 add_714_14_lut (.I0(GND_net), .I1(delay_counter[12]), .I2(n3652[5]), 
            .I3(n39175), .O(delay_counter_15__N_3889[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_714_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_714_14 (.CI(n39175), .I0(delay_counter[12]), .I1(n3652[5]), 
            .CO(n39176));
    SB_LUT4 add_714_13_lut (.I0(GND_net), .I1(delay_counter[11]), .I2(n3652[5]), 
            .I3(n39174), .O(delay_counter_15__N_3889[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_714_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_714_13 (.CI(n39174), .I0(delay_counter[11]), .I1(n3652[5]), 
            .CO(n39175));
    SB_LUT4 add_714_12_lut (.I0(GND_net), .I1(delay_counter[10]), .I2(n3652[5]), 
            .I3(n39173), .O(delay_counter_15__N_3889[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_714_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_714_12 (.CI(n39173), .I0(delay_counter[10]), .I1(n3652[5]), 
            .CO(n39174));
    SB_LUT4 add_714_11_lut (.I0(GND_net), .I1(delay_counter[9]), .I2(n3652[5]), 
            .I3(n39172), .O(delay_counter_15__N_3889[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_714_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_714_11 (.CI(n39172), .I0(delay_counter[9]), .I1(n3652[5]), 
            .CO(n39173));
    SB_LUT4 add_714_10_lut (.I0(GND_net), .I1(delay_counter[8]), .I2(n3652[5]), 
            .I3(n39171), .O(delay_counter_15__N_3889[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_714_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_714_10 (.CI(n39171), .I0(delay_counter[8]), .I1(n3652[5]), 
            .CO(n39172));
    SB_LUT4 add_714_9_lut (.I0(GND_net), .I1(delay_counter[7]), .I2(n3652[5]), 
            .I3(n39170), .O(delay_counter_15__N_3889[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_714_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_714_9 (.CI(n39170), .I0(delay_counter[7]), .I1(n3652[5]), 
            .CO(n39171));
    SB_LUT4 i2_2_lut_adj_846 (.I0(n26478), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n6));   // verilog/eeprom.v(42[12:28])
    defparam i2_2_lut_adj_846.LUT_INIT = 16'heeee;
    SB_LUT4 add_714_8_lut (.I0(GND_net), .I1(delay_counter[6]), .I2(n3652[5]), 
            .I3(n39169), .O(delay_counter_15__N_3889[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_714_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_714_8 (.CI(n39169), .I0(delay_counter[6]), .I1(n3652[5]), 
            .CO(n39170));
    SB_LUT4 add_714_7_lut (.I0(GND_net), .I1(delay_counter[5]), .I2(n3652[5]), 
            .I3(n39168), .O(delay_counter_15__N_3889[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_714_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_714_7 (.CI(n39168), .I0(delay_counter[5]), .I1(n3652[5]), 
            .CO(n39169));
    SB_LUT4 add_714_6_lut (.I0(GND_net), .I1(delay_counter[4]), .I2(n3652[5]), 
            .I3(n39167), .O(delay_counter_15__N_3889[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_714_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_714_6 (.CI(n39167), .I0(delay_counter[4]), .I1(n3652[5]), 
            .CO(n39168));
    SB_LUT4 add_714_5_lut (.I0(GND_net), .I1(delay_counter[3]), .I2(n3652[5]), 
            .I3(n39166), .O(delay_counter_15__N_3889[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_714_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_714_5 (.CI(n39166), .I0(delay_counter[3]), .I1(n3652[5]), 
            .CO(n39167));
    SB_LUT4 add_714_4_lut (.I0(GND_net), .I1(delay_counter[2]), .I2(n3652[5]), 
            .I3(n39165), .O(delay_counter_15__N_3889[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_714_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_714_4 (.CI(n39165), .I0(delay_counter[2]), .I1(n3652[5]), 
            .CO(n39166));
    SB_LUT4 add_714_3_lut (.I0(GND_net), .I1(delay_counter[1]), .I2(n3652[5]), 
            .I3(n39164), .O(delay_counter_15__N_3889[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_714_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_714_3 (.CI(n39164), .I0(delay_counter[1]), .I1(n3652[5]), 
            .CO(n39165));
    SB_LUT4 add_714_2_lut (.I0(GND_net), .I1(delay_counter[0]), .I2(n3652[5]), 
            .I3(GND_net), .O(delay_counter_15__N_3889[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_714_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_714_2 (.CI(GND_net), .I0(delay_counter[0]), .I1(n3652[5]), 
            .CO(n39164));
    SB_DFF rw_43 (.Q(rw), .C(CLK_c), .D(n28217));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF data_ready_42 (.Q(data_ready), .C(CLK_c), .D(n43797));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFFESR delay_counter_i0_i0 (.Q(delay_counter[0]), .C(CLK_c), .E(n27876), 
            .D(delay_counter_15__N_3889[0]), .R(n28073));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i35801_2_lut (.I0(n26478), .I1(enable_slow_N_4090), .I2(GND_net), 
            .I3(GND_net), .O(n3652[5]));   // verilog/eeprom.v(46[18] 48[12])
    defparam i35801_2_lut.LUT_INIT = 16'h2222;
    SB_LUT4 i12_4_lut (.I0(delay_counter[15]), .I1(delay_counter[6]), .I2(delay_counter[2]), 
            .I3(delay_counter[12]), .O(n28));   // verilog/eeprom.v(42[12:28])
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i10_4_lut (.I0(delay_counter[10]), .I1(delay_counter[9]), .I2(delay_counter[8]), 
            .I3(delay_counter[7]), .O(n26));   // verilog/eeprom.v(42[12:28])
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i11_4_lut (.I0(delay_counter[3]), .I1(delay_counter[11]), .I2(delay_counter[1]), 
            .I3(delay_counter[14]), .O(n27));   // verilog/eeprom.v(42[12:28])
    defparam i11_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i9_4_lut (.I0(delay_counter[4]), .I1(delay_counter[0]), .I2(delay_counter[13]), 
            .I3(delay_counter[5]), .O(n25));   // verilog/eeprom.v(42[12:28])
    defparam i9_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i15_4_lut (.I0(n25), .I1(n27), .I2(n26), .I3(n28), .O(n26478));   // verilog/eeprom.v(42[12:28])
    defparam i15_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 mux_906_Mux_0_i1_4_lut (.I0(read), .I1(n26478), .I2(\state[0] ), 
            .I3(enable_slow_N_4090), .O(n4226[0]));   // verilog/eeprom.v(29[3] 57[10])
    defparam mux_906_Mux_0_i1_4_lut.LUT_INIT = 16'h0a3a;
    SB_DFF state__i1 (.Q(\state[1] ), .C(CLK_c), .D(n43693));   // verilog/eeprom.v(26[8] 58[4])
    SB_DFF state__i0 (.Q(\state[0] ), .C(CLK_c), .D(n43685));   // verilog/eeprom.v(26[8] 58[4])
    SB_LUT4 i1_4_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(n44859), 
            .I3(enable_slow_N_4090), .O(n44120));   // verilog/eeprom.v(51[5:9])
    defparam i1_4_lut_4_lut.LUT_INIT = 16'hfcf8;
    SB_LUT4 i21278_2_lut_3_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(enable_slow_N_4090), 
            .I3(GND_net), .O(n34334));   // verilog/eeprom.v(51[5:9])
    defparam i21278_2_lut_3_lut.LUT_INIT = 16'hfbfb;
    i2c_controller i2c (.VCC_net(VCC_net), .GND_net(GND_net), .n5538(n5538), 
            .\state[3] (\state[3] ), .\state[2] (\state[2] ), .\state[1] (state[1]), 
            .CLK_c(CLK_c), .n33769(n33769), .n4(n4), .scl_enable(scl_enable), 
            .\state_7__N_4003[3] (\state_7__N_4003[3] ), .n6014(n6014), 
            .\state_7__N_3987[0] (\state_7__N_3987[0] ), .sda_enable(sda_enable), 
            .n4_adj_1(n4_adj_4), .\saved_addr[0] (\saved_addr[0] ), .\state[0] (\state[0]_adj_5 ), 
            .n10(n10), .n10_adj_2(n10_adj_6), .n8(n8), .n28230(n28230), 
            .data({data}), .n10_adj_3(n10_adj_7), .enable(enable), .enable_slow_N_4090(enable_slow_N_4090), 
            .n28224(n28224), .scl(scl), .sda_out(sda_out), .n28207(n28207), 
            .n28206(n28206), .n28205(n28205), .n28204(n28204), .n28200(n28200), 
            .n28199(n28199), .n28198(n28198), .n26650(n26650), .n26645(n26645), 
            .n49785(n49785)) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;   // verilog/eeprom.v(60[16] 74[4])
    
endmodule
//
// Verilog Description of module i2c_controller
//

module i2c_controller (VCC_net, GND_net, n5538, \state[3] , \state[2] , 
            \state[1] , CLK_c, n33769, n4, scl_enable, \state_7__N_4003[3] , 
            n6014, \state_7__N_3987[0] , sda_enable, n4_adj_1, \saved_addr[0] , 
            \state[0] , n10, n10_adj_2, n8, n28230, data, n10_adj_3, 
            enable, enable_slow_N_4090, n28224, scl, sda_out, n28207, 
            n28206, n28205, n28204, n28200, n28199, n28198, n26650, 
            n26645, n49785) /* synthesis syn_noprune=1, syn_module_defined=1 */ ;
    input VCC_net;
    input GND_net;
    output n5538;
    output \state[3] ;
    output \state[2] ;
    output \state[1] ;
    input CLK_c;
    output n33769;
    output n4;
    output scl_enable;
    input \state_7__N_4003[3] ;
    input n6014;
    output \state_7__N_3987[0] ;
    output sda_enable;
    output n4_adj_1;
    output \saved_addr[0] ;
    output \state[0] ;
    output n10;
    output n10_adj_2;
    input n8;
    input n28230;
    output [7:0]data;
    input n10_adj_3;
    input enable;
    output enable_slow_N_4090;
    input n28224;
    output scl;
    output sda_out;
    input n28207;
    input n28206;
    input n28205;
    input n28204;
    input n28200;
    input n28199;
    input n28198;
    output n26650;
    output n26645;
    output n49785;
    
    wire i2c_clk /* synthesis is_clock=1, SET_AS_NETWORK=\eeprom/i2c/i2c_clk */ ;   // verilog/i2c_controller.v(41[6:13])
    wire CLK_c /* synthesis SET_AS_NETWORK=CLK_c, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(3[9:12])
    wire [7:0]n119;
    wire [7:0]counter;   // verilog/i2c_controller.v(36[12:19])
    
    wire n39363, n39364, n43849, n46193, n33933, n34177, n5, n34447;
    wire [5:0]n29;
    wire [7:0]counter2;   // verilog/i2c_controller.v(37[12:20])
    
    wire n28122, n27956, n28046, n39362, n39361, n39360, n39359, 
        i2c_clk_N_4076, scl_enable_N_4077, n15, n44863, n5531, n37, 
        enable_slow_N_4089, n27854, n40503, n40502, n40501, n40500, 
        n40499, n19384, n5909, n28050, n49887, n43769, sda_out_adj_4092, 
        n10_c, n49774, n49716, n11, n11_adj_4093, n11_adj_4094, 
        n9, n12, n7, state_7__N_3986, n11_adj_4097, n34056, n33_adj_4098, 
        n34_adj_4099, n39, n49793, n39365, n11_adj_4101;
    
    SB_LUT4 sub_39_add_2_7_lut (.I0(GND_net), .I1(counter[5]), .I2(VCC_net), 
            .I3(n39363), .O(n119[5])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_7 (.CI(n39363), .I0(counter[5]), .I1(VCC_net), 
            .CO(n39364));
    SB_DFFESS state_i0_i3 (.Q(\state[3] ), .C(i2c_clk), .E(n5538), .D(n43849), 
            .S(n46193));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i2 (.Q(\state[2] ), .C(i2c_clk), .E(n5538), .D(n33933), 
            .S(n34177));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS state_i0_i1 (.Q(\state[1] ), .C(i2c_clk), .E(n5538), .D(n5), 
            .S(n34447));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_1554_1555__i1 (.Q(counter2[0]), .C(CLK_c), .D(n29[0]), 
            .R(n28122));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFESR counter_i7 (.Q(counter[7]), .C(i2c_clk), .E(n27956), .D(n119[7]), 
            .R(n28046));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i6 (.Q(counter[6]), .C(i2c_clk), .E(n27956), .D(n119[6]), 
            .R(n28046));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i5 (.Q(counter[5]), .C(i2c_clk), .E(n27956), .D(n119[5]), 
            .R(n28046));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i4 (.Q(counter[4]), .C(i2c_clk), .E(n27956), .D(n119[4]), 
            .R(n28046));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESR counter_i3 (.Q(counter[3]), .C(i2c_clk), .E(n27956), .D(n119[3]), 
            .R(n28046));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i2 (.Q(counter[2]), .C(i2c_clk), .E(n27956), .D(n119[2]), 
            .S(n28046));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFESS counter_i1 (.Q(counter[1]), .C(i2c_clk), .E(n27956), .D(n119[1]), 
            .S(n28046));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 sub_39_add_2_6_lut (.I0(GND_net), .I1(counter[4]), .I2(VCC_net), 
            .I3(n39362), .O(n119[4])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_6 (.CI(n39362), .I0(counter[4]), .I1(VCC_net), 
            .CO(n39363));
    SB_LUT4 sub_39_add_2_5_lut (.I0(GND_net), .I1(counter[3]), .I2(VCC_net), 
            .I3(n39361), .O(n119[3])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_5 (.CI(n39361), .I0(counter[3]), .I1(VCC_net), 
            .CO(n39362));
    SB_LUT4 sub_39_add_2_4_lut (.I0(GND_net), .I1(counter[2]), .I2(VCC_net), 
            .I3(n39360), .O(n119[2])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_4 (.CI(n39360), .I0(counter[2]), .I1(VCC_net), 
            .CO(n39361));
    SB_LUT4 sub_39_add_2_3_lut (.I0(GND_net), .I1(counter[1]), .I2(VCC_net), 
            .I3(n39359), .O(n119[1])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i20719_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n33769));
    defparam i20719_2_lut.LUT_INIT = 16'h8888;
    SB_CARRY sub_39_add_2_3 (.CI(n39359), .I0(counter[1]), .I1(VCC_net), 
            .CO(n39360));
    SB_LUT4 sub_39_add_2_2_lut (.I0(GND_net), .I1(counter[0]), .I2(GND_net), 
            .I3(VCC_net), .O(n119[0])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY sub_39_add_2_2 (.CI(VCC_net), .I0(counter[0]), .I1(GND_net), 
            .CO(n39359));
    SB_LUT4 equal_160_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_160_i4_2_lut.LUT_INIT = 16'hbbbb;
    SB_DFF i2c_clk_121 (.Q(i2c_clk), .C(CLK_c), .D(i2c_clk_N_4076));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_DFFN i2c_scl_enable_123 (.Q(scl_enable), .C(i2c_clk), .D(scl_enable_N_4077));   // verilog/i2c_controller.v(76[12] 82[6])
    SB_LUT4 i29978_2_lut (.I0(\state_7__N_4003[3] ), .I1(n15), .I2(GND_net), 
            .I3(GND_net), .O(n44863));
    defparam i29978_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i17_4_lut (.I0(n5531), .I1(n44863), .I2(n6014), .I3(n37), 
            .O(n27956));
    defparam i17_4_lut.LUT_INIT = 16'h3a30;
    SB_DFFE enable_slow_120 (.Q(\state_7__N_3987[0] ), .C(CLK_c), .E(n27854), 
            .D(enable_slow_N_4089));   // verilog/i2c_controller.v(58[9] 71[5])
    SB_LUT4 counter2_1554_1555_add_4_7_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[5]), .I3(n40503), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1554_1555_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 counter2_1554_1555_add_4_6_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[4]), .I3(n40502), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1554_1555_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1554_1555_add_4_6 (.CI(n40502), .I0(GND_net), .I1(counter2[4]), 
            .CO(n40503));
    SB_LUT4 counter2_1554_1555_add_4_5_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[3]), .I3(n40501), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1554_1555_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1554_1555_add_4_5 (.CI(n40501), .I0(GND_net), .I1(counter2[3]), 
            .CO(n40502));
    SB_LUT4 counter2_1554_1555_add_4_4_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[2]), .I3(n40500), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1554_1555_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1554_1555_add_4_4 (.CI(n40500), .I0(GND_net), .I1(counter2[2]), 
            .CO(n40501));
    SB_LUT4 counter2_1554_1555_add_4_3_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[1]), .I3(n40499), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1554_1555_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1554_1555_add_4_3 (.CI(n40499), .I0(GND_net), .I1(counter2[1]), 
            .CO(n40500));
    SB_LUT4 counter2_1554_1555_add_4_2_lut (.I0(GND_net), .I1(GND_net), 
            .I2(counter2[0]), .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam counter2_1554_1555_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY counter2_1554_1555_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(counter2[0]), 
            .CO(n40499));
    SB_DFFNESS write_enable_131 (.Q(sda_enable), .C(i2c_clk), .E(n5909), 
            .D(n19384), .S(n28050));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_LUT4 equal_162_i4_2_lut (.I0(counter[1]), .I1(counter[2]), .I2(GND_net), 
            .I3(GND_net), .O(n4_adj_1));   // verilog/i2c_controller.v(153[6:23])
    defparam equal_162_i4_2_lut.LUT_INIT = 16'hdddd;
    SB_DFFNE sda_out_132 (.Q(sda_out_adj_4092), .C(i2c_clk), .E(n43769), 
            .D(n49887));   // verilog/i2c_controller.v(180[12] 215[6])
    SB_DFFESS counter_i0 (.Q(counter[0]), .C(i2c_clk), .E(n27956), .D(n119[0]), 
            .S(n28046));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i4_4_lut (.I0(counter2[3]), .I1(counter2[5]), .I2(counter2[2]), 
            .I3(counter2[4]), .O(n10_c));
    defparam i4_4_lut.LUT_INIT = 16'h8000;
    SB_LUT4 i5_3_lut (.I0(counter2[1]), .I1(n10_c), .I2(counter2[0]), 
            .I3(GND_net), .O(n28122));
    defparam i5_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i34943_2_lut (.I0(counter[1]), .I1(\saved_addr[0] ), .I2(GND_net), 
            .I3(GND_net), .O(n49774));   // verilog/i2c_controller.v(198[28:35])
    defparam i34943_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 i35087_4_lut (.I0(n49774), .I1(\state[1] ), .I2(counter[0]), 
            .I3(counter[2]), .O(n49716));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i35087_4_lut.LUT_INIT = 16'hc008;
    SB_LUT4 i35148_4_lut (.I0(n49716), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(n11), .O(n49887));   // verilog/i2c_controller.v(181[4] 214[11])
    defparam i35148_4_lut.LUT_INIT = 16'h0322;
    SB_LUT4 i1_4_lut (.I0(n11_adj_4093), .I1(n11_adj_4094), .I2(\state_7__N_4003[3] ), 
            .I3(\saved_addr[0] ), .O(n5));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut.LUT_INIT = 16'h5755;
    SB_LUT4 i35933_2_lut (.I0(\state_7__N_4003[3] ), .I1(n11_adj_4094), 
            .I2(GND_net), .I3(GND_net), .O(n33933));
    defparam i35933_2_lut.LUT_INIT = 16'h1111;
    SB_LUT4 state_7__I_0_143_i9_2_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(GND_net), .I3(GND_net), .O(n9));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i9_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i2_2_lut (.I0(counter[2]), .I1(counter[1]), .I2(GND_net), 
            .I3(GND_net), .O(n10));   // verilog/i2c_controller.v(110[10:22])
    defparam i2_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i5_4_lut (.I0(counter[3]), .I1(counter[5]), .I2(counter[0]), 
            .I3(counter[4]), .O(n12));   // verilog/i2c_controller.v(110[10:22])
    defparam i5_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i6_4_lut (.I0(counter[6]), .I1(n12), .I2(counter[7]), .I3(n10), 
            .O(n5531));   // verilog/i2c_controller.v(110[10:22])
    defparam i6_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(GND_net), 
            .I3(GND_net), .O(n7));
    defparam i1_2_lut.LUT_INIT = 16'h4444;
    SB_LUT4 state_7__I_0_143_i10_2_lut (.I0(\state[2] ), .I1(\state[3] ), 
            .I2(GND_net), .I3(GND_net), .O(n10_adj_2));   // verilog/i2c_controller.v(151[5:14])
    defparam state_7__I_0_143_i10_2_lut.LUT_INIT = 16'hdddd;
    SB_LUT4 i35753_4_lut (.I0(state_7__N_3986), .I1(n5531), .I2(n11_adj_4097), 
            .I3(n34056), .O(n5538));
    defparam i35753_4_lut.LUT_INIT = 16'h5111;
    SB_LUT4 i1_3_lut (.I0(\state[1] ), .I1(n33_adj_4098), .I2(n37), .I3(GND_net), 
            .O(n28050));
    defparam i1_3_lut.LUT_INIT = 16'h5454;
    SB_LUT4 i1_2_lut_adj_841 (.I0(n34_adj_4099), .I1(n37), .I2(GND_net), 
            .I3(GND_net), .O(n39));
    defparam i1_2_lut_adj_841.LUT_INIT = 16'heeee;
    SB_DFFE state_i0_i0 (.Q(\state[0] ), .C(i2c_clk), .E(VCC_net), .D(n8));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i0 (.Q(data[0]), .C(i2c_clk), .D(n28230));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i35012_4_lut (.I0(n10_adj_3), .I1(n10_adj_2), .I2(\state_7__N_4003[3] ), 
            .I3(enable), .O(n49793));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i35012_4_lut.LUT_INIT = 16'h7073;
    SB_LUT4 i35799_2_lut (.I0(\state_7__N_3987[0] ), .I1(enable_slow_N_4090), 
            .I2(GND_net), .I3(GND_net), .O(enable_slow_N_4089));   // verilog/i2c_controller.v(62[6:32])
    defparam i35799_2_lut.LUT_INIT = 16'h7777;
    SB_LUT4 i1_4_lut_adj_842 (.I0(\state[1] ), .I1(n7), .I2(n49793), .I3(\state[0] ), 
            .O(n43849));   // verilog/i2c_controller.v(92[4] 172[11])
    defparam i1_4_lut_adj_842.LUT_INIT = 16'ha088;
    SB_DFF saved_addr__i1 (.Q(\saved_addr[0] ), .C(i2c_clk), .D(n28224));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 i1_2_lut_adj_843 (.I0(i2c_clk), .I1(n28122), .I2(GND_net), 
            .I3(GND_net), .O(i2c_clk_N_4076));
    defparam i1_2_lut_adj_843.LUT_INIT = 16'h6666;
    SB_LUT4 i20617_2_lut (.I0(i2c_clk), .I1(scl_enable), .I2(GND_net), 
            .I3(GND_net), .O(scl));   // verilog/i2c_controller.v(45[19:61])
    defparam i20617_2_lut.LUT_INIT = 16'hbbbb;
    SB_LUT4 i1852_2_lut (.I0(sda_out_adj_4092), .I1(sda_enable), .I2(GND_net), 
            .I3(GND_net), .O(sda_out));   // verilog/i2c_controller.v(46[9:20])
    defparam i1852_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_2_lut_4_lut_4_lut (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(\state[0] ), .O(n34_adj_4099));
    defparam i1_2_lut_4_lut_4_lut.LUT_INIT = 16'h0510;
    SB_DFF data_out_i0_i1 (.Q(data[1]), .C(i2c_clk), .D(n28207));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i2 (.Q(data[2]), .C(i2c_clk), .D(n28206));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_LUT4 equal_103_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n15));   // verilog/i2c_controller.v(77[27:43])
    defparam equal_103_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffd;
    SB_LUT4 state_7__I_0_144_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4093));   // verilog/i2c_controller.v(77[27:43])
    defparam state_7__I_0_144_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hffdf;
    SB_LUT4 state_7__I_0_139_i11_2_lut_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4094));
    defparam state_7__I_0_139_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfff7;
    SB_LUT4 equal_101_i11_2_lut_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(enable_slow_N_4090));
    defparam equal_101_i11_2_lut_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_DFF data_out_i0_i3 (.Q(data[3]), .C(i2c_clk), .D(n28205));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i4 (.Q(data[4]), .C(i2c_clk), .D(n28204));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i5 (.Q(data[5]), .C(i2c_clk), .D(n28200));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i6 (.Q(data[6]), .C(i2c_clk), .D(n28199));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFF data_out_i0_i7 (.Q(data[7]), .C(i2c_clk), .D(n28198));   // verilog/i2c_controller.v(91[8] 173[6])
    SB_DFFSR counter2_1554_1555__i2 (.Q(counter2[1]), .C(CLK_c), .D(n29[1]), 
            .R(n28122));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1554_1555__i3 (.Q(counter2[2]), .C(CLK_c), .D(n29[2]), 
            .R(n28122));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1554_1555__i4 (.Q(counter2[3]), .C(CLK_c), .D(n29[3]), 
            .R(n28122));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1554_1555__i5 (.Q(counter2[4]), .C(CLK_c), .D(n29[4]), 
            .R(n28122));   // verilog/i2c_controller.v(69[20:35])
    SB_DFFSR counter2_1554_1555__i6 (.Q(counter2[5]), .C(CLK_c), .D(n29[5]), 
            .R(n28122));   // verilog/i2c_controller.v(69[20:35])
    SB_LUT4 i22_3_lut_3_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[3] ), 
            .I3(GND_net), .O(n11));
    defparam i22_3_lut_3_lut.LUT_INIT = 16'h1c1c;
    SB_LUT4 i21487_3_lut_4_lut (.I0(\state[1] ), .I1(\state[0] ), .I2(\state[2] ), 
            .I3(n15), .O(scl_enable_N_4077));
    defparam i21487_3_lut_4_lut.LUT_INIT = 16'hfe00;
    SB_LUT4 sub_39_add_2_9_lut (.I0(GND_net), .I1(counter[7]), .I2(VCC_net), 
            .I3(n39365), .O(n119[7])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 sub_39_add_2_8_lut (.I0(GND_net), .I1(counter[6]), .I2(VCC_net), 
            .I3(n39364), .O(n119[6])) /* synthesis syn_instantiated=1 */ ;
    defparam sub_39_add_2_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i35810_4_lut_4_lut (.I0(\state[2] ), .I1(n11), .I2(\state[1] ), 
            .I3(n39), .O(n5909));
    defparam i35810_4_lut_4_lut.LUT_INIT = 16'hef00;
    SB_LUT4 i35835_2_lut_3_lut (.I0(\state[2] ), .I1(n11), .I2(\state[0] ), 
            .I3(GND_net), .O(n19384));
    defparam i35835_2_lut_3_lut.LUT_INIT = 16'h0404;
    SB_LUT4 i21522_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(state_7__N_3986));
    defparam i21522_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 i1_2_lut_3_lut (.I0(n9), .I1(n10_adj_2), .I2(counter[0]), 
            .I3(GND_net), .O(n26650));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hefef;
    SB_LUT4 i1_2_lut_3_lut_adj_844 (.I0(n9), .I1(n10_adj_2), .I2(counter[0]), 
            .I3(GND_net), .O(n26645));   // verilog/i2c_controller.v(151[5:14])
    defparam i1_2_lut_3_lut_adj_844.LUT_INIT = 16'hfefe;
    SB_LUT4 i36098_3_lut_4_lut (.I0(n9), .I1(n10_adj_2), .I2(n11_adj_4101), 
            .I3(n5538), .O(n34177));   // verilog/i2c_controller.v(151[5:14])
    defparam i36098_3_lut_4_lut.LUT_INIT = 16'h1f00;
    SB_CARRY sub_39_add_2_8 (.CI(n39364), .I0(counter[6]), .I1(VCC_net), 
            .CO(n39365));
    SB_LUT4 i2_3_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[3] ), .O(n11_adj_4101));   // verilog/i2c_controller.v(77[27:43])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfdff;
    SB_LUT4 i35094_3_lut_4_lut (.I0(n11_adj_4097), .I1(n11_adj_4101), .I2(enable_slow_N_4090), 
            .I3(\state_7__N_3987[0] ), .O(n49785));
    defparam i35094_3_lut_4_lut.LUT_INIT = 16'h8088;
    SB_LUT4 i35957_3_lut_4_lut (.I0(n11_adj_4097), .I1(n11_adj_4101), .I2(n15), 
            .I3(n5538), .O(n34447));
    defparam i35957_3_lut_4_lut.LUT_INIT = 16'h7f00;
    SB_LUT4 i35804_4_lut_4_lut (.I0(\state[1] ), .I1(\state[2] ), .I2(\state[0] ), 
            .I3(\state[3] ), .O(n43769));
    defparam i35804_4_lut_4_lut.LUT_INIT = 16'h0156;
    SB_LUT4 i1_2_lut_3_lut_adj_845 (.I0(enable), .I1(\state_7__N_3987[0] ), 
            .I2(enable_slow_N_4090), .I3(GND_net), .O(n27854));
    defparam i1_2_lut_3_lut_adj_845.LUT_INIT = 16'heaea;
    SB_LUT4 i56_3_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n33_adj_4098));
    defparam i56_3_lut_3_lut.LUT_INIT = 16'h3434;
    SB_LUT4 i36101_3_lut_4_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[1] ), 
            .I3(n5538), .O(n46193));
    defparam i36101_3_lut_4_lut.LUT_INIT = 16'h0200;
    SB_LUT4 state_7__I_0_138_i11_2_lut_4_lut (.I0(\state[0] ), .I1(\state[1] ), 
            .I2(\state[2] ), .I3(\state[3] ), .O(n11_adj_4097));   // verilog/i2c_controller.v(109[5:12])
    defparam state_7__I_0_138_i11_2_lut_4_lut.LUT_INIT = 16'hfffb;
    SB_LUT4 i21001_2_lut_3_lut (.I0(\state[2] ), .I1(\state[3] ), .I2(\state[0] ), 
            .I3(GND_net), .O(n34056));
    defparam i21001_2_lut_3_lut.LUT_INIT = 16'hfdfd;
    SB_LUT4 i29916_2_lut_4_lut (.I0(\state[0] ), .I1(\state[2] ), .I2(\state[3] ), 
            .I3(n44863), .O(n28046));   // verilog/i2c_controller.v(91[8] 173[6])
    defparam i29916_2_lut_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i1_2_lut_4_lut (.I0(\state[3] ), .I1(\state[1] ), .I2(\state[2] ), 
            .I3(\state[0] ), .O(n37));
    defparam i1_2_lut_4_lut.LUT_INIT = 16'h0554;
    
endmodule
//
// Verilog Description of module pwm
//

module pwm (n50560, VCC_net, INHA_c, clk32MHz, n26492, GND_net, 
            pwm_counter, n26490) /* synthesis syn_module_defined=1 */ ;
    input n50560;
    input VCC_net;
    output INHA_c;
    input clk32MHz;
    input n26492;
    input GND_net;
    output [31:0]pwm_counter;
    input n26490;
    
    wire clk32MHz /* synthesis SET_AS_NETWORK=clk32MHz, is_clock=1 */ ;   // verilog/TinyFPGA_B.v(33[6:14])
    wire [31:0]n133;
    
    wire n40421, n40420, n40419, n40418, n40417, n40416, n40415, 
        n40414, n40413, n40412, n40411, n40410, n40409, n40408, 
        n40407, n40406, n40405, n40404, n40403, n40402, n40401, 
        n40400, n40399, n40398, n40397, n40396, n40395, n40394, 
        n40393, n40392, n40391, pwm_counter_31__N_711, n46147, n18, 
        n24, n22, n26, n21;
    
    SB_DFFESR pwm_out_12 (.Q(INHA_c), .C(clk32MHz), .E(VCC_net), .D(n50560), 
            .R(n26492));   // verilog/pwm.v(16[12] 26[6])
    SB_LUT4 pwm_counter_1547_add_4_33_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[31]), 
            .I3(n40421), .O(n133[31])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_33_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 pwm_counter_1547_add_4_32_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[30]), 
            .I3(n40420), .O(n133[30])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_32_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_32 (.CI(n40420), .I0(GND_net), .I1(pwm_counter[30]), 
            .CO(n40421));
    SB_LUT4 pwm_counter_1547_add_4_31_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[29]), 
            .I3(n40419), .O(n133[29])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_31_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_31 (.CI(n40419), .I0(GND_net), .I1(pwm_counter[29]), 
            .CO(n40420));
    SB_LUT4 pwm_counter_1547_add_4_30_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[28]), 
            .I3(n40418), .O(n133[28])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_30_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_30 (.CI(n40418), .I0(GND_net), .I1(pwm_counter[28]), 
            .CO(n40419));
    SB_LUT4 pwm_counter_1547_add_4_29_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[27]), 
            .I3(n40417), .O(n133[27])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_29_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_29 (.CI(n40417), .I0(GND_net), .I1(pwm_counter[27]), 
            .CO(n40418));
    SB_LUT4 pwm_counter_1547_add_4_28_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[26]), 
            .I3(n40416), .O(n133[26])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_28_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_28 (.CI(n40416), .I0(GND_net), .I1(pwm_counter[26]), 
            .CO(n40417));
    SB_LUT4 pwm_counter_1547_add_4_27_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[25]), 
            .I3(n40415), .O(n133[25])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_27_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_27 (.CI(n40415), .I0(GND_net), .I1(pwm_counter[25]), 
            .CO(n40416));
    SB_LUT4 pwm_counter_1547_add_4_26_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[24]), 
            .I3(n40414), .O(n133[24])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_26_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_26 (.CI(n40414), .I0(GND_net), .I1(pwm_counter[24]), 
            .CO(n40415));
    SB_LUT4 pwm_counter_1547_add_4_25_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[23]), 
            .I3(n40413), .O(n133[23])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_25_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_25 (.CI(n40413), .I0(GND_net), .I1(pwm_counter[23]), 
            .CO(n40414));
    SB_LUT4 pwm_counter_1547_add_4_24_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[22]), 
            .I3(n40412), .O(n133[22])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_24_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_24 (.CI(n40412), .I0(GND_net), .I1(pwm_counter[22]), 
            .CO(n40413));
    SB_LUT4 pwm_counter_1547_add_4_23_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[21]), 
            .I3(n40411), .O(n133[21])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_23_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_23 (.CI(n40411), .I0(GND_net), .I1(pwm_counter[21]), 
            .CO(n40412));
    SB_LUT4 pwm_counter_1547_add_4_22_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[20]), 
            .I3(n40410), .O(n133[20])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_22_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_22 (.CI(n40410), .I0(GND_net), .I1(pwm_counter[20]), 
            .CO(n40411));
    SB_LUT4 pwm_counter_1547_add_4_21_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[19]), 
            .I3(n40409), .O(n133[19])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_21_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_21 (.CI(n40409), .I0(GND_net), .I1(pwm_counter[19]), 
            .CO(n40410));
    SB_LUT4 pwm_counter_1547_add_4_20_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[18]), 
            .I3(n40408), .O(n133[18])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_20_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_20 (.CI(n40408), .I0(GND_net), .I1(pwm_counter[18]), 
            .CO(n40409));
    SB_LUT4 pwm_counter_1547_add_4_19_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[17]), 
            .I3(n40407), .O(n133[17])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_19_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_19 (.CI(n40407), .I0(GND_net), .I1(pwm_counter[17]), 
            .CO(n40408));
    SB_LUT4 pwm_counter_1547_add_4_18_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[16]), 
            .I3(n40406), .O(n133[16])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_18_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_18 (.CI(n40406), .I0(GND_net), .I1(pwm_counter[16]), 
            .CO(n40407));
    SB_LUT4 pwm_counter_1547_add_4_17_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[15]), 
            .I3(n40405), .O(n133[15])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_17_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_17 (.CI(n40405), .I0(GND_net), .I1(pwm_counter[15]), 
            .CO(n40406));
    SB_LUT4 pwm_counter_1547_add_4_16_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[14]), 
            .I3(n40404), .O(n133[14])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_16_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_16 (.CI(n40404), .I0(GND_net), .I1(pwm_counter[14]), 
            .CO(n40405));
    SB_LUT4 pwm_counter_1547_add_4_15_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[13]), 
            .I3(n40403), .O(n133[13])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_15 (.CI(n40403), .I0(GND_net), .I1(pwm_counter[13]), 
            .CO(n40404));
    SB_LUT4 pwm_counter_1547_add_4_14_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[12]), 
            .I3(n40402), .O(n133[12])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_14_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_14 (.CI(n40402), .I0(GND_net), .I1(pwm_counter[12]), 
            .CO(n40403));
    SB_LUT4 pwm_counter_1547_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[11]), 
            .I3(n40401), .O(n133[11])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_13 (.CI(n40401), .I0(GND_net), .I1(pwm_counter[11]), 
            .CO(n40402));
    SB_LUT4 pwm_counter_1547_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[10]), 
            .I3(n40400), .O(n133[10])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_12 (.CI(n40400), .I0(GND_net), .I1(pwm_counter[10]), 
            .CO(n40401));
    SB_LUT4 pwm_counter_1547_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[9]), 
            .I3(n40399), .O(n133[9])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_11 (.CI(n40399), .I0(GND_net), .I1(pwm_counter[9]), 
            .CO(n40400));
    SB_LUT4 pwm_counter_1547_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[8]), 
            .I3(n40398), .O(n133[8])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_10 (.CI(n40398), .I0(GND_net), .I1(pwm_counter[8]), 
            .CO(n40399));
    SB_LUT4 pwm_counter_1547_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[7]), 
            .I3(n40397), .O(n133[7])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_9 (.CI(n40397), .I0(GND_net), .I1(pwm_counter[7]), 
            .CO(n40398));
    SB_LUT4 pwm_counter_1547_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[6]), 
            .I3(n40396), .O(n133[6])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_8 (.CI(n40396), .I0(GND_net), .I1(pwm_counter[6]), 
            .CO(n40397));
    SB_LUT4 pwm_counter_1547_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[5]), 
            .I3(n40395), .O(n133[5])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_7 (.CI(n40395), .I0(GND_net), .I1(pwm_counter[5]), 
            .CO(n40396));
    SB_LUT4 pwm_counter_1547_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[4]), 
            .I3(n40394), .O(n133[4])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_6 (.CI(n40394), .I0(GND_net), .I1(pwm_counter[4]), 
            .CO(n40395));
    SB_LUT4 pwm_counter_1547_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[3]), 
            .I3(n40393), .O(n133[3])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_5 (.CI(n40393), .I0(GND_net), .I1(pwm_counter[3]), 
            .CO(n40394));
    SB_LUT4 pwm_counter_1547_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[2]), 
            .I3(n40392), .O(n133[2])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_4 (.CI(n40392), .I0(GND_net), .I1(pwm_counter[2]), 
            .CO(n40393));
    SB_LUT4 pwm_counter_1547_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[1]), 
            .I3(n40391), .O(n133[1])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_3 (.CI(n40391), .I0(GND_net), .I1(pwm_counter[1]), 
            .CO(n40392));
    SB_LUT4 pwm_counter_1547_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(pwm_counter[0]), 
            .I3(VCC_net), .O(n133[0])) /* synthesis syn_instantiated=1 */ ;
    defparam pwm_counter_1547_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY pwm_counter_1547_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(pwm_counter[0]), 
            .CO(n40391));
    SB_DFFSR pwm_counter_1547__i0 (.Q(pwm_counter[0]), .C(clk32MHz), .D(n133[0]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i1 (.Q(pwm_counter[1]), .C(clk32MHz), .D(n133[1]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i2 (.Q(pwm_counter[2]), .C(clk32MHz), .D(n133[2]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i3 (.Q(pwm_counter[3]), .C(clk32MHz), .D(n133[3]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i4 (.Q(pwm_counter[4]), .C(clk32MHz), .D(n133[4]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i5 (.Q(pwm_counter[5]), .C(clk32MHz), .D(n133[5]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i6 (.Q(pwm_counter[6]), .C(clk32MHz), .D(n133[6]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i7 (.Q(pwm_counter[7]), .C(clk32MHz), .D(n133[7]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i8 (.Q(pwm_counter[8]), .C(clk32MHz), .D(n133[8]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i9 (.Q(pwm_counter[9]), .C(clk32MHz), .D(n133[9]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i10 (.Q(pwm_counter[10]), .C(clk32MHz), .D(n133[10]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i11 (.Q(pwm_counter[11]), .C(clk32MHz), .D(n133[11]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i12 (.Q(pwm_counter[12]), .C(clk32MHz), .D(n133[12]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i13 (.Q(pwm_counter[13]), .C(clk32MHz), .D(n133[13]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i14 (.Q(pwm_counter[14]), .C(clk32MHz), .D(n133[14]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i15 (.Q(pwm_counter[15]), .C(clk32MHz), .D(n133[15]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i16 (.Q(pwm_counter[16]), .C(clk32MHz), .D(n133[16]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i17 (.Q(pwm_counter[17]), .C(clk32MHz), .D(n133[17]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i18 (.Q(pwm_counter[18]), .C(clk32MHz), .D(n133[18]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i19 (.Q(pwm_counter[19]), .C(clk32MHz), .D(n133[19]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i20 (.Q(pwm_counter[20]), .C(clk32MHz), .D(n133[20]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i21 (.Q(pwm_counter[21]), .C(clk32MHz), .D(n133[21]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i22 (.Q(pwm_counter[22]), .C(clk32MHz), .D(n133[22]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i23 (.Q(pwm_counter[23]), .C(clk32MHz), .D(n133[23]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i24 (.Q(pwm_counter[24]), .C(clk32MHz), .D(n133[24]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i25 (.Q(pwm_counter[25]), .C(clk32MHz), .D(n133[25]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i26 (.Q(pwm_counter[26]), .C(clk32MHz), .D(n133[26]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i27 (.Q(pwm_counter[27]), .C(clk32MHz), .D(n133[27]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i28 (.Q(pwm_counter[28]), .C(clk32MHz), .D(n133[28]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i29 (.Q(pwm_counter[29]), .C(clk32MHz), .D(n133[29]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i30 (.Q(pwm_counter[30]), .C(clk32MHz), .D(n133[30]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_DFFSR pwm_counter_1547__i31 (.Q(pwm_counter[31]), .C(clk32MHz), .D(n133[31]), 
            .R(pwm_counter_31__N_711));   // verilog/pwm.v(17[20:33])
    SB_LUT4 i2_3_lut (.I0(pwm_counter[6]), .I1(pwm_counter[8]), .I2(pwm_counter[7]), 
            .I3(GND_net), .O(n46147));
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut (.I0(n46147), .I1(pwm_counter[13]), .I2(pwm_counter[10]), 
            .I3(pwm_counter[9]), .O(n18));
    defparam i4_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i10_4_lut (.I0(pwm_counter[17]), .I1(pwm_counter[22]), .I2(pwm_counter[14]), 
            .I3(pwm_counter[18]), .O(n24));
    defparam i10_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i8_4_lut (.I0(pwm_counter[21]), .I1(n26490), .I2(pwm_counter[16]), 
            .I3(pwm_counter[12]), .O(n22));
    defparam i8_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i12_4_lut (.I0(pwm_counter[15]), .I1(n24), .I2(n18), .I3(pwm_counter[19]), 
            .O(n26));
    defparam i12_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i7_2_lut (.I0(pwm_counter[11]), .I1(pwm_counter[20]), .I2(GND_net), 
            .I3(GND_net), .O(n21));
    defparam i7_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i20814_4_lut (.I0(n21), .I1(pwm_counter[31]), .I2(n26), .I3(n22), 
            .O(pwm_counter_31__N_711));   // verilog/pwm.v(18[8:40])
    defparam i20814_4_lut.LUT_INIT = 16'h3332;
    
endmodule
